-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 755;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (3,0,65,0,215,0,0,0,98,0,60,0,138,0,192,0,0,0,0,0,89,0,62,0,162,0,168,0,132,0,106,0,98,0,67,0,0,0,252,0,204,0,156,0,52,0,253,0,0,0,106,0,0,0,1,0,150,0,0,0,235,0,96,0,65,0,116,0,89,0,131,0,71,0,202,0,157,0,27,0,54,0,201,0,176,0,59,0,98,0,0,0,201,0,147,0,0,0,33,0,223,0,206,0,137,0,163,0,26,0,253,0,0,0,0,0,151,0,84,0,219,0,52,0,96,0,0,0,0,0,51,0,0,0,0,0,41,0,2,0,207,0,0,0,132,0,1,0,109,0,146,0,0,0,0,0,0,0,79,0,169,0,137,0,138,0,0,0,131,0,0,0,189,0,0,0,157,0,183,0,0,0,246,0,0,0,0,0,111,0,79,0,195,0,0,0,8,0,147,0,141,0,70,0,0,0,187,0,131,0,196,0,0,0,166,0,123,0,46,0,122,0,79,0,0,0,192,0,180,0,0,0,107,0,69,0,44,0,87,0,199,0,57,0,253,0,0,0,101,0,60,0,155,0,0,0,222,0,22,0,0,0,134,0,254,0,20,0,126,0,0,0,0,0,218,0,143,0,205,0,107,0,20,0,141,0,213,0,0,0,249,0,12,0,76,0,242,0,254,0,67,0,168,0,98,0,45,0,0,0,32,0,0,0,120,0,83,0,123,0,131,0,152,0,213,0,0,0,15,0,186,0,9,0,0,0,217,0,0,0,232,0,161,0,73,0,0,0,92,0,239,0,177,0,1,0,0,0,11,0,24,0,29,0,0,0,0,0,0,0,1,0,58,0,29,0,160,0,59,0,147,0,17,0,114,0,8,0,14,0,200,0,99,0,173,0,170,0,50,0,63,0,34,0,0,0,167,0,225,0,45,0,171,0,251,0,0,0,0,0,0,0,227,0,104,0,125,0,93,0,14,0,61,0,178,0,138,0,0,0,78,0,0,0,245,0,0,0,0,0,255,0,136,0,19,0,148,0,0,0,0,0,191,0,77,0,0,0,166,0,0,0,252,0,0,0,45,0,0,0,0,0,7,0,170,0,171,0,199,0,123,0,90,0,46,0,25,0,116,0,218,0,9,0,0,0,204,0,103,0,71,0,194,0,0,0,51,0,60,0,0,0,142,0,47,0,0,0,0,0,50,0,223,0,208,0,78,0,205,0,0,0,116,0,37,0,0,0,0,0,138,0,255,0,147,0,103,0,7,0,93,0,150,0,167,0,90,0,67,0,0,0,249,0,0,0,123,0,14,0,246,0,130,0,169,0,175,0,213,0,14,0,102,0,216,0,0,0,0,0,15,0,0,0,159,0,15,0,0,0,0,0,79,0,254,0,148,0,0,0,50,0,0,0,244,0,114,0,81,0,134,0,0,0,0,0,33,0,27,0,0,0,252,0,130,0,85,0,82,0,190,0,149,0,222,0,119,0,126,0,81,0,98,0,120,0,38,0,80,0,12,0,105,0,1,0,45,0,135,0,70,0,199,0,224,0,86,0,0,0,0,0,0,0,178,0,32,0,123,0,209,0,22,0,0,0,27,0,249,0,8,0,159,0,238,0,232,0,83,0,0,0,128,0,82,0,227,0,43,0,148,0,169,0,119,0,0,0,145,0,17,0,78,0,253,0,226,0,41,0,163,0,0,0,113,0,6,0,0,0,0,0,0,0,151,0,120,0,176,0,120,0,251,0,69,0,205,0,103,0,0,0,31,0,0,0,13,0,0,0,53,0,129,0,57,0,0,0,122,0,40,0,188,0,0,0,0,0,158,0,43,0,120,0,0,0,207,0,0,0,0,0,0,0,177,0,47,0,0,0,230,0,77,0,143,0,28,0,0,0,141,0,165,0,244,0,25,0,54,0,54,0,0,0,248,0,0,0,255,0,79,0,121,0,0,0,72,0,228,0,0,0,0,0,99,0,0,0,126,0,67,0,206,0,0,0,2,0,0,0,229,0,238,0,110,0,132,0,72,0,116,0,43,0,123,0,189,0,137,0,153,0,0,0,148,0,17,0,0,0,118,0,0,0,3,0,0,0,0,0,226,0,98,0,0,0,238,0,22,0,113,0,51,0,0,0,171,0,0,0,133,0,30,0,162,0,0,0,234,0,170,0,0,0,77,0,0,0,243,0,64,0,47,0,72,0,245,0,172,0,11,0,77,0,151,0,171,0,15,0,121,0,0,0,252,0,59,0,0,0,71,0,0,0,125,0,35,0,59,0,119,0,219,0,90,0,193,0,84,0,14,0,0,0,166,0,35,0,123,0,0,0,59,0,0,0,27,0,160,0,0,0,114,0,38,0,69,0,241,0,46,0,187,0,202,0,149,0,164,0,0,0,73,0,200,0,168,0,112,0,235,0,35,0,0,0,0,0,178,0,0,0,0,0,0,0,168,0,0,0,42,0,0,0,20,0,184,0,90,0,0,0,0,0,15,0,198,0,2,0,0,0,191,0,160,0,0,0,126,0,98,0,243,0,137,0,151,0,134,0,236,0,126,0,0,0,205,0,24,0,22,0,114,0,0,0,216,0,200,0,26,0,91,0,26,0,126,0,112,0,32,0,125,0,89,0,0,0,215,0,156,0,122,0,79,0,204,0,0,0,9,0,0,0,25,0,0,0,0,0,55,0,224,0,11,0,0,0,249,0,0,0,42,0,188,0,42,0,0,0,86,0,179,0,3,0,89,0,5,0,144,0,18,0,241,0,171,0,229,0,77,0,0,0,216,0,161,0,0,0,136,0,16,0,149,0,0,0,3,0,210,0,197,0,103,0,8,0,225,0,0,0,90,0,142,0,237,0,98,0,6,0,0,0,43,0,254,0,239,0,0,0,54,0,104,0,87,0,149,0,2,0,0,0,242,0,0,0,254,0,178,0,0,0,52,0,0,0,10,0,148,0,29,0,0,0,189,0,182,0,65,0,0,0,147,0,114,0,190,0,83,0,86,0,0,0,0,0,140,0,7,0,0,0,0,0,0,0,73,0,147,0,155,0,32,0,119,0,0,0,0,0,154,0,0,0,0,0,40,0,0,0,0,0,0,0,0,0,177,0,184,0,163,0,123,0,233,0,208,0,184,0,217,0,59,0,229,0,24,0,134,0,13,0,198,0,159,0,0,0,0,0,247,0,187,0,0,0,31,0,194,0,19,0,85,0,25,0,215,0,70,0,185,0,0,0,155,0,223,0,150,0,103,0,0,0,248,0,0,0,40,0,115,0,111,0,103,0,119,0,151,0,0,0,249,0,188,0,108,0,35,0,0,0,0,0,165,0,0,0,84,0,0,0,26,0,0,0,231,0,157,0,11,0,70,0,14,0,226,0,10,0,162,0,112,0,62,0,208,0);
signal scenario_full  : scenario_type := (3,31,65,31,215,31,215,30,98,31,60,31,138,31,192,31,192,30,192,29,89,31,62,31,162,31,168,31,132,31,106,31,98,31,67,31,67,30,252,31,204,31,156,31,52,31,253,31,253,30,106,31,106,30,1,31,150,31,150,30,235,31,96,31,65,31,116,31,89,31,131,31,71,31,202,31,157,31,27,31,54,31,201,31,176,31,59,31,98,31,98,30,201,31,147,31,147,30,33,31,223,31,206,31,137,31,163,31,26,31,253,31,253,30,253,29,151,31,84,31,219,31,52,31,96,31,96,30,96,29,51,31,51,30,51,29,41,31,2,31,207,31,207,30,132,31,1,31,109,31,146,31,146,30,146,29,146,28,79,31,169,31,137,31,138,31,138,30,131,31,131,30,189,31,189,30,157,31,183,31,183,30,246,31,246,30,246,29,111,31,79,31,195,31,195,30,8,31,147,31,141,31,70,31,70,30,187,31,131,31,196,31,196,30,166,31,123,31,46,31,122,31,79,31,79,30,192,31,180,31,180,30,107,31,69,31,44,31,87,31,199,31,57,31,253,31,253,30,101,31,60,31,155,31,155,30,222,31,22,31,22,30,134,31,254,31,20,31,126,31,126,30,126,29,218,31,143,31,205,31,107,31,20,31,141,31,213,31,213,30,249,31,12,31,76,31,242,31,254,31,67,31,168,31,98,31,45,31,45,30,32,31,32,30,120,31,83,31,123,31,131,31,152,31,213,31,213,30,15,31,186,31,9,31,9,30,217,31,217,30,232,31,161,31,73,31,73,30,92,31,239,31,177,31,1,31,1,30,11,31,24,31,29,31,29,30,29,29,29,28,1,31,58,31,29,31,160,31,59,31,147,31,17,31,114,31,8,31,14,31,200,31,99,31,173,31,170,31,50,31,63,31,34,31,34,30,167,31,225,31,45,31,171,31,251,31,251,30,251,29,251,28,227,31,104,31,125,31,93,31,14,31,61,31,178,31,138,31,138,30,78,31,78,30,245,31,245,30,245,29,255,31,136,31,19,31,148,31,148,30,148,29,191,31,77,31,77,30,166,31,166,30,252,31,252,30,45,31,45,30,45,29,7,31,170,31,171,31,199,31,123,31,90,31,46,31,25,31,116,31,218,31,9,31,9,30,204,31,103,31,71,31,194,31,194,30,51,31,60,31,60,30,142,31,47,31,47,30,47,29,50,31,223,31,208,31,78,31,205,31,205,30,116,31,37,31,37,30,37,29,138,31,255,31,147,31,103,31,7,31,93,31,150,31,167,31,90,31,67,31,67,30,249,31,249,30,123,31,14,31,246,31,130,31,169,31,175,31,213,31,14,31,102,31,216,31,216,30,216,29,15,31,15,30,159,31,15,31,15,30,15,29,79,31,254,31,148,31,148,30,50,31,50,30,244,31,114,31,81,31,134,31,134,30,134,29,33,31,27,31,27,30,252,31,130,31,85,31,82,31,190,31,149,31,222,31,119,31,126,31,81,31,98,31,120,31,38,31,80,31,12,31,105,31,1,31,45,31,135,31,70,31,199,31,224,31,86,31,86,30,86,29,86,28,178,31,32,31,123,31,209,31,22,31,22,30,27,31,249,31,8,31,159,31,238,31,232,31,83,31,83,30,128,31,82,31,227,31,43,31,148,31,169,31,119,31,119,30,145,31,17,31,78,31,253,31,226,31,41,31,163,31,163,30,113,31,6,31,6,30,6,29,6,28,151,31,120,31,176,31,120,31,251,31,69,31,205,31,103,31,103,30,31,31,31,30,13,31,13,30,53,31,129,31,57,31,57,30,122,31,40,31,188,31,188,30,188,29,158,31,43,31,120,31,120,30,207,31,207,30,207,29,207,28,177,31,47,31,47,30,230,31,77,31,143,31,28,31,28,30,141,31,165,31,244,31,25,31,54,31,54,31,54,30,248,31,248,30,255,31,79,31,121,31,121,30,72,31,228,31,228,30,228,29,99,31,99,30,126,31,67,31,206,31,206,30,2,31,2,30,229,31,238,31,110,31,132,31,72,31,116,31,43,31,123,31,189,31,137,31,153,31,153,30,148,31,17,31,17,30,118,31,118,30,3,31,3,30,3,29,226,31,98,31,98,30,238,31,22,31,113,31,51,31,51,30,171,31,171,30,133,31,30,31,162,31,162,30,234,31,170,31,170,30,77,31,77,30,243,31,64,31,47,31,72,31,245,31,172,31,11,31,77,31,151,31,171,31,15,31,121,31,121,30,252,31,59,31,59,30,71,31,71,30,125,31,35,31,59,31,119,31,219,31,90,31,193,31,84,31,14,31,14,30,166,31,35,31,123,31,123,30,59,31,59,30,27,31,160,31,160,30,114,31,38,31,69,31,241,31,46,31,187,31,202,31,149,31,164,31,164,30,73,31,200,31,168,31,112,31,235,31,35,31,35,30,35,29,178,31,178,30,178,29,178,28,168,31,168,30,42,31,42,30,20,31,184,31,90,31,90,30,90,29,15,31,198,31,2,31,2,30,191,31,160,31,160,30,126,31,98,31,243,31,137,31,151,31,134,31,236,31,126,31,126,30,205,31,24,31,22,31,114,31,114,30,216,31,200,31,26,31,91,31,26,31,126,31,112,31,32,31,125,31,89,31,89,30,215,31,156,31,122,31,79,31,204,31,204,30,9,31,9,30,25,31,25,30,25,29,55,31,224,31,11,31,11,30,249,31,249,30,42,31,188,31,42,31,42,30,86,31,179,31,3,31,89,31,5,31,144,31,18,31,241,31,171,31,229,31,77,31,77,30,216,31,161,31,161,30,136,31,16,31,149,31,149,30,3,31,210,31,197,31,103,31,8,31,225,31,225,30,90,31,142,31,237,31,98,31,6,31,6,30,43,31,254,31,239,31,239,30,54,31,104,31,87,31,149,31,2,31,2,30,242,31,242,30,254,31,178,31,178,30,52,31,52,30,10,31,148,31,29,31,29,30,189,31,182,31,65,31,65,30,147,31,114,31,190,31,83,31,86,31,86,30,86,29,140,31,7,31,7,30,7,29,7,28,73,31,147,31,155,31,32,31,119,31,119,30,119,29,154,31,154,30,154,29,40,31,40,30,40,29,40,28,40,27,177,31,184,31,163,31,123,31,233,31,208,31,184,31,217,31,59,31,229,31,24,31,134,31,13,31,198,31,159,31,159,30,159,29,247,31,187,31,187,30,31,31,194,31,19,31,85,31,25,31,215,31,70,31,185,31,185,30,155,31,223,31,150,31,103,31,103,30,248,31,248,30,40,31,115,31,111,31,103,31,119,31,151,31,151,30,249,31,188,31,108,31,35,31,35,30,35,29,165,31,165,30,84,31,84,30,26,31,26,30,231,31,157,31,11,31,70,31,14,31,226,31,10,31,162,31,112,31,62,31,208,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
