-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 953;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (24,0,138,0,9,0,33,0,130,0,167,0,66,0,8,0,0,0,37,0,62,0,0,0,230,0,68,0,50,0,71,0,130,0,10,0,45,0,118,0,0,0,98,0,38,0,224,0,59,0,0,0,180,0,0,0,0,0,0,0,115,0,88,0,0,0,103,0,255,0,21,0,0,0,94,0,0,0,89,0,0,0,5,0,3,0,0,0,0,0,206,0,215,0,156,0,0,0,158,0,127,0,189,0,99,0,0,0,82,0,0,0,43,0,46,0,196,0,182,0,74,0,29,0,0,0,38,0,150,0,137,0,0,0,89,0,60,0,0,0,0,0,79,0,241,0,181,0,170,0,243,0,164,0,129,0,115,0,169,0,0,0,55,0,238,0,191,0,13,0,0,0,214,0,44,0,0,0,104,0,167,0,168,0,228,0,172,0,185,0,0,0,74,0,0,0,240,0,159,0,0,0,0,0,163,0,43,0,10,0,0,0,250,0,162,0,0,0,115,0,255,0,67,0,156,0,235,0,219,0,0,0,57,0,142,0,16,0,160,0,129,0,0,0,0,0,0,0,30,0,0,0,215,0,140,0,223,0,136,0,192,0,171,0,15,0,28,0,62,0,80,0,91,0,0,0,242,0,136,0,6,0,138,0,120,0,223,0,22,0,114,0,137,0,0,0,0,0,118,0,0,0,47,0,225,0,253,0,216,0,92,0,168,0,9,0,53,0,191,0,237,0,0,0,138,0,182,0,214,0,196,0,79,0,150,0,178,0,252,0,36,0,243,0,229,0,253,0,19,0,60,0,0,0,96,0,0,0,135,0,0,0,0,0,96,0,88,0,0,0,167,0,25,0,61,0,101,0,0,0,28,0,53,0,234,0,171,0,64,0,173,0,29,0,43,0,150,0,42,0,0,0,109,0,0,0,128,0,158,0,217,0,120,0,0,0,184,0,182,0,29,0,81,0,0,0,0,0,130,0,167,0,210,0,164,0,94,0,236,0,167,0,49,0,230,0,167,0,0,0,130,0,0,0,11,0,104,0,249,0,115,0,63,0,80,0,45,0,111,0,77,0,96,0,0,0,160,0,183,0,133,0,146,0,178,0,54,0,42,0,0,0,188,0,255,0,223,0,230,0,203,0,0,0,0,0,168,0,151,0,175,0,172,0,65,0,14,0,68,0,74,0,105,0,202,0,112,0,63,0,234,0,0,0,0,0,159,0,150,0,213,0,208,0,43,0,159,0,118,0,0,0,221,0,187,0,0,0,235,0,227,0,75,0,0,0,0,0,0,0,135,0,70,0,115,0,0,0,172,0,166,0,0,0,58,0,0,0,0,0,0,0,214,0,93,0,0,0,247,0,240,0,188,0,0,0,85,0,67,0,135,0,43,0,0,0,141,0,50,0,247,0,0,0,0,0,117,0,0,0,0,0,141,0,7,0,0,0,69,0,132,0,171,0,183,0,214,0,0,0,153,0,130,0,39,0,254,0,0,0,164,0,109,0,215,0,98,0,64,0,33,0,255,0,27,0,0,0,0,0,112,0,12,0,29,0,122,0,0,0,93,0,179,0,101,0,137,0,210,0,47,0,0,0,131,0,101,0,72,0,228,0,106,0,203,0,0,0,59,0,149,0,196,0,49,0,111,0,159,0,192,0,0,0,255,0,29,0,105,0,58,0,25,0,67,0,23,0,46,0,132,0,205,0,0,0,159,0,220,0,190,0,166,0,68,0,20,0,160,0,155,0,250,0,106,0,152,0,0,0,149,0,241,0,207,0,147,0,70,0,78,0,29,0,159,0,0,0,0,0,141,0,10,0,127,0,86,0,80,0,23,0,0,0,10,0,0,0,200,0,61,0,0,0,0,0,248,0,25,0,182,0,0,0,198,0,0,0,225,0,249,0,29,0,151,0,252,0,187,0,9,0,178,0,174,0,248,0,223,0,82,0,12,0,157,0,13,0,232,0,140,0,125,0,17,0,252,0,104,0,71,0,40,0,160,0,10,0,59,0,133,0,159,0,0,0,168,0,59,0,150,0,43,0,70,0,0,0,46,0,151,0,0,0,55,0,244,0,5,0,0,0,203,0,160,0,122,0,126,0,224,0,197,0,0,0,93,0,0,0,17,0,180,0,148,0,219,0,202,0,0,0,0,0,101,0,60,0,125,0,191,0,198,0,64,0,0,0,138,0,0,0,144,0,60,0,198,0,120,0,227,0,0,0,151,0,139,0,0,0,206,0,238,0,29,0,0,0,190,0,177,0,157,0,185,0,15,0,57,0,7,0,0,0,123,0,48,0,163,0,123,0,234,0,203,0,0,0,98,0,148,0,211,0,253,0,81,0,0,0,0,0,109,0,247,0,196,0,82,0,30,0,36,0,222,0,38,0,111,0,89,0,246,0,16,0,236,0,71,0,0,0,66,0,82,0,192,0,98,0,166,0,0,0,20,0,113,0,11,0,204,0,50,0,1,0,0,0,149,0,251,0,147,0,167,0,133,0,30,0,47,0,0,0,11,0,0,0,138,0,176,0,0,0,79,0,179,0,0,0,0,0,57,0,0,0,239,0,69,0,29,0,83,0,239,0,8,0,119,0,33,0,0,0,186,0,0,0,156,0,218,0,209,0,0,0,82,0,222,0,0,0,190,0,48,0,49,0,6,0,29,0,123,0,0,0,130,0,32,0,145,0,101,0,1,0,38,0,39,0,150,0,0,0,0,0,98,0,253,0,86,0,105,0,15,0,84,0,126,0,0,0,210,0,176,0,168,0,216,0,159,0,243,0,0,0,237,0,224,0,214,0,232,0,85,0,164,0,59,0,162,0,153,0,17,0,151,0,71,0,150,0,179,0,19,0,185,0,219,0,0,0,113,0,87,0,28,0,71,0,13,0,232,0,201,0,87,0,39,0,131,0,180,0,161,0,251,0,0,0,0,0,246,0,31,0,59,0,88,0,93,0,95,0,35,0,70,0,181,0,171,0,41,0,253,0,0,0,67,0,129,0,59,0,33,0,161,0,12,0,25,0,57,0,13,0,234,0,234,0,183,0,75,0,0,0,92,0,64,0,175,0,65,0,153,0,172,0,164,0,144,0,120,0,0,0,22,0,112,0,124,0,44,0,69,0,0,0,0,0,0,0,157,0,148,0,0,0,208,0,15,0,24,0,0,0,2,0,184,0,218,0,49,0,103,0,0,0,157,0,226,0,113,0,57,0,233,0,62,0,191,0,88,0,91,0,0,0,0,0,59,0,0,0,0,0,0,0,0,0,159,0,0,0,11,0,134,0,0,0,0,0,93,0,104,0,196,0,19,0,239,0,180,0,197,0,241,0,20,0,19,0,219,0,180,0,211,0,248,0,0,0,0,0,105,0,62,0,25,0,14,0,201,0,155,0,0,0,137,0,0,0,199,0,245,0,247,0,204,0,0,0,4,0,177,0,113,0,115,0,32,0,0,0,0,0,145,0,63,0,71,0,0,0,159,0,0,0,0,0,247,0,126,0,203,0,225,0,209,0,238,0,251,0,216,0,109,0,0,0,51,0,54,0,30,0,251,0,82,0,21,0,0,0,127,0,124,0,91,0,35,0,175,0,220,0,227,0,18,0,0,0,0,0,0,0,135,0,227,0,49,0,130,0,0,0,5,0,92,0,143,0,0,0,124,0,102,0,251,0,0,0,229,0,192,0,142,0,127,0,0,0,100,0,0,0,0,0,229,0,175,0,104,0,67,0,108,0,76,0,128,0,63,0,85,0,125,0,0,0,0,0,0,0,0,0,111,0,224,0,38,0,23,0,82,0,182,0,238,0,84,0,38,0,115,0,166,0,249,0,147,0,63,0,138,0,108,0,225,0,197,0,206,0,11,0,94,0,0,0,102,0,24,0,121,0,192,0,26,0,137,0,62,0,213,0,0,0,45,0,136,0,167,0,225,0,148,0,201,0,244,0,122,0,36,0,122,0,114,0,50,0,51,0,130,0,156,0,30,0,68,0,50,0,171,0,98,0,0,0,124,0,207,0,57,0,0,0,148,0,9,0,128,0,4,0,84,0,87,0,156,0,242,0,228,0,229,0,177,0,0,0,48,0,158,0,48,0,136,0,147,0,247,0,103,0,57,0,201,0,0,0,227,0,0,0,55,0,196,0,148,0,193,0,164,0,0,0,220,0,162,0,246,0,0,0,241,0,70,0,0,0,241,0,172,0,0,0,56,0,164,0,0,0,252,0,85,0,176,0,90,0,220,0,73,0,123,0,218,0,39,0,0,0,31,0,92,0,229,0,0,0,0,0,96,0);
signal scenario_full  : scenario_type := (24,31,138,31,9,31,33,31,130,31,167,31,66,31,8,31,8,30,37,31,62,31,62,30,230,31,68,31,50,31,71,31,130,31,10,31,45,31,118,31,118,30,98,31,38,31,224,31,59,31,59,30,180,31,180,30,180,29,180,28,115,31,88,31,88,30,103,31,255,31,21,31,21,30,94,31,94,30,89,31,89,30,5,31,3,31,3,30,3,29,206,31,215,31,156,31,156,30,158,31,127,31,189,31,99,31,99,30,82,31,82,30,43,31,46,31,196,31,182,31,74,31,29,31,29,30,38,31,150,31,137,31,137,30,89,31,60,31,60,30,60,29,79,31,241,31,181,31,170,31,243,31,164,31,129,31,115,31,169,31,169,30,55,31,238,31,191,31,13,31,13,30,214,31,44,31,44,30,104,31,167,31,168,31,228,31,172,31,185,31,185,30,74,31,74,30,240,31,159,31,159,30,159,29,163,31,43,31,10,31,10,30,250,31,162,31,162,30,115,31,255,31,67,31,156,31,235,31,219,31,219,30,57,31,142,31,16,31,160,31,129,31,129,30,129,29,129,28,30,31,30,30,215,31,140,31,223,31,136,31,192,31,171,31,15,31,28,31,62,31,80,31,91,31,91,30,242,31,136,31,6,31,138,31,120,31,223,31,22,31,114,31,137,31,137,30,137,29,118,31,118,30,47,31,225,31,253,31,216,31,92,31,168,31,9,31,53,31,191,31,237,31,237,30,138,31,182,31,214,31,196,31,79,31,150,31,178,31,252,31,36,31,243,31,229,31,253,31,19,31,60,31,60,30,96,31,96,30,135,31,135,30,135,29,96,31,88,31,88,30,167,31,25,31,61,31,101,31,101,30,28,31,53,31,234,31,171,31,64,31,173,31,29,31,43,31,150,31,42,31,42,30,109,31,109,30,128,31,158,31,217,31,120,31,120,30,184,31,182,31,29,31,81,31,81,30,81,29,130,31,167,31,210,31,164,31,94,31,236,31,167,31,49,31,230,31,167,31,167,30,130,31,130,30,11,31,104,31,249,31,115,31,63,31,80,31,45,31,111,31,77,31,96,31,96,30,160,31,183,31,133,31,146,31,178,31,54,31,42,31,42,30,188,31,255,31,223,31,230,31,203,31,203,30,203,29,168,31,151,31,175,31,172,31,65,31,14,31,68,31,74,31,105,31,202,31,112,31,63,31,234,31,234,30,234,29,159,31,150,31,213,31,208,31,43,31,159,31,118,31,118,30,221,31,187,31,187,30,235,31,227,31,75,31,75,30,75,29,75,28,135,31,70,31,115,31,115,30,172,31,166,31,166,30,58,31,58,30,58,29,58,28,214,31,93,31,93,30,247,31,240,31,188,31,188,30,85,31,67,31,135,31,43,31,43,30,141,31,50,31,247,31,247,30,247,29,117,31,117,30,117,29,141,31,7,31,7,30,69,31,132,31,171,31,183,31,214,31,214,30,153,31,130,31,39,31,254,31,254,30,164,31,109,31,215,31,98,31,64,31,33,31,255,31,27,31,27,30,27,29,112,31,12,31,29,31,122,31,122,30,93,31,179,31,101,31,137,31,210,31,47,31,47,30,131,31,101,31,72,31,228,31,106,31,203,31,203,30,59,31,149,31,196,31,49,31,111,31,159,31,192,31,192,30,255,31,29,31,105,31,58,31,25,31,67,31,23,31,46,31,132,31,205,31,205,30,159,31,220,31,190,31,166,31,68,31,20,31,160,31,155,31,250,31,106,31,152,31,152,30,149,31,241,31,207,31,147,31,70,31,78,31,29,31,159,31,159,30,159,29,141,31,10,31,127,31,86,31,80,31,23,31,23,30,10,31,10,30,200,31,61,31,61,30,61,29,248,31,25,31,182,31,182,30,198,31,198,30,225,31,249,31,29,31,151,31,252,31,187,31,9,31,178,31,174,31,248,31,223,31,82,31,12,31,157,31,13,31,232,31,140,31,125,31,17,31,252,31,104,31,71,31,40,31,160,31,10,31,59,31,133,31,159,31,159,30,168,31,59,31,150,31,43,31,70,31,70,30,46,31,151,31,151,30,55,31,244,31,5,31,5,30,203,31,160,31,122,31,126,31,224,31,197,31,197,30,93,31,93,30,17,31,180,31,148,31,219,31,202,31,202,30,202,29,101,31,60,31,125,31,191,31,198,31,64,31,64,30,138,31,138,30,144,31,60,31,198,31,120,31,227,31,227,30,151,31,139,31,139,30,206,31,238,31,29,31,29,30,190,31,177,31,157,31,185,31,15,31,57,31,7,31,7,30,123,31,48,31,163,31,123,31,234,31,203,31,203,30,98,31,148,31,211,31,253,31,81,31,81,30,81,29,109,31,247,31,196,31,82,31,30,31,36,31,222,31,38,31,111,31,89,31,246,31,16,31,236,31,71,31,71,30,66,31,82,31,192,31,98,31,166,31,166,30,20,31,113,31,11,31,204,31,50,31,1,31,1,30,149,31,251,31,147,31,167,31,133,31,30,31,47,31,47,30,11,31,11,30,138,31,176,31,176,30,79,31,179,31,179,30,179,29,57,31,57,30,239,31,69,31,29,31,83,31,239,31,8,31,119,31,33,31,33,30,186,31,186,30,156,31,218,31,209,31,209,30,82,31,222,31,222,30,190,31,48,31,49,31,6,31,29,31,123,31,123,30,130,31,32,31,145,31,101,31,1,31,38,31,39,31,150,31,150,30,150,29,98,31,253,31,86,31,105,31,15,31,84,31,126,31,126,30,210,31,176,31,168,31,216,31,159,31,243,31,243,30,237,31,224,31,214,31,232,31,85,31,164,31,59,31,162,31,153,31,17,31,151,31,71,31,150,31,179,31,19,31,185,31,219,31,219,30,113,31,87,31,28,31,71,31,13,31,232,31,201,31,87,31,39,31,131,31,180,31,161,31,251,31,251,30,251,29,246,31,31,31,59,31,88,31,93,31,95,31,35,31,70,31,181,31,171,31,41,31,253,31,253,30,67,31,129,31,59,31,33,31,161,31,12,31,25,31,57,31,13,31,234,31,234,31,183,31,75,31,75,30,92,31,64,31,175,31,65,31,153,31,172,31,164,31,144,31,120,31,120,30,22,31,112,31,124,31,44,31,69,31,69,30,69,29,69,28,157,31,148,31,148,30,208,31,15,31,24,31,24,30,2,31,184,31,218,31,49,31,103,31,103,30,157,31,226,31,113,31,57,31,233,31,62,31,191,31,88,31,91,31,91,30,91,29,59,31,59,30,59,29,59,28,59,27,159,31,159,30,11,31,134,31,134,30,134,29,93,31,104,31,196,31,19,31,239,31,180,31,197,31,241,31,20,31,19,31,219,31,180,31,211,31,248,31,248,30,248,29,105,31,62,31,25,31,14,31,201,31,155,31,155,30,137,31,137,30,199,31,245,31,247,31,204,31,204,30,4,31,177,31,113,31,115,31,32,31,32,30,32,29,145,31,63,31,71,31,71,30,159,31,159,30,159,29,247,31,126,31,203,31,225,31,209,31,238,31,251,31,216,31,109,31,109,30,51,31,54,31,30,31,251,31,82,31,21,31,21,30,127,31,124,31,91,31,35,31,175,31,220,31,227,31,18,31,18,30,18,29,18,28,135,31,227,31,49,31,130,31,130,30,5,31,92,31,143,31,143,30,124,31,102,31,251,31,251,30,229,31,192,31,142,31,127,31,127,30,100,31,100,30,100,29,229,31,175,31,104,31,67,31,108,31,76,31,128,31,63,31,85,31,125,31,125,30,125,29,125,28,125,27,111,31,224,31,38,31,23,31,82,31,182,31,238,31,84,31,38,31,115,31,166,31,249,31,147,31,63,31,138,31,108,31,225,31,197,31,206,31,11,31,94,31,94,30,102,31,24,31,121,31,192,31,26,31,137,31,62,31,213,31,213,30,45,31,136,31,167,31,225,31,148,31,201,31,244,31,122,31,36,31,122,31,114,31,50,31,51,31,130,31,156,31,30,31,68,31,50,31,171,31,98,31,98,30,124,31,207,31,57,31,57,30,148,31,9,31,128,31,4,31,84,31,87,31,156,31,242,31,228,31,229,31,177,31,177,30,48,31,158,31,48,31,136,31,147,31,247,31,103,31,57,31,201,31,201,30,227,31,227,30,55,31,196,31,148,31,193,31,164,31,164,30,220,31,162,31,246,31,246,30,241,31,70,31,70,30,241,31,172,31,172,30,56,31,164,31,164,30,252,31,85,31,176,31,90,31,220,31,73,31,123,31,218,31,39,31,39,30,31,31,92,31,229,31,229,30,229,29,96,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
