-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_958 is
end project_tb_958;

architecture project_tb_arch_958 of project_tb_958 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 813;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (252,0,0,0,45,0,96,0,166,0,0,0,0,0,88,0,0,0,25,0,201,0,230,0,0,0,59,0,100,0,0,0,193,0,3,0,0,0,149,0,207,0,243,0,0,0,0,0,236,0,122,0,102,0,33,0,180,0,92,0,2,0,101,0,195,0,231,0,137,0,73,0,213,0,131,0,218,0,0,0,175,0,138,0,110,0,146,0,218,0,0,0,251,0,127,0,0,0,43,0,109,0,131,0,99,0,0,0,128,0,97,0,152,0,60,0,56,0,106,0,242,0,96,0,92,0,192,0,139,0,74,0,0,0,187,0,60,0,197,0,9,0,133,0,149,0,82,0,255,0,190,0,181,0,236,0,0,0,87,0,0,0,30,0,210,0,146,0,116,0,0,0,31,0,0,0,247,0,0,0,0,0,57,0,26,0,78,0,155,0,53,0,65,0,73,0,152,0,53,0,91,0,0,0,113,0,7,0,94,0,232,0,0,0,8,0,55,0,0,0,43,0,86,0,2,0,111,0,217,0,0,0,131,0,197,0,190,0,197,0,168,0,182,0,0,0,213,0,180,0,80,0,184,0,172,0,205,0,157,0,50,0,212,0,0,0,246,0,152,0,106,0,83,0,243,0,29,0,77,0,14,0,0,0,75,0,62,0,54,0,119,0,30,0,90,0,146,0,51,0,188,0,157,0,158,0,54,0,170,0,161,0,20,0,173,0,0,0,160,0,0,0,55,0,9,0,45,0,84,0,106,0,0,0,49,0,184,0,36,0,231,0,77,0,139,0,0,0,74,0,176,0,149,0,0,0,235,0,129,0,253,0,83,0,205,0,22,0,160,0,0,0,0,0,231,0,113,0,249,0,249,0,169,0,113,0,176,0,212,0,234,0,237,0,0,0,255,0,223,0,55,0,222,0,101,0,49,0,0,0,251,0,53,0,0,0,0,0,183,0,244,0,11,0,0,0,98,0,0,0,251,0,0,0,155,0,200,0,0,0,216,0,99,0,92,0,1,0,0,0,80,0,44,0,74,0,8,0,7,0,69,0,182,0,40,0,81,0,105,0,217,0,70,0,49,0,0,0,10,0,0,0,154,0,254,0,186,0,234,0,175,0,0,0,28,0,173,0,63,0,0,0,0,0,0,0,212,0,7,0,118,0,217,0,205,0,0,0,10,0,4,0,207,0,0,0,2,0,148,0,131,0,25,0,0,0,0,0,87,0,116,0,242,0,149,0,57,0,65,0,74,0,120,0,223,0,116,0,239,0,101,0,0,0,0,0,0,0,138,0,78,0,122,0,114,0,0,0,114,0,0,0,165,0,219,0,17,0,142,0,249,0,96,0,139,0,74,0,102,0,108,0,183,0,255,0,187,0,126,0,0,0,108,0,74,0,232,0,0,0,132,0,0,0,181,0,62,0,80,0,0,0,157,0,229,0,142,0,141,0,0,0,0,0,0,0,159,0,51,0,0,0,5,0,134,0,220,0,135,0,162,0,4,0,121,0,249,0,91,0,0,0,235,0,38,0,184,0,0,0,184,0,137,0,230,0,111,0,166,0,123,0,0,0,0,0,163,0,167,0,91,0,134,0,171,0,0,0,254,0,148,0,70,0,0,0,0,0,0,0,160,0,198,0,237,0,124,0,117,0,0,0,0,0,197,0,35,0,0,0,183,0,220,0,144,0,141,0,0,0,188,0,35,0,140,0,153,0,200,0,133,0,119,0,132,0,236,0,19,0,51,0,196,0,0,0,8,0,89,0,83,0,7,0,4,0,227,0,0,0,0,0,188,0,152,0,37,0,132,0,152,0,242,0,0,0,0,0,111,0,226,0,163,0,0,0,181,0,238,0,0,0,104,0,76,0,152,0,39,0,139,0,54,0,203,0,174,0,100,0,85,0,16,0,73,0,67,0,49,0,212,0,68,0,8,0,0,0,235,0,71,0,41,0,23,0,224,0,136,0,59,0,1,0,47,0,105,0,249,0,230,0,246,0,163,0,179,0,151,0,192,0,224,0,53,0,222,0,78,0,34,0,59,0,254,0,5,0,27,0,0,0,59,0,0,0,239,0,0,0,42,0,34,0,53,0,78,0,39,0,13,0,100,0,42,0,128,0,30,0,115,0,76,0,151,0,200,0,29,0,0,0,0,0,168,0,232,0,0,0,0,0,58,0,81,0,251,0,116,0,246,0,68,0,167,0,40,0,114,0,243,0,26,0,0,0,71,0,133,0,128,0,18,0,79,0,52,0,30,0,88,0,238,0,147,0,0,0,6,0,54,0,246,0,0,0,151,0,131,0,78,0,245,0,66,0,130,0,0,0,206,0,0,0,69,0,60,0,187,0,87,0,82,0,0,0,238,0,236,0,101,0,228,0,0,0,77,0,245,0,158,0,75,0,6,0,0,0,195,0,233,0,0,0,0,0,88,0,0,0,109,0,30,0,9,0,223,0,181,0,44,0,2,0,0,0,0,0,54,0,0,0,247,0,149,0,85,0,0,0,110,0,113,0,55,0,9,0,235,0,218,0,190,0,119,0,213,0,203,0,30,0,47,0,47,0,78,0,127,0,30,0,72,0,235,0,46,0,184,0,252,0,67,0,147,0,0,0,156,0,253,0,1,0,21,0,0,0,103,0,88,0,0,0,24,0,0,0,29,0,0,0,239,0,0,0,0,0,66,0,31,0,139,0,34,0,0,0,199,0,101,0,214,0,78,0,64,0,237,0,255,0,232,0,0,0,152,0,228,0,0,0,141,0,166,0,161,0,46,0,27,0,198,0,63,0,133,0,99,0,77,0,238,0,108,0,110,0,230,0,0,0,28,0,2,0,101,0,0,0,0,0,242,0,90,0,113,0,0,0,225,0,10,0,239,0,104,0,210,0,118,0,244,0,0,0,204,0,0,0,161,0,7,0,91,0,11,0,88,0,104,0,155,0,164,0,240,0,80,0,12,0,149,0,204,0,179,0,64,0,188,0,227,0,13,0,0,0,191,0,206,0,207,0,211,0,0,0,242,0,194,0,28,0,0,0,222,0,0,0,207,0,74,0,21,0,109,0,76,0,109,0,93,0,145,0,139,0,77,0,51,0,180,0,55,0,45,0,9,0,0,0,0,0,114,0,93,0,0,0,161,0,2,0,195,0,11,0,117,0,0,0,164,0,201,0,183,0,124,0,215,0,132,0,17,0,0,0,146,0,0,0,130,0,61,0,60,0,233,0,15,0,143,0,66,0,106,0,167,0,41,0,248,0,23,0,143,0,244,0,127,0,86,0,89,0,54,0,167,0,85,0,17,0,85,0,205,0,56,0,70,0,224,0,53,0,118,0,92,0,171,0,70,0,177,0,10,0,233,0,0,0,0,0,140,0,121,0,159,0,52,0,52,0,179,0,244,0,44,0,80,0,187,0,162,0,223,0,0,0,243,0,120,0,150,0,109,0,144,0,0,0,0,0,202,0,245,0,212,0,186,0,0,0,104,0,144,0,212,0,18,0,0,0,64,0,93,0,0,0,119,0,206,0,6,0,115,0,135,0,0,0,188,0,146,0,253,0,61,0,14,0,71,0,93,0,0,0,33,0,0,0,127,0,0,0,111,0,65,0,0,0,171,0,0,0,253,0,168,0,105,0,192,0,7,0,0,0,187,0,224,0,89,0,97,0);
signal scenario_full  : scenario_type := (252,31,252,30,45,31,96,31,166,31,166,30,166,29,88,31,88,30,25,31,201,31,230,31,230,30,59,31,100,31,100,30,193,31,3,31,3,30,149,31,207,31,243,31,243,30,243,29,236,31,122,31,102,31,33,31,180,31,92,31,2,31,101,31,195,31,231,31,137,31,73,31,213,31,131,31,218,31,218,30,175,31,138,31,110,31,146,31,218,31,218,30,251,31,127,31,127,30,43,31,109,31,131,31,99,31,99,30,128,31,97,31,152,31,60,31,56,31,106,31,242,31,96,31,92,31,192,31,139,31,74,31,74,30,187,31,60,31,197,31,9,31,133,31,149,31,82,31,255,31,190,31,181,31,236,31,236,30,87,31,87,30,30,31,210,31,146,31,116,31,116,30,31,31,31,30,247,31,247,30,247,29,57,31,26,31,78,31,155,31,53,31,65,31,73,31,152,31,53,31,91,31,91,30,113,31,7,31,94,31,232,31,232,30,8,31,55,31,55,30,43,31,86,31,2,31,111,31,217,31,217,30,131,31,197,31,190,31,197,31,168,31,182,31,182,30,213,31,180,31,80,31,184,31,172,31,205,31,157,31,50,31,212,31,212,30,246,31,152,31,106,31,83,31,243,31,29,31,77,31,14,31,14,30,75,31,62,31,54,31,119,31,30,31,90,31,146,31,51,31,188,31,157,31,158,31,54,31,170,31,161,31,20,31,173,31,173,30,160,31,160,30,55,31,9,31,45,31,84,31,106,31,106,30,49,31,184,31,36,31,231,31,77,31,139,31,139,30,74,31,176,31,149,31,149,30,235,31,129,31,253,31,83,31,205,31,22,31,160,31,160,30,160,29,231,31,113,31,249,31,249,31,169,31,113,31,176,31,212,31,234,31,237,31,237,30,255,31,223,31,55,31,222,31,101,31,49,31,49,30,251,31,53,31,53,30,53,29,183,31,244,31,11,31,11,30,98,31,98,30,251,31,251,30,155,31,200,31,200,30,216,31,99,31,92,31,1,31,1,30,80,31,44,31,74,31,8,31,7,31,69,31,182,31,40,31,81,31,105,31,217,31,70,31,49,31,49,30,10,31,10,30,154,31,254,31,186,31,234,31,175,31,175,30,28,31,173,31,63,31,63,30,63,29,63,28,212,31,7,31,118,31,217,31,205,31,205,30,10,31,4,31,207,31,207,30,2,31,148,31,131,31,25,31,25,30,25,29,87,31,116,31,242,31,149,31,57,31,65,31,74,31,120,31,223,31,116,31,239,31,101,31,101,30,101,29,101,28,138,31,78,31,122,31,114,31,114,30,114,31,114,30,165,31,219,31,17,31,142,31,249,31,96,31,139,31,74,31,102,31,108,31,183,31,255,31,187,31,126,31,126,30,108,31,74,31,232,31,232,30,132,31,132,30,181,31,62,31,80,31,80,30,157,31,229,31,142,31,141,31,141,30,141,29,141,28,159,31,51,31,51,30,5,31,134,31,220,31,135,31,162,31,4,31,121,31,249,31,91,31,91,30,235,31,38,31,184,31,184,30,184,31,137,31,230,31,111,31,166,31,123,31,123,30,123,29,163,31,167,31,91,31,134,31,171,31,171,30,254,31,148,31,70,31,70,30,70,29,70,28,160,31,198,31,237,31,124,31,117,31,117,30,117,29,197,31,35,31,35,30,183,31,220,31,144,31,141,31,141,30,188,31,35,31,140,31,153,31,200,31,133,31,119,31,132,31,236,31,19,31,51,31,196,31,196,30,8,31,89,31,83,31,7,31,4,31,227,31,227,30,227,29,188,31,152,31,37,31,132,31,152,31,242,31,242,30,242,29,111,31,226,31,163,31,163,30,181,31,238,31,238,30,104,31,76,31,152,31,39,31,139,31,54,31,203,31,174,31,100,31,85,31,16,31,73,31,67,31,49,31,212,31,68,31,8,31,8,30,235,31,71,31,41,31,23,31,224,31,136,31,59,31,1,31,47,31,105,31,249,31,230,31,246,31,163,31,179,31,151,31,192,31,224,31,53,31,222,31,78,31,34,31,59,31,254,31,5,31,27,31,27,30,59,31,59,30,239,31,239,30,42,31,34,31,53,31,78,31,39,31,13,31,100,31,42,31,128,31,30,31,115,31,76,31,151,31,200,31,29,31,29,30,29,29,168,31,232,31,232,30,232,29,58,31,81,31,251,31,116,31,246,31,68,31,167,31,40,31,114,31,243,31,26,31,26,30,71,31,133,31,128,31,18,31,79,31,52,31,30,31,88,31,238,31,147,31,147,30,6,31,54,31,246,31,246,30,151,31,131,31,78,31,245,31,66,31,130,31,130,30,206,31,206,30,69,31,60,31,187,31,87,31,82,31,82,30,238,31,236,31,101,31,228,31,228,30,77,31,245,31,158,31,75,31,6,31,6,30,195,31,233,31,233,30,233,29,88,31,88,30,109,31,30,31,9,31,223,31,181,31,44,31,2,31,2,30,2,29,54,31,54,30,247,31,149,31,85,31,85,30,110,31,113,31,55,31,9,31,235,31,218,31,190,31,119,31,213,31,203,31,30,31,47,31,47,31,78,31,127,31,30,31,72,31,235,31,46,31,184,31,252,31,67,31,147,31,147,30,156,31,253,31,1,31,21,31,21,30,103,31,88,31,88,30,24,31,24,30,29,31,29,30,239,31,239,30,239,29,66,31,31,31,139,31,34,31,34,30,199,31,101,31,214,31,78,31,64,31,237,31,255,31,232,31,232,30,152,31,228,31,228,30,141,31,166,31,161,31,46,31,27,31,198,31,63,31,133,31,99,31,77,31,238,31,108,31,110,31,230,31,230,30,28,31,2,31,101,31,101,30,101,29,242,31,90,31,113,31,113,30,225,31,10,31,239,31,104,31,210,31,118,31,244,31,244,30,204,31,204,30,161,31,7,31,91,31,11,31,88,31,104,31,155,31,164,31,240,31,80,31,12,31,149,31,204,31,179,31,64,31,188,31,227,31,13,31,13,30,191,31,206,31,207,31,211,31,211,30,242,31,194,31,28,31,28,30,222,31,222,30,207,31,74,31,21,31,109,31,76,31,109,31,93,31,145,31,139,31,77,31,51,31,180,31,55,31,45,31,9,31,9,30,9,29,114,31,93,31,93,30,161,31,2,31,195,31,11,31,117,31,117,30,164,31,201,31,183,31,124,31,215,31,132,31,17,31,17,30,146,31,146,30,130,31,61,31,60,31,233,31,15,31,143,31,66,31,106,31,167,31,41,31,248,31,23,31,143,31,244,31,127,31,86,31,89,31,54,31,167,31,85,31,17,31,85,31,205,31,56,31,70,31,224,31,53,31,118,31,92,31,171,31,70,31,177,31,10,31,233,31,233,30,233,29,140,31,121,31,159,31,52,31,52,31,179,31,244,31,44,31,80,31,187,31,162,31,223,31,223,30,243,31,120,31,150,31,109,31,144,31,144,30,144,29,202,31,245,31,212,31,186,31,186,30,104,31,144,31,212,31,18,31,18,30,64,31,93,31,93,30,119,31,206,31,6,31,115,31,135,31,135,30,188,31,146,31,253,31,61,31,14,31,71,31,93,31,93,30,33,31,33,30,127,31,127,30,111,31,65,31,65,30,171,31,171,30,253,31,168,31,105,31,192,31,7,31,7,30,187,31,224,31,89,31,97,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
