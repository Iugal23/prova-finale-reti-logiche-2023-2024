-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 689;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (197,0,244,0,58,0,66,0,184,0,45,0,84,0,172,0,86,0,166,0,250,0,108,0,0,0,69,0,220,0,0,0,4,0,0,0,136,0,203,0,160,0,161,0,0,0,0,0,216,0,0,0,192,0,0,0,16,0,13,0,166,0,47,0,0,0,0,0,0,0,254,0,32,0,65,0,77,0,68,0,216,0,67,0,165,0,150,0,3,0,84,0,40,0,37,0,171,0,24,0,211,0,164,0,174,0,69,0,234,0,90,0,153,0,115,0,18,0,165,0,0,0,83,0,34,0,0,0,234,0,206,0,114,0,94,0,189,0,17,0,60,0,62,0,0,0,203,0,124,0,150,0,184,0,0,0,91,0,149,0,59,0,51,0,0,0,176,0,183,0,147,0,220,0,68,0,0,0,5,0,253,0,247,0,118,0,253,0,240,0,66,0,179,0,197,0,128,0,0,0,141,0,77,0,18,0,157,0,206,0,0,0,11,0,78,0,112,0,47,0,115,0,0,0,18,0,49,0,9,0,108,0,20,0,122,0,123,0,222,0,0,0,30,0,209,0,18,0,13,0,11,0,0,0,120,0,0,0,0,0,6,0,228,0,232,0,0,0,203,0,10,0,0,0,93,0,99,0,57,0,221,0,91,0,0,0,135,0,171,0,27,0,0,0,0,0,151,0,63,0,0,0,169,0,104,0,100,0,112,0,56,0,125,0,252,0,120,0,134,0,48,0,0,0,0,0,185,0,9,0,0,0,0,0,131,0,0,0,3,0,0,0,57,0,76,0,50,0,43,0,241,0,252,0,0,0,34,0,214,0,194,0,230,0,64,0,0,0,81,0,43,0,219,0,73,0,0,0,93,0,0,0,124,0,24,0,73,0,198,0,199,0,89,0,156,0,81,0,155,0,62,0,140,0,0,0,0,0,241,0,48,0,183,0,234,0,0,0,212,0,251,0,0,0,0,0,124,0,0,0,86,0,100,0,0,0,187,0,218,0,0,0,0,0,148,0,244,0,68,0,147,0,26,0,227,0,226,0,49,0,114,0,67,0,11,0,245,0,214,0,203,0,81,0,239,0,12,0,0,0,48,0,139,0,0,0,168,0,39,0,20,0,0,0,157,0,165,0,0,0,129,0,0,0,99,0,173,0,46,0,0,0,99,0,63,0,142,0,25,0,82,0,126,0,216,0,82,0,37,0,0,0,0,0,57,0,203,0,0,0,0,0,62,0,72,0,60,0,137,0,231,0,18,0,247,0,220,0,213,0,103,0,3,0,56,0,0,0,84,0,246,0,59,0,0,0,65,0,132,0,161,0,91,0,65,0,178,0,73,0,143,0,0,0,23,0,181,0,170,0,55,0,29,0,148,0,172,0,134,0,84,0,44,0,78,0,18,0,96,0,181,0,0,0,0,0,163,0,0,0,0,0,189,0,246,0,70,0,24,0,0,0,163,0,129,0,0,0,0,0,245,0,0,0,126,0,57,0,83,0,178,0,65,0,201,0,26,0,210,0,165,0,37,0,174,0,109,0,0,0,103,0,120,0,106,0,168,0,149,0,31,0,76,0,233,0,7,0,211,0,219,0,59,0,149,0,0,0,59,0,198,0,176,0,0,0,218,0,199,0,0,0,97,0,85,0,63,0,139,0,211,0,0,0,0,0,25,0,159,0,45,0,95,0,16,0,39,0,235,0,88,0,214,0,190,0,225,0,37,0,0,0,25,0,0,0,215,0,0,0,66,0,194,0,116,0,46,0,0,0,0,0,103,0,0,0,246,0,1,0,228,0,170,0,0,0,228,0,0,0,158,0,1,0,0,0,67,0,153,0,196,0,68,0,116,0,52,0,0,0,230,0,24,0,247,0,78,0,152,0,14,0,180,0,220,0,112,0,187,0,0,0,209,0,236,0,33,0,0,0,163,0,43,0,118,0,192,0,23,0,198,0,0,0,42,0,242,0,0,0,146,0,0,0,164,0,122,0,41,0,15,0,35,0,206,0,45,0,149,0,196,0,144,0,0,0,27,0,132,0,52,0,141,0,0,0,132,0,0,0,0,0,42,0,51,0,94,0,163,0,245,0,32,0,125,0,147,0,0,0,244,0,139,0,118,0,127,0,241,0,221,0,165,0,73,0,0,0,50,0,139,0,35,0,182,0,80,0,243,0,203,0,125,0,226,0,28,0,0,0,0,0,205,0,227,0,151,0,11,0,133,0,205,0,107,0,0,0,51,0,0,0,0,0,184,0,5,0,108,0,35,0,101,0,97,0,229,0,0,0,195,0,57,0,194,0,29,0,24,0,0,0,133,0,102,0,35,0,252,0,225,0,61,0,244,0,152,0,211,0,221,0,20,0,7,0,253,0,145,0,151,0,53,0,5,0,69,0,66,0,0,0,211,0,193,0,82,0,10,0,199,0,166,0,48,0,0,0,0,0,30,0,41,0,0,0,136,0,0,0,18,0,61,0,0,0,173,0,0,0,0,0,86,0,74,0,149,0,127,0,13,0,0,0,22,0,0,0,133,0,0,0,169,0,7,0,0,0,0,0,75,0,63,0,77,0,186,0,0,0,0,0,237,0,236,0,42,0,40,0,201,0,73,0,151,0,0,0,17,0,126,0,167,0,156,0,41,0,230,0,185,0,79,0,0,0,21,0,121,0,235,0,130,0,160,0,183,0,250,0,92,0,224,0,200,0,53,0,84,0,0,0,28,0,0,0,212,0,35,0,18,0,196,0,147,0,100,0,217,0,46,0,67,0,150,0,20,0,0,0,88,0,66,0,8,0,0,0,28,0,180,0,80,0,0,0,182,0,0,0,87,0,0,0,212,0,35,0,0,0,249,0,87,0,127,0,155,0,0,0,75,0,69,0,145,0,72,0,0,0,58,0,87,0,42,0,0,0,236,0,146,0,177,0,204,0,0,0,39,0,23,0,69,0,228,0,0,0,43,0,0,0,163,0,210,0,122,0,0,0,33,0,172,0,0,0,68,0,49,0,181,0,52,0,178,0,183,0,0,0,0,0,244,0,255,0,136,0,7,0,242,0,0,0,0,0,0,0,75,0,147,0,231,0,66,0,222,0,92,0,76,0,0,0,21,0,0,0);
signal scenario_full  : scenario_type := (197,31,244,31,58,31,66,31,184,31,45,31,84,31,172,31,86,31,166,31,250,31,108,31,108,30,69,31,220,31,220,30,4,31,4,30,136,31,203,31,160,31,161,31,161,30,161,29,216,31,216,30,192,31,192,30,16,31,13,31,166,31,47,31,47,30,47,29,47,28,254,31,32,31,65,31,77,31,68,31,216,31,67,31,165,31,150,31,3,31,84,31,40,31,37,31,171,31,24,31,211,31,164,31,174,31,69,31,234,31,90,31,153,31,115,31,18,31,165,31,165,30,83,31,34,31,34,30,234,31,206,31,114,31,94,31,189,31,17,31,60,31,62,31,62,30,203,31,124,31,150,31,184,31,184,30,91,31,149,31,59,31,51,31,51,30,176,31,183,31,147,31,220,31,68,31,68,30,5,31,253,31,247,31,118,31,253,31,240,31,66,31,179,31,197,31,128,31,128,30,141,31,77,31,18,31,157,31,206,31,206,30,11,31,78,31,112,31,47,31,115,31,115,30,18,31,49,31,9,31,108,31,20,31,122,31,123,31,222,31,222,30,30,31,209,31,18,31,13,31,11,31,11,30,120,31,120,30,120,29,6,31,228,31,232,31,232,30,203,31,10,31,10,30,93,31,99,31,57,31,221,31,91,31,91,30,135,31,171,31,27,31,27,30,27,29,151,31,63,31,63,30,169,31,104,31,100,31,112,31,56,31,125,31,252,31,120,31,134,31,48,31,48,30,48,29,185,31,9,31,9,30,9,29,131,31,131,30,3,31,3,30,57,31,76,31,50,31,43,31,241,31,252,31,252,30,34,31,214,31,194,31,230,31,64,31,64,30,81,31,43,31,219,31,73,31,73,30,93,31,93,30,124,31,24,31,73,31,198,31,199,31,89,31,156,31,81,31,155,31,62,31,140,31,140,30,140,29,241,31,48,31,183,31,234,31,234,30,212,31,251,31,251,30,251,29,124,31,124,30,86,31,100,31,100,30,187,31,218,31,218,30,218,29,148,31,244,31,68,31,147,31,26,31,227,31,226,31,49,31,114,31,67,31,11,31,245,31,214,31,203,31,81,31,239,31,12,31,12,30,48,31,139,31,139,30,168,31,39,31,20,31,20,30,157,31,165,31,165,30,129,31,129,30,99,31,173,31,46,31,46,30,99,31,63,31,142,31,25,31,82,31,126,31,216,31,82,31,37,31,37,30,37,29,57,31,203,31,203,30,203,29,62,31,72,31,60,31,137,31,231,31,18,31,247,31,220,31,213,31,103,31,3,31,56,31,56,30,84,31,246,31,59,31,59,30,65,31,132,31,161,31,91,31,65,31,178,31,73,31,143,31,143,30,23,31,181,31,170,31,55,31,29,31,148,31,172,31,134,31,84,31,44,31,78,31,18,31,96,31,181,31,181,30,181,29,163,31,163,30,163,29,189,31,246,31,70,31,24,31,24,30,163,31,129,31,129,30,129,29,245,31,245,30,126,31,57,31,83,31,178,31,65,31,201,31,26,31,210,31,165,31,37,31,174,31,109,31,109,30,103,31,120,31,106,31,168,31,149,31,31,31,76,31,233,31,7,31,211,31,219,31,59,31,149,31,149,30,59,31,198,31,176,31,176,30,218,31,199,31,199,30,97,31,85,31,63,31,139,31,211,31,211,30,211,29,25,31,159,31,45,31,95,31,16,31,39,31,235,31,88,31,214,31,190,31,225,31,37,31,37,30,25,31,25,30,215,31,215,30,66,31,194,31,116,31,46,31,46,30,46,29,103,31,103,30,246,31,1,31,228,31,170,31,170,30,228,31,228,30,158,31,1,31,1,30,67,31,153,31,196,31,68,31,116,31,52,31,52,30,230,31,24,31,247,31,78,31,152,31,14,31,180,31,220,31,112,31,187,31,187,30,209,31,236,31,33,31,33,30,163,31,43,31,118,31,192,31,23,31,198,31,198,30,42,31,242,31,242,30,146,31,146,30,164,31,122,31,41,31,15,31,35,31,206,31,45,31,149,31,196,31,144,31,144,30,27,31,132,31,52,31,141,31,141,30,132,31,132,30,132,29,42,31,51,31,94,31,163,31,245,31,32,31,125,31,147,31,147,30,244,31,139,31,118,31,127,31,241,31,221,31,165,31,73,31,73,30,50,31,139,31,35,31,182,31,80,31,243,31,203,31,125,31,226,31,28,31,28,30,28,29,205,31,227,31,151,31,11,31,133,31,205,31,107,31,107,30,51,31,51,30,51,29,184,31,5,31,108,31,35,31,101,31,97,31,229,31,229,30,195,31,57,31,194,31,29,31,24,31,24,30,133,31,102,31,35,31,252,31,225,31,61,31,244,31,152,31,211,31,221,31,20,31,7,31,253,31,145,31,151,31,53,31,5,31,69,31,66,31,66,30,211,31,193,31,82,31,10,31,199,31,166,31,48,31,48,30,48,29,30,31,41,31,41,30,136,31,136,30,18,31,61,31,61,30,173,31,173,30,173,29,86,31,74,31,149,31,127,31,13,31,13,30,22,31,22,30,133,31,133,30,169,31,7,31,7,30,7,29,75,31,63,31,77,31,186,31,186,30,186,29,237,31,236,31,42,31,40,31,201,31,73,31,151,31,151,30,17,31,126,31,167,31,156,31,41,31,230,31,185,31,79,31,79,30,21,31,121,31,235,31,130,31,160,31,183,31,250,31,92,31,224,31,200,31,53,31,84,31,84,30,28,31,28,30,212,31,35,31,18,31,196,31,147,31,100,31,217,31,46,31,67,31,150,31,20,31,20,30,88,31,66,31,8,31,8,30,28,31,180,31,80,31,80,30,182,31,182,30,87,31,87,30,212,31,35,31,35,30,249,31,87,31,127,31,155,31,155,30,75,31,69,31,145,31,72,31,72,30,58,31,87,31,42,31,42,30,236,31,146,31,177,31,204,31,204,30,39,31,23,31,69,31,228,31,228,30,43,31,43,30,163,31,210,31,122,31,122,30,33,31,172,31,172,30,68,31,49,31,181,31,52,31,178,31,183,31,183,30,183,29,244,31,255,31,136,31,7,31,242,31,242,30,242,29,242,28,75,31,147,31,231,31,66,31,222,31,92,31,76,31,76,30,21,31,21,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
