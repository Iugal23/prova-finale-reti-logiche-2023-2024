-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_930 is
end project_tb_930;

architecture project_tb_arch_930 of project_tb_930 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 171;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (34,0,192,0,0,0,221,0,0,0,141,0,0,0,253,0,186,0,0,0,93,0,68,0,42,0,25,0,0,0,25,0,0,0,165,0,0,0,0,0,0,0,0,0,163,0,62,0,104,0,248,0,152,0,4,0,7,0,46,0,164,0,236,0,152,0,21,0,76,0,92,0,25,0,224,0,220,0,0,0,5,0,164,0,120,0,87,0,0,0,108,0,0,0,0,0,127,0,17,0,0,0,0,0,0,0,0,0,208,0,163,0,78,0,133,0,194,0,8,0,28,0,0,0,0,0,230,0,197,0,0,0,11,0,3,0,200,0,0,0,162,0,218,0,212,0,90,0,0,0,109,0,24,0,0,0,174,0,0,0,26,0,107,0,83,0,29,0,37,0,79,0,224,0,78,0,0,0,83,0,22,0,52,0,186,0,157,0,44,0,144,0,246,0,0,0,62,0,216,0,221,0,164,0,0,0,99,0,147,0,139,0,74,0,197,0,138,0,176,0,244,0,185,0,188,0,14,0,139,0,0,0,120,0,33,0,194,0,177,0,140,0,95,0,87,0,149,0,25,0,176,0,0,0,76,0,46,0,115,0,107,0,2,0,23,0,139,0,0,0,104,0,189,0,252,0,0,0,12,0,127,0,248,0,88,0,118,0,150,0,228,0,104,0,0,0,216,0,89,0,189,0,194,0,239,0,120,0,0,0,0,0,217,0,0,0,78,0,198,0,0,0,20,0,239,0,48,0,0,0,63,0,105,0,207,0,0,0,88,0,169,0);
signal scenario_full  : scenario_type := (34,31,192,31,192,30,221,31,221,30,141,31,141,30,253,31,186,31,186,30,93,31,68,31,42,31,25,31,25,30,25,31,25,30,165,31,165,30,165,29,165,28,165,27,163,31,62,31,104,31,248,31,152,31,4,31,7,31,46,31,164,31,236,31,152,31,21,31,76,31,92,31,25,31,224,31,220,31,220,30,5,31,164,31,120,31,87,31,87,30,108,31,108,30,108,29,127,31,17,31,17,30,17,29,17,28,17,27,208,31,163,31,78,31,133,31,194,31,8,31,28,31,28,30,28,29,230,31,197,31,197,30,11,31,3,31,200,31,200,30,162,31,218,31,212,31,90,31,90,30,109,31,24,31,24,30,174,31,174,30,26,31,107,31,83,31,29,31,37,31,79,31,224,31,78,31,78,30,83,31,22,31,52,31,186,31,157,31,44,31,144,31,246,31,246,30,62,31,216,31,221,31,164,31,164,30,99,31,147,31,139,31,74,31,197,31,138,31,176,31,244,31,185,31,188,31,14,31,139,31,139,30,120,31,33,31,194,31,177,31,140,31,95,31,87,31,149,31,25,31,176,31,176,30,76,31,46,31,115,31,107,31,2,31,23,31,139,31,139,30,104,31,189,31,252,31,252,30,12,31,127,31,248,31,88,31,118,31,150,31,228,31,104,31,104,30,216,31,89,31,189,31,194,31,239,31,120,31,120,30,120,29,217,31,217,30,78,31,198,31,198,30,20,31,239,31,48,31,48,30,63,31,105,31,207,31,207,30,88,31,169,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
