-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 368;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,107,0,0,0,115,0,22,0,177,0,59,0,56,0,132,0,97,0,64,0,0,0,0,0,0,0,220,0,0,0,173,0,177,0,85,0,249,0,177,0,8,0,135,0,238,0,0,0,11,0,36,0,160,0,43,0,182,0,201,0,18,0,0,0,90,0,31,0,63,0,0,0,26,0,121,0,0,0,242,0,0,0,211,0,0,0,128,0,6,0,207,0,154,0,193,0,0,0,145,0,54,0,157,0,29,0,17,0,46,0,131,0,251,0,50,0,187,0,212,0,82,0,0,0,176,0,200,0,49,0,83,0,0,0,72,0,20,0,166,0,23,0,219,0,95,0,135,0,105,0,14,0,0,0,0,0,0,0,197,0,118,0,105,0,114,0,94,0,65,0,59,0,168,0,127,0,110,0,248,0,21,0,0,0,142,0,179,0,176,0,213,0,28,0,225,0,0,0,251,0,87,0,156,0,234,0,67,0,54,0,0,0,244,0,0,0,176,0,41,0,161,0,249,0,0,0,185,0,84,0,111,0,52,0,84,0,87,0,220,0,0,0,124,0,171,0,102,0,139,0,0,0,91,0,0,0,117,0,92,0,20,0,0,0,34,0,116,0,0,0,87,0,158,0,49,0,0,0,243,0,196,0,237,0,0,0,48,0,81,0,254,0,47,0,198,0,109,0,41,0,124,0,0,0,26,0,0,0,204,0,42,0,69,0,0,0,144,0,53,0,138,0,50,0,69,0,152,0,48,0,252,0,0,0,16,0,240,0,51,0,99,0,36,0,187,0,82,0,31,0,109,0,0,0,202,0,193,0,145,0,0,0,138,0,1,0,202,0,107,0,222,0,0,0,48,0,181,0,76,0,26,0,200,0,113,0,28,0,6,0,192,0,5,0,0,0,42,0,146,0,2,0,0,0,0,0,104,0,210,0,135,0,30,0,107,0,58,0,0,0,7,0,0,0,170,0,70,0,212,0,140,0,107,0,0,0,219,0,38,0,113,0,64,0,182,0,0,0,216,0,0,0,132,0,74,0,133,0,222,0,0,0,0,0,70,0,248,0,34,0,111,0,0,0,214,0,145,0,209,0,161,0,11,0,230,0,53,0,224,0,159,0,198,0,140,0,167,0,0,0,54,0,28,0,63,0,0,0,86,0,129,0,155,0,102,0,161,0,254,0,17,0,155,0,136,0,0,0,0,0,193,0,96,0,219,0,116,0,0,0,155,0,215,0,124,0,236,0,208,0,37,0,0,0,203,0,0,0,73,0,166,0,0,0,21,0,215,0,2,0,43,0,31,0,152,0,240,0,236,0,0,0,49,0,219,0,225,0,230,0,143,0,241,0,0,0,0,0,179,0,202,0,138,0,158,0,87,0,138,0,70,0,51,0,168,0,0,0,252,0,173,0,129,0,240,0,111,0,158,0,195,0,0,0,0,0,134,0,0,0,177,0,76,0,115,0,44,0,0,0,175,0,48,0,1,0,164,0,0,0,128,0,149,0,86,0,224,0,244,0,145,0,102,0,7,0,126,0,10,0,185,0,0,0,214,0,118,0,81,0,120,0,105,0,48,0,18,0,53,0,0,0,46,0,0,0,119,0,182,0,251,0,0,0,250,0,43,0,214,0,106,0,106,0,237,0,110,0,230,0,205,0,84,0);
signal scenario_full  : scenario_type := (0,0,107,31,107,30,115,31,22,31,177,31,59,31,56,31,132,31,97,31,64,31,64,30,64,29,64,28,220,31,220,30,173,31,177,31,85,31,249,31,177,31,8,31,135,31,238,31,238,30,11,31,36,31,160,31,43,31,182,31,201,31,18,31,18,30,90,31,31,31,63,31,63,30,26,31,121,31,121,30,242,31,242,30,211,31,211,30,128,31,6,31,207,31,154,31,193,31,193,30,145,31,54,31,157,31,29,31,17,31,46,31,131,31,251,31,50,31,187,31,212,31,82,31,82,30,176,31,200,31,49,31,83,31,83,30,72,31,20,31,166,31,23,31,219,31,95,31,135,31,105,31,14,31,14,30,14,29,14,28,197,31,118,31,105,31,114,31,94,31,65,31,59,31,168,31,127,31,110,31,248,31,21,31,21,30,142,31,179,31,176,31,213,31,28,31,225,31,225,30,251,31,87,31,156,31,234,31,67,31,54,31,54,30,244,31,244,30,176,31,41,31,161,31,249,31,249,30,185,31,84,31,111,31,52,31,84,31,87,31,220,31,220,30,124,31,171,31,102,31,139,31,139,30,91,31,91,30,117,31,92,31,20,31,20,30,34,31,116,31,116,30,87,31,158,31,49,31,49,30,243,31,196,31,237,31,237,30,48,31,81,31,254,31,47,31,198,31,109,31,41,31,124,31,124,30,26,31,26,30,204,31,42,31,69,31,69,30,144,31,53,31,138,31,50,31,69,31,152,31,48,31,252,31,252,30,16,31,240,31,51,31,99,31,36,31,187,31,82,31,31,31,109,31,109,30,202,31,193,31,145,31,145,30,138,31,1,31,202,31,107,31,222,31,222,30,48,31,181,31,76,31,26,31,200,31,113,31,28,31,6,31,192,31,5,31,5,30,42,31,146,31,2,31,2,30,2,29,104,31,210,31,135,31,30,31,107,31,58,31,58,30,7,31,7,30,170,31,70,31,212,31,140,31,107,31,107,30,219,31,38,31,113,31,64,31,182,31,182,30,216,31,216,30,132,31,74,31,133,31,222,31,222,30,222,29,70,31,248,31,34,31,111,31,111,30,214,31,145,31,209,31,161,31,11,31,230,31,53,31,224,31,159,31,198,31,140,31,167,31,167,30,54,31,28,31,63,31,63,30,86,31,129,31,155,31,102,31,161,31,254,31,17,31,155,31,136,31,136,30,136,29,193,31,96,31,219,31,116,31,116,30,155,31,215,31,124,31,236,31,208,31,37,31,37,30,203,31,203,30,73,31,166,31,166,30,21,31,215,31,2,31,43,31,31,31,152,31,240,31,236,31,236,30,49,31,219,31,225,31,230,31,143,31,241,31,241,30,241,29,179,31,202,31,138,31,158,31,87,31,138,31,70,31,51,31,168,31,168,30,252,31,173,31,129,31,240,31,111,31,158,31,195,31,195,30,195,29,134,31,134,30,177,31,76,31,115,31,44,31,44,30,175,31,48,31,1,31,164,31,164,30,128,31,149,31,86,31,224,31,244,31,145,31,102,31,7,31,126,31,10,31,185,31,185,30,214,31,118,31,81,31,120,31,105,31,48,31,18,31,53,31,53,30,46,31,46,30,119,31,182,31,251,31,251,30,250,31,43,31,214,31,106,31,106,31,237,31,110,31,230,31,205,31,84,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
