-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_232 is
end project_tb_232;

architecture project_tb_arch_232 of project_tb_232 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 208;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,64,0,112,0,165,0,199,0,254,0,135,0,0,0,204,0,98,0,210,0,3,0,0,0,44,0,104,0,90,0,36,0,175,0,51,0,0,0,208,0,161,0,183,0,0,0,212,0,0,0,84,0,115,0,62,0,118,0,0,0,54,0,0,0,63,0,0,0,223,0,175,0,116,0,201,0,164,0,223,0,114,0,49,0,0,0,0,0,0,0,174,0,253,0,139,0,226,0,210,0,200,0,64,0,196,0,130,0,0,0,59,0,24,0,20,0,151,0,52,0,143,0,178,0,18,0,196,0,103,0,196,0,136,0,248,0,93,0,234,0,144,0,121,0,18,0,172,0,48,0,48,0,0,0,33,0,44,0,255,0,201,0,0,0,130,0,23,0,22,0,246,0,175,0,0,0,0,0,0,0,37,0,227,0,46,0,131,0,209,0,46,0,0,0,231,0,253,0,0,0,12,0,70,0,0,0,61,0,238,0,201,0,221,0,231,0,39,0,175,0,105,0,31,0,207,0,203,0,29,0,141,0,119,0,104,0,1,0,0,0,0,0,162,0,47,0,158,0,0,0,188,0,77,0,237,0,68,0,230,0,81,0,206,0,205,0,77,0,0,0,154,0,103,0,28,0,162,0,205,0,225,0,0,0,148,0,21,0,158,0,54,0,145,0,143,0,61,0,216,0,197,0,251,0,250,0,239,0,124,0,129,0,21,0,113,0,51,0,166,0,136,0,24,0,180,0,191,0,103,0,96,0,250,0,161,0,202,0,110,0,115,0,39,0,70,0,119,0,164,0,66,0,40,0,84,0,60,0,149,0,189,0,0,0,78,0,44,0,16,0,0,0,208,0,136,0,0,0,68,0,0,0,185,0,36,0,136,0,96,0,207,0,185,0,205,0,252,0,59,0,163,0,0,0,48,0,2,0,16,0,52,0,158,0);
signal scenario_full  : scenario_type := (0,0,64,31,112,31,165,31,199,31,254,31,135,31,135,30,204,31,98,31,210,31,3,31,3,30,44,31,104,31,90,31,36,31,175,31,51,31,51,30,208,31,161,31,183,31,183,30,212,31,212,30,84,31,115,31,62,31,118,31,118,30,54,31,54,30,63,31,63,30,223,31,175,31,116,31,201,31,164,31,223,31,114,31,49,31,49,30,49,29,49,28,174,31,253,31,139,31,226,31,210,31,200,31,64,31,196,31,130,31,130,30,59,31,24,31,20,31,151,31,52,31,143,31,178,31,18,31,196,31,103,31,196,31,136,31,248,31,93,31,234,31,144,31,121,31,18,31,172,31,48,31,48,31,48,30,33,31,44,31,255,31,201,31,201,30,130,31,23,31,22,31,246,31,175,31,175,30,175,29,175,28,37,31,227,31,46,31,131,31,209,31,46,31,46,30,231,31,253,31,253,30,12,31,70,31,70,30,61,31,238,31,201,31,221,31,231,31,39,31,175,31,105,31,31,31,207,31,203,31,29,31,141,31,119,31,104,31,1,31,1,30,1,29,162,31,47,31,158,31,158,30,188,31,77,31,237,31,68,31,230,31,81,31,206,31,205,31,77,31,77,30,154,31,103,31,28,31,162,31,205,31,225,31,225,30,148,31,21,31,158,31,54,31,145,31,143,31,61,31,216,31,197,31,251,31,250,31,239,31,124,31,129,31,21,31,113,31,51,31,166,31,136,31,24,31,180,31,191,31,103,31,96,31,250,31,161,31,202,31,110,31,115,31,39,31,70,31,119,31,164,31,66,31,40,31,84,31,60,31,149,31,189,31,189,30,78,31,44,31,16,31,16,30,208,31,136,31,136,30,68,31,68,30,185,31,36,31,136,31,96,31,207,31,185,31,205,31,252,31,59,31,163,31,163,30,48,31,2,31,16,31,52,31,158,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
