-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 453;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (86,0,0,0,204,0,19,0,110,0,203,0,101,0,18,0,75,0,224,0,75,0,58,0,253,0,143,0,198,0,193,0,30,0,108,0,243,0,156,0,0,0,0,0,0,0,0,0,0,0,164,0,101,0,103,0,0,0,110,0,227,0,39,0,0,0,243,0,240,0,0,0,204,0,0,0,7,0,63,0,247,0,0,0,127,0,147,0,99,0,9,0,2,0,62,0,0,0,221,0,19,0,0,0,230,0,4,0,106,0,36,0,118,0,169,0,183,0,239,0,0,0,212,0,0,0,149,0,55,0,60,0,204,0,22,0,71,0,0,0,115,0,120,0,229,0,217,0,43,0,205,0,28,0,162,0,200,0,239,0,109,0,44,0,68,0,85,0,185,0,159,0,0,0,252,0,247,0,0,0,0,0,54,0,243,0,142,0,119,0,144,0,79,0,0,0,207,0,1,0,251,0,187,0,67,0,243,0,149,0,117,0,146,0,114,0,3,0,0,0,50,0,0,0,48,0,131,0,150,0,77,0,107,0,23,0,127,0,254,0,89,0,114,0,106,0,243,0,22,0,54,0,50,0,178,0,167,0,113,0,70,0,130,0,78,0,235,0,82,0,205,0,38,0,66,0,1,0,188,0,193,0,207,0,27,0,121,0,206,0,170,0,25,0,0,0,0,0,44,0,0,0,35,0,105,0,228,0,117,0,95,0,0,0,0,0,246,0,148,0,6,0,201,0,36,0,66,0,131,0,209,0,102,0,196,0,141,0,160,0,21,0,181,0,154,0,74,0,104,0,161,0,14,0,41,0,0,0,118,0,50,0,58,0,0,0,191,0,250,0,79,0,0,0,31,0,66,0,24,0,0,0,177,0,247,0,36,0,30,0,170,0,229,0,76,0,173,0,138,0,11,0,208,0,0,0,100,0,70,0,185,0,179,0,182,0,232,0,210,0,40,0,63,0,0,0,0,0,59,0,155,0,0,0,177,0,156,0,2,0,243,0,166,0,55,0,32,0,0,0,49,0,85,0,134,0,97,0,212,0,27,0,0,0,8,0,13,0,0,0,157,0,14,0,222,0,182,0,107,0,3,0,254,0,98,0,0,0,227,0,0,0,0,0,100,0,153,0,72,0,42,0,94,0,0,0,1,0,28,0,125,0,42,0,203,0,105,0,87,0,165,0,0,0,79,0,226,0,102,0,106,0,16,0,78,0,0,0,223,0,116,0,243,0,92,0,0,0,114,0,140,0,44,0,203,0,64,0,92,0,92,0,241,0,9,0,248,0,4,0,205,0,60,0,150,0,169,0,0,0,119,0,117,0,0,0,216,0,231,0,171,0,0,0,165,0,134,0,119,0,63,0,149,0,0,0,211,0,0,0,134,0,0,0,36,0,0,0,28,0,233,0,237,0,236,0,185,0,0,0,109,0,0,0,0,0,168,0,131,0,122,0,126,0,186,0,91,0,216,0,113,0,104,0,238,0,224,0,249,0,172,0,108,0,61,0,144,0,43,0,123,0,0,0,116,0,232,0,246,0,230,0,54,0,168,0,75,0,195,0,178,0,126,0,0,0,244,0,31,0,29,0,136,0,177,0,226,0,146,0,77,0,140,0,233,0,104,0,36,0,170,0,166,0,65,0,182,0,121,0,121,0,69,0,168,0,0,0,90,0,69,0,189,0,180,0,246,0,182,0,3,0,36,0,0,0,61,0,162,0,87,0,26,0,40,0,171,0,217,0,168,0,129,0,186,0,0,0,230,0,82,0,133,0,0,0,166,0,0,0,173,0,183,0,44,0,205,0,3,0,225,0,248,0,235,0,191,0,58,0,62,0,59,0,202,0,110,0,0,0,254,0,37,0,95,0,146,0,69,0,244,0,211,0,218,0,188,0,243,0,20,0,0,0,238,0,197,0,70,0,63,0,72,0,99,0,157,0,53,0,254,0,230,0,0,0,99,0,0,0,0,0,211,0,179,0,0,0,41,0,113,0,0,0,0,0,86,0,0,0,89,0,0,0,0,0,104,0,24,0,199,0,160,0,73,0);
signal scenario_full  : scenario_type := (86,31,86,30,204,31,19,31,110,31,203,31,101,31,18,31,75,31,224,31,75,31,58,31,253,31,143,31,198,31,193,31,30,31,108,31,243,31,156,31,156,30,156,29,156,28,156,27,156,26,164,31,101,31,103,31,103,30,110,31,227,31,39,31,39,30,243,31,240,31,240,30,204,31,204,30,7,31,63,31,247,31,247,30,127,31,147,31,99,31,9,31,2,31,62,31,62,30,221,31,19,31,19,30,230,31,4,31,106,31,36,31,118,31,169,31,183,31,239,31,239,30,212,31,212,30,149,31,55,31,60,31,204,31,22,31,71,31,71,30,115,31,120,31,229,31,217,31,43,31,205,31,28,31,162,31,200,31,239,31,109,31,44,31,68,31,85,31,185,31,159,31,159,30,252,31,247,31,247,30,247,29,54,31,243,31,142,31,119,31,144,31,79,31,79,30,207,31,1,31,251,31,187,31,67,31,243,31,149,31,117,31,146,31,114,31,3,31,3,30,50,31,50,30,48,31,131,31,150,31,77,31,107,31,23,31,127,31,254,31,89,31,114,31,106,31,243,31,22,31,54,31,50,31,178,31,167,31,113,31,70,31,130,31,78,31,235,31,82,31,205,31,38,31,66,31,1,31,188,31,193,31,207,31,27,31,121,31,206,31,170,31,25,31,25,30,25,29,44,31,44,30,35,31,105,31,228,31,117,31,95,31,95,30,95,29,246,31,148,31,6,31,201,31,36,31,66,31,131,31,209,31,102,31,196,31,141,31,160,31,21,31,181,31,154,31,74,31,104,31,161,31,14,31,41,31,41,30,118,31,50,31,58,31,58,30,191,31,250,31,79,31,79,30,31,31,66,31,24,31,24,30,177,31,247,31,36,31,30,31,170,31,229,31,76,31,173,31,138,31,11,31,208,31,208,30,100,31,70,31,185,31,179,31,182,31,232,31,210,31,40,31,63,31,63,30,63,29,59,31,155,31,155,30,177,31,156,31,2,31,243,31,166,31,55,31,32,31,32,30,49,31,85,31,134,31,97,31,212,31,27,31,27,30,8,31,13,31,13,30,157,31,14,31,222,31,182,31,107,31,3,31,254,31,98,31,98,30,227,31,227,30,227,29,100,31,153,31,72,31,42,31,94,31,94,30,1,31,28,31,125,31,42,31,203,31,105,31,87,31,165,31,165,30,79,31,226,31,102,31,106,31,16,31,78,31,78,30,223,31,116,31,243,31,92,31,92,30,114,31,140,31,44,31,203,31,64,31,92,31,92,31,241,31,9,31,248,31,4,31,205,31,60,31,150,31,169,31,169,30,119,31,117,31,117,30,216,31,231,31,171,31,171,30,165,31,134,31,119,31,63,31,149,31,149,30,211,31,211,30,134,31,134,30,36,31,36,30,28,31,233,31,237,31,236,31,185,31,185,30,109,31,109,30,109,29,168,31,131,31,122,31,126,31,186,31,91,31,216,31,113,31,104,31,238,31,224,31,249,31,172,31,108,31,61,31,144,31,43,31,123,31,123,30,116,31,232,31,246,31,230,31,54,31,168,31,75,31,195,31,178,31,126,31,126,30,244,31,31,31,29,31,136,31,177,31,226,31,146,31,77,31,140,31,233,31,104,31,36,31,170,31,166,31,65,31,182,31,121,31,121,31,69,31,168,31,168,30,90,31,69,31,189,31,180,31,246,31,182,31,3,31,36,31,36,30,61,31,162,31,87,31,26,31,40,31,171,31,217,31,168,31,129,31,186,31,186,30,230,31,82,31,133,31,133,30,166,31,166,30,173,31,183,31,44,31,205,31,3,31,225,31,248,31,235,31,191,31,58,31,62,31,59,31,202,31,110,31,110,30,254,31,37,31,95,31,146,31,69,31,244,31,211,31,218,31,188,31,243,31,20,31,20,30,238,31,197,31,70,31,63,31,72,31,99,31,157,31,53,31,254,31,230,31,230,30,99,31,99,30,99,29,211,31,179,31,179,30,41,31,113,31,113,30,113,29,86,31,86,30,89,31,89,30,89,29,104,31,24,31,199,31,160,31,73,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
