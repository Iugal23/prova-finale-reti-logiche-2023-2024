-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_374 is
end project_tb_374;

architecture project_tb_arch_374 of project_tb_374 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 770;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (199,0,242,0,241,0,48,0,232,0,96,0,186,0,0,0,113,0,23,0,28,0,236,0,220,0,213,0,13,0,209,0,10,0,92,0,0,0,189,0,177,0,226,0,247,0,119,0,136,0,205,0,30,0,178,0,44,0,134,0,194,0,94,0,146,0,0,0,0,0,238,0,66,0,227,0,0,0,98,0,37,0,162,0,10,0,0,0,0,0,22,0,78,0,25,0,6,0,59,0,140,0,87,0,11,0,162,0,78,0,242,0,151,0,0,0,35,0,171,0,149,0,196,0,139,0,29,0,215,0,32,0,152,0,149,0,108,0,118,0,163,0,203,0,237,0,61,0,231,0,20,0,0,0,92,0,177,0,120,0,88,0,65,0,108,0,161,0,68,0,172,0,85,0,84,0,53,0,188,0,94,0,184,0,0,0,0,0,135,0,253,0,139,0,52,0,0,0,0,0,0,0,165,0,0,0,166,0,93,0,120,0,36,0,175,0,22,0,114,0,0,0,67,0,239,0,44,0,239,0,105,0,0,0,0,0,97,0,104,0,178,0,0,0,0,0,0,0,131,0,0,0,111,0,95,0,13,0,5,0,242,0,10,0,126,0,0,0,235,0,51,0,242,0,242,0,18,0,206,0,212,0,161,0,43,0,170,0,231,0,121,0,129,0,241,0,6,0,189,0,247,0,92,0,96,0,44,0,49,0,106,0,130,0,0,0,192,0,252,0,0,0,51,0,140,0,28,0,12,0,44,0,0,0,196,0,216,0,89,0,0,0,0,0,146,0,88,0,61,0,89,0,34,0,24,0,73,0,213,0,0,0,0,0,0,0,31,0,251,0,0,0,33,0,174,0,8,0,0,0,0,0,169,0,84,0,79,0,63,0,174,0,65,0,82,0,0,0,231,0,98,0,240,0,204,0,105,0,0,0,38,0,0,0,82,0,249,0,122,0,173,0,13,0,46,0,226,0,44,0,125,0,0,0,77,0,28,0,201,0,190,0,54,0,0,0,255,0,0,0,0,0,172,0,94,0,0,0,156,0,127,0,254,0,0,0,238,0,237,0,115,0,103,0,238,0,131,0,132,0,208,0,105,0,112,0,0,0,147,0,137,0,37,0,188,0,57,0,232,0,0,0,210,0,52,0,138,0,20,0,164,0,161,0,233,0,0,0,51,0,249,0,186,0,204,0,77,0,153,0,139,0,0,0,98,0,0,0,52,0,0,0,78,0,0,0,124,0,86,0,192,0,215,0,208,0,94,0,225,0,206,0,0,0,134,0,221,0,108,0,174,0,182,0,17,0,252,0,221,0,206,0,69,0,0,0,48,0,164,0,46,0,239,0,0,0,175,0,144,0,46,0,0,0,1,0,39,0,80,0,20,0,211,0,0,0,111,0,0,0,90,0,172,0,53,0,0,0,103,0,0,0,0,0,103,0,47,0,0,0,39,0,0,0,0,0,123,0,0,0,56,0,121,0,176,0,71,0,0,0,69,0,0,0,0,0,255,0,18,0,0,0,200,0,111,0,161,0,5,0,50,0,44,0,159,0,21,0,0,0,0,0,0,0,85,0,127,0,134,0,67,0,152,0,98,0,16,0,0,0,0,0,155,0,0,0,197,0,92,0,180,0,11,0,13,0,0,0,132,0,112,0,13,0,164,0,150,0,202,0,190,0,178,0,0,0,102,0,27,0,0,0,139,0,58,0,12,0,61,0,89,0,21,0,37,0,2,0,152,0,249,0,0,0,0,0,85,0,40,0,225,0,108,0,99,0,43,0,109,0,0,0,178,0,34,0,0,0,16,0,107,0,45,0,210,0,0,0,249,0,122,0,238,0,5,0,219,0,80,0,157,0,57,0,239,0,41,0,0,0,0,0,228,0,18,0,154,0,115,0,55,0,100,0,85,0,0,0,0,0,0,0,0,0,227,0,144,0,13,0,2,0,45,0,105,0,97,0,220,0,109,0,181,0,230,0,10,0,0,0,139,0,191,0,163,0,88,0,186,0,123,0,106,0,235,0,116,0,121,0,190,0,246,0,114,0,0,0,138,0,163,0,187,0,0,0,36,0,3,0,60,0,156,0,212,0,180,0,246,0,162,0,63,0,109,0,181,0,0,0,228,0,19,0,230,0,243,0,83,0,232,0,166,0,122,0,147,0,65,0,75,0,37,0,39,0,99,0,75,0,242,0,226,0,0,0,14,0,105,0,158,0,254,0,25,0,0,0,0,0,197,0,45,0,95,0,245,0,54,0,148,0,70,0,99,0,243,0,209,0,254,0,100,0,0,0,178,0,212,0,83,0,255,0,0,0,0,0,46,0,224,0,26,0,137,0,21,0,56,0,0,0,16,0,30,0,230,0,0,0,0,0,0,0,0,0,233,0,13,0,87,0,156,0,239,0,167,0,17,0,68,0,38,0,101,0,125,0,55,0,145,0,99,0,233,0,145,0,142,0,137,0,0,0,197,0,89,0,34,0,67,0,53,0,0,0,17,0,0,0,43,0,145,0,242,0,38,0,26,0,0,0,211,0,0,0,100,0,216,0,17,0,26,0,194,0,4,0,77,0,75,0,14,0,37,0,42,0,132,0,16,0,151,0,66,0,192,0,0,0,242,0,106,0,86,0,0,0,211,0,28,0,217,0,67,0,228,0,0,0,76,0,133,0,68,0,215,0,1,0,0,0,0,0,211,0,20,0,226,0,226,0,21,0,0,0,121,0,217,0,208,0,177,0,46,0,255,0,0,0,236,0,0,0,22,0,0,0,0,0,0,0,68,0,13,0,231,0,5,0,150,0,14,0,34,0,134,0,186,0,0,0,0,0,206,0,137,0,172,0,125,0,232,0,63,0,223,0,32,0,191,0,216,0,51,0,215,0,224,0,244,0,0,0,45,0,3,0,0,0,65,0,158,0,0,0,254,0,17,0,0,0,106,0,214,0,182,0,19,0,182,0,120,0,98,0,0,0,0,0,37,0,119,0,254,0,189,0,100,0,231,0,187,0,176,0,0,0,248,0,63,0,30,0,218,0,170,0,55,0,0,0,0,0,0,0,40,0,198,0,35,0,217,0,249,0,111,0,0,0,96,0,185,0,66,0,168,0,0,0,61,0,191,0,97,0,0,0,10,0,59,0,175,0,61,0,115,0,142,0,138,0,224,0,14,0,177,0,0,0,0,0,134,0,5,0,194,0,236,0,99,0,231,0,45,0,155,0,177,0,55,0,62,0,110,0,0,0,218,0,145,0,118,0,226,0,0,0,43,0,0,0,0,0,122,0,225,0,241,0,211,0,122,0,236,0,0,0,2,0,12,0,0,0,57,0,4,0,212,0,0,0,66,0,171,0,250,0,167,0,0,0,14,0,0,0,88,0,200,0,41,0,134,0,8,0,41,0,0,0,108,0,152,0,9,0,98,0,135,0,130,0,141,0,0,0,0,0,0,0,7,0,46,0,5,0,220,0,62,0);
signal scenario_full  : scenario_type := (199,31,242,31,241,31,48,31,232,31,96,31,186,31,186,30,113,31,23,31,28,31,236,31,220,31,213,31,13,31,209,31,10,31,92,31,92,30,189,31,177,31,226,31,247,31,119,31,136,31,205,31,30,31,178,31,44,31,134,31,194,31,94,31,146,31,146,30,146,29,238,31,66,31,227,31,227,30,98,31,37,31,162,31,10,31,10,30,10,29,22,31,78,31,25,31,6,31,59,31,140,31,87,31,11,31,162,31,78,31,242,31,151,31,151,30,35,31,171,31,149,31,196,31,139,31,29,31,215,31,32,31,152,31,149,31,108,31,118,31,163,31,203,31,237,31,61,31,231,31,20,31,20,30,92,31,177,31,120,31,88,31,65,31,108,31,161,31,68,31,172,31,85,31,84,31,53,31,188,31,94,31,184,31,184,30,184,29,135,31,253,31,139,31,52,31,52,30,52,29,52,28,165,31,165,30,166,31,93,31,120,31,36,31,175,31,22,31,114,31,114,30,67,31,239,31,44,31,239,31,105,31,105,30,105,29,97,31,104,31,178,31,178,30,178,29,178,28,131,31,131,30,111,31,95,31,13,31,5,31,242,31,10,31,126,31,126,30,235,31,51,31,242,31,242,31,18,31,206,31,212,31,161,31,43,31,170,31,231,31,121,31,129,31,241,31,6,31,189,31,247,31,92,31,96,31,44,31,49,31,106,31,130,31,130,30,192,31,252,31,252,30,51,31,140,31,28,31,12,31,44,31,44,30,196,31,216,31,89,31,89,30,89,29,146,31,88,31,61,31,89,31,34,31,24,31,73,31,213,31,213,30,213,29,213,28,31,31,251,31,251,30,33,31,174,31,8,31,8,30,8,29,169,31,84,31,79,31,63,31,174,31,65,31,82,31,82,30,231,31,98,31,240,31,204,31,105,31,105,30,38,31,38,30,82,31,249,31,122,31,173,31,13,31,46,31,226,31,44,31,125,31,125,30,77,31,28,31,201,31,190,31,54,31,54,30,255,31,255,30,255,29,172,31,94,31,94,30,156,31,127,31,254,31,254,30,238,31,237,31,115,31,103,31,238,31,131,31,132,31,208,31,105,31,112,31,112,30,147,31,137,31,37,31,188,31,57,31,232,31,232,30,210,31,52,31,138,31,20,31,164,31,161,31,233,31,233,30,51,31,249,31,186,31,204,31,77,31,153,31,139,31,139,30,98,31,98,30,52,31,52,30,78,31,78,30,124,31,86,31,192,31,215,31,208,31,94,31,225,31,206,31,206,30,134,31,221,31,108,31,174,31,182,31,17,31,252,31,221,31,206,31,69,31,69,30,48,31,164,31,46,31,239,31,239,30,175,31,144,31,46,31,46,30,1,31,39,31,80,31,20,31,211,31,211,30,111,31,111,30,90,31,172,31,53,31,53,30,103,31,103,30,103,29,103,31,47,31,47,30,39,31,39,30,39,29,123,31,123,30,56,31,121,31,176,31,71,31,71,30,69,31,69,30,69,29,255,31,18,31,18,30,200,31,111,31,161,31,5,31,50,31,44,31,159,31,21,31,21,30,21,29,21,28,85,31,127,31,134,31,67,31,152,31,98,31,16,31,16,30,16,29,155,31,155,30,197,31,92,31,180,31,11,31,13,31,13,30,132,31,112,31,13,31,164,31,150,31,202,31,190,31,178,31,178,30,102,31,27,31,27,30,139,31,58,31,12,31,61,31,89,31,21,31,37,31,2,31,152,31,249,31,249,30,249,29,85,31,40,31,225,31,108,31,99,31,43,31,109,31,109,30,178,31,34,31,34,30,16,31,107,31,45,31,210,31,210,30,249,31,122,31,238,31,5,31,219,31,80,31,157,31,57,31,239,31,41,31,41,30,41,29,228,31,18,31,154,31,115,31,55,31,100,31,85,31,85,30,85,29,85,28,85,27,227,31,144,31,13,31,2,31,45,31,105,31,97,31,220,31,109,31,181,31,230,31,10,31,10,30,139,31,191,31,163,31,88,31,186,31,123,31,106,31,235,31,116,31,121,31,190,31,246,31,114,31,114,30,138,31,163,31,187,31,187,30,36,31,3,31,60,31,156,31,212,31,180,31,246,31,162,31,63,31,109,31,181,31,181,30,228,31,19,31,230,31,243,31,83,31,232,31,166,31,122,31,147,31,65,31,75,31,37,31,39,31,99,31,75,31,242,31,226,31,226,30,14,31,105,31,158,31,254,31,25,31,25,30,25,29,197,31,45,31,95,31,245,31,54,31,148,31,70,31,99,31,243,31,209,31,254,31,100,31,100,30,178,31,212,31,83,31,255,31,255,30,255,29,46,31,224,31,26,31,137,31,21,31,56,31,56,30,16,31,30,31,230,31,230,30,230,29,230,28,230,27,233,31,13,31,87,31,156,31,239,31,167,31,17,31,68,31,38,31,101,31,125,31,55,31,145,31,99,31,233,31,145,31,142,31,137,31,137,30,197,31,89,31,34,31,67,31,53,31,53,30,17,31,17,30,43,31,145,31,242,31,38,31,26,31,26,30,211,31,211,30,100,31,216,31,17,31,26,31,194,31,4,31,77,31,75,31,14,31,37,31,42,31,132,31,16,31,151,31,66,31,192,31,192,30,242,31,106,31,86,31,86,30,211,31,28,31,217,31,67,31,228,31,228,30,76,31,133,31,68,31,215,31,1,31,1,30,1,29,211,31,20,31,226,31,226,31,21,31,21,30,121,31,217,31,208,31,177,31,46,31,255,31,255,30,236,31,236,30,22,31,22,30,22,29,22,28,68,31,13,31,231,31,5,31,150,31,14,31,34,31,134,31,186,31,186,30,186,29,206,31,137,31,172,31,125,31,232,31,63,31,223,31,32,31,191,31,216,31,51,31,215,31,224,31,244,31,244,30,45,31,3,31,3,30,65,31,158,31,158,30,254,31,17,31,17,30,106,31,214,31,182,31,19,31,182,31,120,31,98,31,98,30,98,29,37,31,119,31,254,31,189,31,100,31,231,31,187,31,176,31,176,30,248,31,63,31,30,31,218,31,170,31,55,31,55,30,55,29,55,28,40,31,198,31,35,31,217,31,249,31,111,31,111,30,96,31,185,31,66,31,168,31,168,30,61,31,191,31,97,31,97,30,10,31,59,31,175,31,61,31,115,31,142,31,138,31,224,31,14,31,177,31,177,30,177,29,134,31,5,31,194,31,236,31,99,31,231,31,45,31,155,31,177,31,55,31,62,31,110,31,110,30,218,31,145,31,118,31,226,31,226,30,43,31,43,30,43,29,122,31,225,31,241,31,211,31,122,31,236,31,236,30,2,31,12,31,12,30,57,31,4,31,212,31,212,30,66,31,171,31,250,31,167,31,167,30,14,31,14,30,88,31,200,31,41,31,134,31,8,31,41,31,41,30,108,31,152,31,9,31,98,31,135,31,130,31,141,31,141,30,141,29,141,28,7,31,46,31,5,31,220,31,62,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
