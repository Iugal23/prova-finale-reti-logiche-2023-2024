-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 646;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (6,0,17,0,140,0,125,0,0,0,179,0,117,0,0,0,91,0,0,0,247,0,194,0,74,0,0,0,179,0,0,0,165,0,141,0,0,0,0,0,133,0,0,0,0,0,0,0,68,0,0,0,233,0,184,0,142,0,0,0,0,0,229,0,233,0,233,0,17,0,95,0,112,0,172,0,71,0,247,0,106,0,0,0,176,0,16,0,0,0,0,0,135,0,0,0,138,0,118,0,4,0,0,0,139,0,125,0,45,0,198,0,0,0,137,0,0,0,159,0,166,0,124,0,104,0,137,0,0,0,55,0,117,0,180,0,172,0,87,0,172,0,24,0,186,0,186,0,49,0,0,0,194,0,102,0,72,0,53,0,0,0,0,0,0,0,58,0,0,0,185,0,211,0,0,0,216,0,101,0,230,0,166,0,0,0,47,0,16,0,0,0,0,0,205,0,32,0,208,0,152,0,233,0,219,0,134,0,191,0,0,0,117,0,1,0,68,0,60,0,0,0,217,0,186,0,170,0,113,0,121,0,18,0,0,0,92,0,65,0,0,0,0,0,146,0,134,0,238,0,0,0,0,0,82,0,75,0,104,0,72,0,17,0,83,0,254,0,0,0,58,0,248,0,93,0,110,0,0,0,5,0,117,0,33,0,216,0,154,0,0,0,167,0,63,0,250,0,36,0,222,0,68,0,153,0,0,0,107,0,51,0,82,0,28,0,175,0,0,0,224,0,2,0,0,0,196,0,181,0,90,0,102,0,0,0,135,0,249,0,0,0,139,0,69,0,0,0,235,0,141,0,0,0,62,0,0,0,250,0,153,0,232,0,46,0,117,0,68,0,242,0,121,0,0,0,54,0,202,0,169,0,155,0,15,0,103,0,26,0,114,0,165,0,99,0,224,0,0,0,203,0,0,0,108,0,152,0,0,0,253,0,255,0,207,0,0,0,200,0,45,0,247,0,208,0,254,0,172,0,115,0,121,0,103,0,148,0,22,0,0,0,56,0,104,0,184,0,48,0,17,0,102,0,38,0,40,0,68,0,103,0,106,0,253,0,202,0,105,0,55,0,110,0,234,0,193,0,0,0,238,0,184,0,253,0,110,0,147,0,189,0,146,0,175,0,136,0,154,0,31,0,63,0,63,0,142,0,187,0,0,0,173,0,106,0,101,0,186,0,0,0,0,0,115,0,50,0,0,0,0,0,64,0,31,0,185,0,185,0,226,0,0,0,15,0,209,0,0,0,0,0,189,0,185,0,26,0,25,0,48,0,67,0,135,0,0,0,174,0,3,0,145,0,43,0,19,0,1,0,199,0,183,0,0,0,242,0,126,0,57,0,0,0,170,0,216,0,178,0,143,0,180,0,188,0,23,0,85,0,0,0,68,0,39,0,0,0,0,0,122,0,234,0,2,0,0,0,151,0,0,0,157,0,24,0,67,0,15,0,184,0,133,0,205,0,7,0,230,0,193,0,26,0,240,0,114,0,17,0,0,0,146,0,140,0,49,0,149,0,223,0,0,0,83,0,26,0,49,0,41,0,0,0,10,0,116,0,125,0,0,0,68,0,81,0,241,0,200,0,0,0,195,0,170,0,198,0,0,0,0,0,106,0,41,0,122,0,254,0,134,0,0,0,153,0,18,0,94,0,35,0,162,0,91,0,2,0,52,0,92,0,111,0,89,0,49,0,199,0,146,0,34,0,39,0,0,0,46,0,165,0,231,0,75,0,238,0,234,0,6,0,155,0,35,0,109,0,178,0,203,0,106,0,210,0,0,0,18,0,48,0,172,0,2,0,99,0,145,0,74,0,230,0,111,0,113,0,33,0,146,0,234,0,149,0,180,0,55,0,0,0,0,0,178,0,210,0,0,0,208,0,0,0,171,0,214,0,47,0,157,0,130,0,87,0,65,0,0,0,45,0,57,0,0,0,58,0,0,0,251,0,14,0,10,0,140,0,29,0,187,0,40,0,0,0,169,0,149,0,100,0,168,0,11,0,147,0,155,0,178,0,149,0,162,0,185,0,231,0,173,0,19,0,0,0,0,0,3,0,88,0,214,0,0,0,173,0,0,0,0,0,107,0,131,0,151,0,158,0,158,0,0,0,90,0,215,0,41,0,0,0,4,0,194,0,211,0,149,0,26,0,2,0,239,0,175,0,0,0,0,0,168,0,132,0,223,0,114,0,94,0,220,0,101,0,0,0,0,0,243,0,165,0,248,0,164,0,10,0,0,0,73,0,172,0,0,0,0,0,99,0,0,0,23,0,228,0,206,0,8,0,0,0,232,0,11,0,62,0,0,0,5,0,0,0,251,0,55,0,204,0,144,0,2,0,0,0,201,0,0,0,139,0,222,0,254,0,97,0,0,0,37,0,57,0,48,0,171,0,0,0,73,0,147,0,95,0,102,0,0,0,63,0,31,0,240,0,53,0,172,0,252,0,30,0,221,0,0,0,234,0,247,0,1,0,139,0,66,0,254,0,0,0,100,0,24,0,0,0,89,0,11,0,146,0,223,0,168,0,124,0,145,0,242,0,103,0,0,0,144,0,228,0,0,0,95,0,0,0,8,0,172,0,55,0,64,0,0,0,15,0,78,0,107,0,147,0,237,0,252,0,124,0,68,0,178,0,36,0,173,0,0,0,160,0,195,0,248,0,0,0,241,0,117,0,0,0,15,0,145,0,0,0,33,0,15,0,0,0,26,0,67,0,255,0,10,0,0,0,0,0,74,0,227,0,93,0,0,0,0,0,181,0,1,0,107,0,153,0,185,0,141,0,125,0,74,0,112,0,31,0,11,0,0,0,26,0,0,0,96,0,133,0,14,0,226,0,0,0,191,0,0,0,164,0,60,0,158,0,161,0,0,0,0,0,0,0,0,0,67,0,18,0,245,0,122,0,199,0,0,0);
signal scenario_full  : scenario_type := (6,31,17,31,140,31,125,31,125,30,179,31,117,31,117,30,91,31,91,30,247,31,194,31,74,31,74,30,179,31,179,30,165,31,141,31,141,30,141,29,133,31,133,30,133,29,133,28,68,31,68,30,233,31,184,31,142,31,142,30,142,29,229,31,233,31,233,31,17,31,95,31,112,31,172,31,71,31,247,31,106,31,106,30,176,31,16,31,16,30,16,29,135,31,135,30,138,31,118,31,4,31,4,30,139,31,125,31,45,31,198,31,198,30,137,31,137,30,159,31,166,31,124,31,104,31,137,31,137,30,55,31,117,31,180,31,172,31,87,31,172,31,24,31,186,31,186,31,49,31,49,30,194,31,102,31,72,31,53,31,53,30,53,29,53,28,58,31,58,30,185,31,211,31,211,30,216,31,101,31,230,31,166,31,166,30,47,31,16,31,16,30,16,29,205,31,32,31,208,31,152,31,233,31,219,31,134,31,191,31,191,30,117,31,1,31,68,31,60,31,60,30,217,31,186,31,170,31,113,31,121,31,18,31,18,30,92,31,65,31,65,30,65,29,146,31,134,31,238,31,238,30,238,29,82,31,75,31,104,31,72,31,17,31,83,31,254,31,254,30,58,31,248,31,93,31,110,31,110,30,5,31,117,31,33,31,216,31,154,31,154,30,167,31,63,31,250,31,36,31,222,31,68,31,153,31,153,30,107,31,51,31,82,31,28,31,175,31,175,30,224,31,2,31,2,30,196,31,181,31,90,31,102,31,102,30,135,31,249,31,249,30,139,31,69,31,69,30,235,31,141,31,141,30,62,31,62,30,250,31,153,31,232,31,46,31,117,31,68,31,242,31,121,31,121,30,54,31,202,31,169,31,155,31,15,31,103,31,26,31,114,31,165,31,99,31,224,31,224,30,203,31,203,30,108,31,152,31,152,30,253,31,255,31,207,31,207,30,200,31,45,31,247,31,208,31,254,31,172,31,115,31,121,31,103,31,148,31,22,31,22,30,56,31,104,31,184,31,48,31,17,31,102,31,38,31,40,31,68,31,103,31,106,31,253,31,202,31,105,31,55,31,110,31,234,31,193,31,193,30,238,31,184,31,253,31,110,31,147,31,189,31,146,31,175,31,136,31,154,31,31,31,63,31,63,31,142,31,187,31,187,30,173,31,106,31,101,31,186,31,186,30,186,29,115,31,50,31,50,30,50,29,64,31,31,31,185,31,185,31,226,31,226,30,15,31,209,31,209,30,209,29,189,31,185,31,26,31,25,31,48,31,67,31,135,31,135,30,174,31,3,31,145,31,43,31,19,31,1,31,199,31,183,31,183,30,242,31,126,31,57,31,57,30,170,31,216,31,178,31,143,31,180,31,188,31,23,31,85,31,85,30,68,31,39,31,39,30,39,29,122,31,234,31,2,31,2,30,151,31,151,30,157,31,24,31,67,31,15,31,184,31,133,31,205,31,7,31,230,31,193,31,26,31,240,31,114,31,17,31,17,30,146,31,140,31,49,31,149,31,223,31,223,30,83,31,26,31,49,31,41,31,41,30,10,31,116,31,125,31,125,30,68,31,81,31,241,31,200,31,200,30,195,31,170,31,198,31,198,30,198,29,106,31,41,31,122,31,254,31,134,31,134,30,153,31,18,31,94,31,35,31,162,31,91,31,2,31,52,31,92,31,111,31,89,31,49,31,199,31,146,31,34,31,39,31,39,30,46,31,165,31,231,31,75,31,238,31,234,31,6,31,155,31,35,31,109,31,178,31,203,31,106,31,210,31,210,30,18,31,48,31,172,31,2,31,99,31,145,31,74,31,230,31,111,31,113,31,33,31,146,31,234,31,149,31,180,31,55,31,55,30,55,29,178,31,210,31,210,30,208,31,208,30,171,31,214,31,47,31,157,31,130,31,87,31,65,31,65,30,45,31,57,31,57,30,58,31,58,30,251,31,14,31,10,31,140,31,29,31,187,31,40,31,40,30,169,31,149,31,100,31,168,31,11,31,147,31,155,31,178,31,149,31,162,31,185,31,231,31,173,31,19,31,19,30,19,29,3,31,88,31,214,31,214,30,173,31,173,30,173,29,107,31,131,31,151,31,158,31,158,31,158,30,90,31,215,31,41,31,41,30,4,31,194,31,211,31,149,31,26,31,2,31,239,31,175,31,175,30,175,29,168,31,132,31,223,31,114,31,94,31,220,31,101,31,101,30,101,29,243,31,165,31,248,31,164,31,10,31,10,30,73,31,172,31,172,30,172,29,99,31,99,30,23,31,228,31,206,31,8,31,8,30,232,31,11,31,62,31,62,30,5,31,5,30,251,31,55,31,204,31,144,31,2,31,2,30,201,31,201,30,139,31,222,31,254,31,97,31,97,30,37,31,57,31,48,31,171,31,171,30,73,31,147,31,95,31,102,31,102,30,63,31,31,31,240,31,53,31,172,31,252,31,30,31,221,31,221,30,234,31,247,31,1,31,139,31,66,31,254,31,254,30,100,31,24,31,24,30,89,31,11,31,146,31,223,31,168,31,124,31,145,31,242,31,103,31,103,30,144,31,228,31,228,30,95,31,95,30,8,31,172,31,55,31,64,31,64,30,15,31,78,31,107,31,147,31,237,31,252,31,124,31,68,31,178,31,36,31,173,31,173,30,160,31,195,31,248,31,248,30,241,31,117,31,117,30,15,31,145,31,145,30,33,31,15,31,15,30,26,31,67,31,255,31,10,31,10,30,10,29,74,31,227,31,93,31,93,30,93,29,181,31,1,31,107,31,153,31,185,31,141,31,125,31,74,31,112,31,31,31,11,31,11,30,26,31,26,30,96,31,133,31,14,31,226,31,226,30,191,31,191,30,164,31,60,31,158,31,161,31,161,30,161,29,161,28,161,27,67,31,18,31,245,31,122,31,199,31,199,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
