-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 502;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (103,0,169,0,92,0,110,0,213,0,62,0,30,0,90,0,73,0,0,0,0,0,97,0,237,0,136,0,31,0,60,0,251,0,95,0,0,0,82,0,150,0,138,0,20,0,90,0,151,0,0,0,159,0,220,0,246,0,64,0,36,0,0,0,0,0,64,0,108,0,113,0,218,0,24,0,245,0,247,0,0,0,144,0,0,0,130,0,175,0,164,0,8,0,11,0,38,0,138,0,0,0,173,0,191,0,99,0,155,0,0,0,75,0,246,0,0,0,190,0,251,0,169,0,145,0,251,0,0,0,175,0,0,0,41,0,32,0,86,0,152,0,57,0,153,0,0,0,207,0,138,0,131,0,251,0,167,0,66,0,235,0,206,0,162,0,84,0,247,0,111,0,53,0,167,0,71,0,104,0,53,0,214,0,107,0,11,0,121,0,76,0,120,0,6,0,44,0,96,0,80,0,187,0,87,0,25,0,26,0,132,0,13,0,240,0,122,0,153,0,101,0,180,0,187,0,236,0,172,0,208,0,0,0,231,0,214,0,0,0,109,0,37,0,221,0,133,0,196,0,0,0,89,0,18,0,46,0,220,0,159,0,161,0,230,0,217,0,0,0,61,0,213,0,15,0,44,0,73,0,209,0,226,0,198,0,35,0,68,0,180,0,0,0,238,0,103,0,55,0,0,0,0,0,209,0,176,0,88,0,120,0,255,0,0,0,238,0,169,0,235,0,88,0,0,0,0,0,0,0,80,0,0,0,0,0,130,0,70,0,131,0,0,0,237,0,54,0,255,0,129,0,246,0,34,0,60,0,42,0,167,0,0,0,0,0,0,0,61,0,0,0,0,0,255,0,0,0,155,0,0,0,0,0,47,0,211,0,14,0,1,0,181,0,32,0,0,0,16,0,3,0,0,0,185,0,32,0,63,0,185,0,53,0,142,0,79,0,125,0,121,0,210,0,0,0,89,0,0,0,59,0,164,0,198,0,233,0,148,0,0,0,138,0,30,0,247,0,216,0,130,0,61,0,38,0,0,0,74,0,145,0,250,0,0,0,197,0,181,0,0,0,182,0,215,0,69,0,85,0,0,0,202,0,0,0,195,0,0,0,225,0,218,0,252,0,0,0,210,0,0,0,161,0,0,0,104,0,203,0,47,0,66,0,234,0,0,0,0,0,0,0,0,0,126,0,171,0,0,0,173,0,67,0,0,0,0,0,88,0,126,0,188,0,0,0,189,0,121,0,130,0,111,0,39,0,37,0,176,0,125,0,101,0,235,0,55,0,251,0,55,0,38,0,83,0,140,0,114,0,210,0,176,0,187,0,0,0,245,0,215,0,18,0,125,0,60,0,11,0,252,0,0,0,252,0,8,0,98,0,241,0,183,0,141,0,0,0,38,0,0,0,194,0,0,0,93,0,9,0,0,0,129,0,17,0,11,0,0,0,0,0,66,0,201,0,0,0,175,0,91,0,31,0,112,0,94,0,252,0,221,0,0,0,14,0,45,0,221,0,226,0,144,0,0,0,227,0,93,0,214,0,153,0,0,0,141,0,0,0,75,0,233,0,214,0,148,0,83,0,0,0,183,0,40,0,93,0,176,0,126,0,39,0,80,0,0,0,39,0,0,0,180,0,6,0,50,0,0,0,37,0,25,0,116,0,7,0,157,0,244,0,242,0,0,0,149,0,8,0,41,0,31,0,0,0,129,0,137,0,195,0,177,0,85,0,150,0,0,0,152,0,217,0,47,0,0,0,173,0,78,0,23,0,93,0,146,0,227,0,252,0,28,0,7,0,51,0,115,0,213,0,214,0,157,0,44,0,253,0,86,0,218,0,0,0,213,0,22,0,0,0,131,0,126,0,0,0,144,0,215,0,75,0,120,0,123,0,0,0,137,0,211,0,141,0,148,0,155,0,138,0,212,0,67,0,111,0,235,0,0,0,67,0,126,0,2,0,1,0,43,0,74,0,0,0,192,0,0,0,85,0,159,0,167,0,232,0,69,0,0,0,29,0,236,0,255,0,213,0,160,0,0,0,6,0,38,0,32,0,0,0,190,0,70,0,105,0,95,0,82,0,182,0,82,0,224,0,0,0,93,0,229,0,77,0,109,0,151,0,0,0,17,0,251,0,192,0,28,0,41,0,142,0,255,0,196,0,148,0,40,0,0,0,194,0,0,0,154,0,190,0,59,0,156,0,88,0,58,0,16,0,205,0,187,0,91,0,215,0,0,0,136,0,0,0,0,0,238,0,210,0,0,0);
signal scenario_full  : scenario_type := (103,31,169,31,92,31,110,31,213,31,62,31,30,31,90,31,73,31,73,30,73,29,97,31,237,31,136,31,31,31,60,31,251,31,95,31,95,30,82,31,150,31,138,31,20,31,90,31,151,31,151,30,159,31,220,31,246,31,64,31,36,31,36,30,36,29,64,31,108,31,113,31,218,31,24,31,245,31,247,31,247,30,144,31,144,30,130,31,175,31,164,31,8,31,11,31,38,31,138,31,138,30,173,31,191,31,99,31,155,31,155,30,75,31,246,31,246,30,190,31,251,31,169,31,145,31,251,31,251,30,175,31,175,30,41,31,32,31,86,31,152,31,57,31,153,31,153,30,207,31,138,31,131,31,251,31,167,31,66,31,235,31,206,31,162,31,84,31,247,31,111,31,53,31,167,31,71,31,104,31,53,31,214,31,107,31,11,31,121,31,76,31,120,31,6,31,44,31,96,31,80,31,187,31,87,31,25,31,26,31,132,31,13,31,240,31,122,31,153,31,101,31,180,31,187,31,236,31,172,31,208,31,208,30,231,31,214,31,214,30,109,31,37,31,221,31,133,31,196,31,196,30,89,31,18,31,46,31,220,31,159,31,161,31,230,31,217,31,217,30,61,31,213,31,15,31,44,31,73,31,209,31,226,31,198,31,35,31,68,31,180,31,180,30,238,31,103,31,55,31,55,30,55,29,209,31,176,31,88,31,120,31,255,31,255,30,238,31,169,31,235,31,88,31,88,30,88,29,88,28,80,31,80,30,80,29,130,31,70,31,131,31,131,30,237,31,54,31,255,31,129,31,246,31,34,31,60,31,42,31,167,31,167,30,167,29,167,28,61,31,61,30,61,29,255,31,255,30,155,31,155,30,155,29,47,31,211,31,14,31,1,31,181,31,32,31,32,30,16,31,3,31,3,30,185,31,32,31,63,31,185,31,53,31,142,31,79,31,125,31,121,31,210,31,210,30,89,31,89,30,59,31,164,31,198,31,233,31,148,31,148,30,138,31,30,31,247,31,216,31,130,31,61,31,38,31,38,30,74,31,145,31,250,31,250,30,197,31,181,31,181,30,182,31,215,31,69,31,85,31,85,30,202,31,202,30,195,31,195,30,225,31,218,31,252,31,252,30,210,31,210,30,161,31,161,30,104,31,203,31,47,31,66,31,234,31,234,30,234,29,234,28,234,27,126,31,171,31,171,30,173,31,67,31,67,30,67,29,88,31,126,31,188,31,188,30,189,31,121,31,130,31,111,31,39,31,37,31,176,31,125,31,101,31,235,31,55,31,251,31,55,31,38,31,83,31,140,31,114,31,210,31,176,31,187,31,187,30,245,31,215,31,18,31,125,31,60,31,11,31,252,31,252,30,252,31,8,31,98,31,241,31,183,31,141,31,141,30,38,31,38,30,194,31,194,30,93,31,9,31,9,30,129,31,17,31,11,31,11,30,11,29,66,31,201,31,201,30,175,31,91,31,31,31,112,31,94,31,252,31,221,31,221,30,14,31,45,31,221,31,226,31,144,31,144,30,227,31,93,31,214,31,153,31,153,30,141,31,141,30,75,31,233,31,214,31,148,31,83,31,83,30,183,31,40,31,93,31,176,31,126,31,39,31,80,31,80,30,39,31,39,30,180,31,6,31,50,31,50,30,37,31,25,31,116,31,7,31,157,31,244,31,242,31,242,30,149,31,8,31,41,31,31,31,31,30,129,31,137,31,195,31,177,31,85,31,150,31,150,30,152,31,217,31,47,31,47,30,173,31,78,31,23,31,93,31,146,31,227,31,252,31,28,31,7,31,51,31,115,31,213,31,214,31,157,31,44,31,253,31,86,31,218,31,218,30,213,31,22,31,22,30,131,31,126,31,126,30,144,31,215,31,75,31,120,31,123,31,123,30,137,31,211,31,141,31,148,31,155,31,138,31,212,31,67,31,111,31,235,31,235,30,67,31,126,31,2,31,1,31,43,31,74,31,74,30,192,31,192,30,85,31,159,31,167,31,232,31,69,31,69,30,29,31,236,31,255,31,213,31,160,31,160,30,6,31,38,31,32,31,32,30,190,31,70,31,105,31,95,31,82,31,182,31,82,31,224,31,224,30,93,31,229,31,77,31,109,31,151,31,151,30,17,31,251,31,192,31,28,31,41,31,142,31,255,31,196,31,148,31,40,31,40,30,194,31,194,30,154,31,190,31,59,31,156,31,88,31,58,31,16,31,205,31,187,31,91,31,215,31,215,30,136,31,136,30,136,29,238,31,210,31,210,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
