-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_851 is
end project_tb_851;

architecture project_tb_arch_851 of project_tb_851 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 796;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (171,0,58,0,161,0,56,0,8,0,77,0,0,0,176,0,21,0,134,0,61,0,222,0,182,0,194,0,9,0,170,0,96,0,143,0,230,0,157,0,38,0,75,0,0,0,0,0,225,0,87,0,0,0,121,0,130,0,166,0,28,0,202,0,27,0,103,0,0,0,229,0,18,0,85,0,113,0,214,0,6,0,62,0,123,0,32,0,138,0,236,0,206,0,33,0,0,0,220,0,176,0,165,0,105,0,247,0,163,0,144,0,76,0,0,0,147,0,252,0,181,0,92,0,230,0,44,0,142,0,44,0,0,0,30,0,0,0,215,0,164,0,249,0,132,0,219,0,0,0,0,0,227,0,61,0,67,0,135,0,137,0,234,0,0,0,142,0,12,0,50,0,179,0,142,0,52,0,190,0,74,0,0,0,60,0,30,0,253,0,249,0,180,0,0,0,91,0,133,0,249,0,185,0,70,0,73,0,241,0,0,0,63,0,131,0,160,0,117,0,99,0,0,0,86,0,145,0,26,0,160,0,74,0,32,0,160,0,233,0,0,0,0,0,0,0,130,0,110,0,119,0,152,0,183,0,73,0,190,0,0,0,209,0,186,0,35,0,245,0,178,0,0,0,0,0,227,0,43,0,0,0,232,0,48,0,135,0,170,0,196,0,0,0,147,0,82,0,154,0,222,0,88,0,49,0,0,0,0,0,87,0,52,0,7,0,0,0,227,0,59,0,72,0,0,0,0,0,240,0,101,0,114,0,148,0,93,0,212,0,3,0,28,0,210,0,35,0,69,0,91,0,95,0,146,0,0,0,219,0,86,0,0,0,46,0,96,0,50,0,80,0,15,0,221,0,168,0,235,0,75,0,20,0,91,0,142,0,0,0,144,0,119,0,220,0,0,0,132,0,255,0,155,0,158,0,0,0,247,0,0,0,251,0,0,0,223,0,250,0,18,0,23,0,37,0,187,0,115,0,118,0,133,0,212,0,72,0,26,0,129,0,0,0,111,0,0,0,59,0,7,0,100,0,0,0,0,0,144,0,47,0,33,0,194,0,90,0,6,0,23,0,31,0,145,0,161,0,102,0,137,0,104,0,28,0,53,0,236,0,67,0,0,0,41,0,90,0,94,0,200,0,0,0,161,0,149,0,140,0,252,0,0,0,182,0,98,0,0,0,182,0,51,0,30,0,88,0,176,0,29,0,58,0,126,0,232,0,68,0,142,0,58,0,0,0,28,0,5,0,74,0,148,0,0,0,211,0,157,0,10,0,0,0,250,0,195,0,31,0,17,0,143,0,67,0,0,0,95,0,219,0,93,0,0,0,179,0,37,0,0,0,234,0,0,0,75,0,84,0,0,0,96,0,0,0,0,0,0,0,196,0,45,0,213,0,15,0,0,0,227,0,60,0,143,0,214,0,18,0,106,0,235,0,138,0,73,0,146,0,201,0,100,0,3,0,237,0,255,0,172,0,151,0,92,0,203,0,17,0,99,0,0,0,209,0,202,0,74,0,221,0,6,0,99,0,61,0,85,0,0,0,14,0,170,0,99,0,29,0,182,0,158,0,89,0,0,0,135,0,65,0,247,0,30,0,0,0,0,0,60,0,96,0,220,0,249,0,159,0,58,0,142,0,159,0,0,0,0,0,101,0,193,0,162,0,0,0,77,0,99,0,0,0,0,0,203,0,0,0,0,0,203,0,89,0,0,0,25,0,245,0,142,0,219,0,0,0,0,0,97,0,117,0,0,0,0,0,140,0,0,0,247,0,0,0,201,0,0,0,219,0,29,0,136,0,70,0,0,0,116,0,139,0,0,0,0,0,38,0,0,0,45,0,57,0,0,0,235,0,192,0,155,0,110,0,0,0,0,0,251,0,133,0,46,0,229,0,34,0,31,0,228,0,99,0,155,0,46,0,252,0,0,0,62,0,110,0,0,0,217,0,84,0,0,0,100,0,171,0,143,0,65,0,71,0,0,0,0,0,251,0,244,0,88,0,244,0,0,0,28,0,152,0,191,0,185,0,2,0,211,0,13,0,89,0,0,0,75,0,250,0,203,0,209,0,216,0,113,0,215,0,105,0,0,0,80,0,72,0,80,0,197,0,82,0,81,0,108,0,120,0,176,0,128,0,0,0,0,0,55,0,58,0,252,0,52,0,22,0,0,0,47,0,149,0,34,0,48,0,250,0,32,0,179,0,0,0,52,0,220,0,0,0,35,0,214,0,25,0,160,0,184,0,71,0,250,0,0,0,89,0,67,0,74,0,208,0,219,0,0,0,65,0,247,0,212,0,0,0,67,0,246,0,161,0,118,0,232,0,220,0,169,0,49,0,235,0,0,0,108,0,24,0,28,0,108,0,131,0,105,0,0,0,77,0,0,0,55,0,141,0,74,0,79,0,181,0,147,0,30,0,240,0,65,0,116,0,216,0,93,0,217,0,200,0,88,0,0,0,0,0,186,0,197,0,107,0,46,0,176,0,0,0,49,0,206,0,0,0,87,0,20,0,94,0,96,0,0,0,0,0,37,0,56,0,32,0,170,0,225,0,223,0,134,0,142,0,178,0,0,0,176,0,10,0,180,0,16,0,138,0,247,0,0,0,123,0,158,0,84,0,116,0,55,0,0,0,250,0,0,0,117,0,181,0,60,0,0,0,4,0,115,0,215,0,69,0,169,0,0,0,221,0,180,0,98,0,0,0,30,0,154,0,82,0,0,0,0,0,81,0,223,0,40,0,111,0,219,0,0,0,83,0,142,0,87,0,32,0,0,0,52,0,1,0,43,0,244,0,73,0,0,0,50,0,0,0,244,0,194,0,187,0,92,0,250,0,234,0,43,0,208,0,72,0,212,0,0,0,233,0,195,0,135,0,112,0,11,0,0,0,110,0,6,0,65,0,80,0,51,0,214,0,0,0,212,0,27,0,147,0,61,0,178,0,48,0,81,0,98,0,138,0,207,0,81,0,43,0,0,0,0,0,247,0,49,0,52,0,26,0,9,0,220,0,203,0,182,0,83,0,83,0,232,0,199,0,59,0,87,0,190,0,162,0,207,0,26,0,0,0,234,0,0,0,77,0,17,0,0,0,136,0,61,0,0,0,214,0,118,0,9,0,6,0,229,0,7,0,45,0,107,0,120,0,231,0,252,0,2,0,128,0,208,0,0,0,126,0,0,0,145,0,0,0,0,0,103,0,0,0,0,0,199,0,0,0,135,0,0,0,233,0,101,0,0,0,0,0,60,0,226,0,108,0,239,0,190,0,77,0,171,0,249,0,169,0,0,0,0,0,65,0,152,0,85,0,243,0,83,0,42,0,0,0,21,0,175,0,208,0,74,0,0,0,106,0,70,0,0,0,181,0,207,0,0,0,160,0,158,0,172,0,35,0,15,0,246,0,169,0,126,0,134,0,158,0,173,0,0,0,244,0,0,0,61,0,97,0,147,0,104,0,0,0,217,0,52,0,77,0,184,0,200,0,238,0,0,0,0,0,231,0,0,0,166,0,128,0,250,0,11,0,232,0,20,0,0,0,29,0,0,0,0,0,177,0,72,0,218,0,50,0,170,0,245,0,43,0,0,0);
signal scenario_full  : scenario_type := (171,31,58,31,161,31,56,31,8,31,77,31,77,30,176,31,21,31,134,31,61,31,222,31,182,31,194,31,9,31,170,31,96,31,143,31,230,31,157,31,38,31,75,31,75,30,75,29,225,31,87,31,87,30,121,31,130,31,166,31,28,31,202,31,27,31,103,31,103,30,229,31,18,31,85,31,113,31,214,31,6,31,62,31,123,31,32,31,138,31,236,31,206,31,33,31,33,30,220,31,176,31,165,31,105,31,247,31,163,31,144,31,76,31,76,30,147,31,252,31,181,31,92,31,230,31,44,31,142,31,44,31,44,30,30,31,30,30,215,31,164,31,249,31,132,31,219,31,219,30,219,29,227,31,61,31,67,31,135,31,137,31,234,31,234,30,142,31,12,31,50,31,179,31,142,31,52,31,190,31,74,31,74,30,60,31,30,31,253,31,249,31,180,31,180,30,91,31,133,31,249,31,185,31,70,31,73,31,241,31,241,30,63,31,131,31,160,31,117,31,99,31,99,30,86,31,145,31,26,31,160,31,74,31,32,31,160,31,233,31,233,30,233,29,233,28,130,31,110,31,119,31,152,31,183,31,73,31,190,31,190,30,209,31,186,31,35,31,245,31,178,31,178,30,178,29,227,31,43,31,43,30,232,31,48,31,135,31,170,31,196,31,196,30,147,31,82,31,154,31,222,31,88,31,49,31,49,30,49,29,87,31,52,31,7,31,7,30,227,31,59,31,72,31,72,30,72,29,240,31,101,31,114,31,148,31,93,31,212,31,3,31,28,31,210,31,35,31,69,31,91,31,95,31,146,31,146,30,219,31,86,31,86,30,46,31,96,31,50,31,80,31,15,31,221,31,168,31,235,31,75,31,20,31,91,31,142,31,142,30,144,31,119,31,220,31,220,30,132,31,255,31,155,31,158,31,158,30,247,31,247,30,251,31,251,30,223,31,250,31,18,31,23,31,37,31,187,31,115,31,118,31,133,31,212,31,72,31,26,31,129,31,129,30,111,31,111,30,59,31,7,31,100,31,100,30,100,29,144,31,47,31,33,31,194,31,90,31,6,31,23,31,31,31,145,31,161,31,102,31,137,31,104,31,28,31,53,31,236,31,67,31,67,30,41,31,90,31,94,31,200,31,200,30,161,31,149,31,140,31,252,31,252,30,182,31,98,31,98,30,182,31,51,31,30,31,88,31,176,31,29,31,58,31,126,31,232,31,68,31,142,31,58,31,58,30,28,31,5,31,74,31,148,31,148,30,211,31,157,31,10,31,10,30,250,31,195,31,31,31,17,31,143,31,67,31,67,30,95,31,219,31,93,31,93,30,179,31,37,31,37,30,234,31,234,30,75,31,84,31,84,30,96,31,96,30,96,29,96,28,196,31,45,31,213,31,15,31,15,30,227,31,60,31,143,31,214,31,18,31,106,31,235,31,138,31,73,31,146,31,201,31,100,31,3,31,237,31,255,31,172,31,151,31,92,31,203,31,17,31,99,31,99,30,209,31,202,31,74,31,221,31,6,31,99,31,61,31,85,31,85,30,14,31,170,31,99,31,29,31,182,31,158,31,89,31,89,30,135,31,65,31,247,31,30,31,30,30,30,29,60,31,96,31,220,31,249,31,159,31,58,31,142,31,159,31,159,30,159,29,101,31,193,31,162,31,162,30,77,31,99,31,99,30,99,29,203,31,203,30,203,29,203,31,89,31,89,30,25,31,245,31,142,31,219,31,219,30,219,29,97,31,117,31,117,30,117,29,140,31,140,30,247,31,247,30,201,31,201,30,219,31,29,31,136,31,70,31,70,30,116,31,139,31,139,30,139,29,38,31,38,30,45,31,57,31,57,30,235,31,192,31,155,31,110,31,110,30,110,29,251,31,133,31,46,31,229,31,34,31,31,31,228,31,99,31,155,31,46,31,252,31,252,30,62,31,110,31,110,30,217,31,84,31,84,30,100,31,171,31,143,31,65,31,71,31,71,30,71,29,251,31,244,31,88,31,244,31,244,30,28,31,152,31,191,31,185,31,2,31,211,31,13,31,89,31,89,30,75,31,250,31,203,31,209,31,216,31,113,31,215,31,105,31,105,30,80,31,72,31,80,31,197,31,82,31,81,31,108,31,120,31,176,31,128,31,128,30,128,29,55,31,58,31,252,31,52,31,22,31,22,30,47,31,149,31,34,31,48,31,250,31,32,31,179,31,179,30,52,31,220,31,220,30,35,31,214,31,25,31,160,31,184,31,71,31,250,31,250,30,89,31,67,31,74,31,208,31,219,31,219,30,65,31,247,31,212,31,212,30,67,31,246,31,161,31,118,31,232,31,220,31,169,31,49,31,235,31,235,30,108,31,24,31,28,31,108,31,131,31,105,31,105,30,77,31,77,30,55,31,141,31,74,31,79,31,181,31,147,31,30,31,240,31,65,31,116,31,216,31,93,31,217,31,200,31,88,31,88,30,88,29,186,31,197,31,107,31,46,31,176,31,176,30,49,31,206,31,206,30,87,31,20,31,94,31,96,31,96,30,96,29,37,31,56,31,32,31,170,31,225,31,223,31,134,31,142,31,178,31,178,30,176,31,10,31,180,31,16,31,138,31,247,31,247,30,123,31,158,31,84,31,116,31,55,31,55,30,250,31,250,30,117,31,181,31,60,31,60,30,4,31,115,31,215,31,69,31,169,31,169,30,221,31,180,31,98,31,98,30,30,31,154,31,82,31,82,30,82,29,81,31,223,31,40,31,111,31,219,31,219,30,83,31,142,31,87,31,32,31,32,30,52,31,1,31,43,31,244,31,73,31,73,30,50,31,50,30,244,31,194,31,187,31,92,31,250,31,234,31,43,31,208,31,72,31,212,31,212,30,233,31,195,31,135,31,112,31,11,31,11,30,110,31,6,31,65,31,80,31,51,31,214,31,214,30,212,31,27,31,147,31,61,31,178,31,48,31,81,31,98,31,138,31,207,31,81,31,43,31,43,30,43,29,247,31,49,31,52,31,26,31,9,31,220,31,203,31,182,31,83,31,83,31,232,31,199,31,59,31,87,31,190,31,162,31,207,31,26,31,26,30,234,31,234,30,77,31,17,31,17,30,136,31,61,31,61,30,214,31,118,31,9,31,6,31,229,31,7,31,45,31,107,31,120,31,231,31,252,31,2,31,128,31,208,31,208,30,126,31,126,30,145,31,145,30,145,29,103,31,103,30,103,29,199,31,199,30,135,31,135,30,233,31,101,31,101,30,101,29,60,31,226,31,108,31,239,31,190,31,77,31,171,31,249,31,169,31,169,30,169,29,65,31,152,31,85,31,243,31,83,31,42,31,42,30,21,31,175,31,208,31,74,31,74,30,106,31,70,31,70,30,181,31,207,31,207,30,160,31,158,31,172,31,35,31,15,31,246,31,169,31,126,31,134,31,158,31,173,31,173,30,244,31,244,30,61,31,97,31,147,31,104,31,104,30,217,31,52,31,77,31,184,31,200,31,238,31,238,30,238,29,231,31,231,30,166,31,128,31,250,31,11,31,232,31,20,31,20,30,29,31,29,30,29,29,177,31,72,31,218,31,50,31,170,31,245,31,43,31,43,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
