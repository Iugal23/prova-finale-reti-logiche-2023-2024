-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 623;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (18,0,31,0,165,0,248,0,0,0,0,0,46,0,52,0,197,0,145,0,150,0,51,0,90,0,103,0,187,0,158,0,216,0,137,0,26,0,10,0,56,0,0,0,0,0,244,0,208,0,71,0,94,0,51,0,0,0,169,0,33,0,212,0,0,0,23,0,10,0,143,0,117,0,95,0,186,0,252,0,0,0,200,0,49,0,0,0,97,0,8,0,97,0,0,0,180,0,0,0,205,0,107,0,142,0,156,0,167,0,39,0,126,0,32,0,0,0,0,0,172,0,0,0,208,0,146,0,0,0,0,0,247,0,176,0,197,0,175,0,197,0,0,0,97,0,95,0,218,0,0,0,0,0,9,0,16,0,2,0,142,0,221,0,98,0,120,0,208,0,82,0,18,0,235,0,0,0,65,0,0,0,253,0,160,0,106,0,122,0,0,0,251,0,37,0,145,0,162,0,189,0,0,0,133,0,225,0,83,0,238,0,46,0,2,0,116,0,137,0,0,0,126,0,210,0,140,0,223,0,160,0,0,0,205,0,212,0,191,0,170,0,150,0,76,0,123,0,193,0,138,0,185,0,102,0,43,0,0,0,123,0,0,0,198,0,8,0,119,0,0,0,154,0,23,0,0,0,153,0,228,0,0,0,3,0,57,0,33,0,19,0,234,0,185,0,83,0,24,0,4,0,95,0,12,0,46,0,244,0,124,0,7,0,138,0,117,0,70,0,0,0,58,0,107,0,150,0,0,0,60,0,230,0,0,0,157,0,175,0,51,0,169,0,0,0,7,0,180,0,13,0,78,0,120,0,0,0,203,0,0,0,216,0,169,0,0,0,0,0,144,0,167,0,58,0,113,0,0,0,125,0,216,0,191,0,18,0,65,0,215,0,0,0,101,0,75,0,88,0,158,0,0,0,167,0,136,0,133,0,57,0,0,0,110,0,0,0,49,0,158,0,0,0,233,0,198,0,23,0,1,0,211,0,110,0,40,0,147,0,171,0,181,0,123,0,167,0,0,0,0,0,76,0,88,0,237,0,221,0,79,0,132,0,36,0,32,0,0,0,1,0,52,0,82,0,0,0,214,0,227,0,182,0,112,0,224,0,142,0,48,0,0,0,164,0,48,0,156,0,174,0,58,0,0,0,238,0,225,0,175,0,117,0,29,0,0,0,35,0,231,0,5,0,77,0,0,0,0,0,39,0,50,0,118,0,72,0,201,0,90,0,128,0,122,0,104,0,195,0,71,0,70,0,0,0,196,0,166,0,143,0,169,0,220,0,250,0,0,0,14,0,0,0,71,0,221,0,32,0,179,0,119,0,0,0,104,0,35,0,138,0,244,0,199,0,58,0,241,0,55,0,0,0,0,0,50,0,137,0,201,0,0,0,0,0,0,0,62,0,94,0,217,0,179,0,14,0,191,0,244,0,222,0,144,0,15,0,131,0,0,0,109,0,0,0,152,0,196,0,52,0,0,0,228,0,194,0,34,0,80,0,105,0,0,0,243,0,20,0,61,0,224,0,135,0,185,0,59,0,79,0,0,0,213,0,149,0,241,0,223,0,120,0,97,0,200,0,233,0,0,0,227,0,236,0,28,0,74,0,108,0,63,0,71,0,107,0,69,0,0,0,56,0,217,0,81,0,86,0,51,0,138,0,172,0,213,0,183,0,206,0,22,0,93,0,140,0,29,0,108,0,148,0,157,0,0,0,211,0,182,0,222,0,80,0,251,0,34,0,108,0,33,0,79,0,203,0,240,0,12,0,27,0,188,0,94,0,143,0,47,0,140,0,161,0,79,0,23,0,167,0,0,0,195,0,5,0,24,0,33,0,45,0,217,0,194,0,138,0,236,0,109,0,201,0,7,0,187,0,0,0,98,0,0,0,90,0,145,0,0,0,47,0,210,0,161,0,13,0,210,0,0,0,116,0,156,0,114,0,177,0,201,0,62,0,204,0,16,0,78,0,0,0,56,0,42,0,0,0,48,0,64,0,112,0,87,0,155,0,0,0,191,0,216,0,192,0,0,0,75,0,184,0,83,0,205,0,44,0,94,0,171,0,33,0,17,0,0,0,109,0,99,0,237,0,191,0,237,0,52,0,194,0,0,0,0,0,0,0,195,0,32,0,67,0,0,0,0,0,114,0,144,0,21,0,60,0,216,0,255,0,60,0,0,0,0,0,30,0,0,0,0,0,128,0,223,0,143,0,0,0,23,0,229,0,92,0,161,0,215,0,253,0,0,0,191,0,54,0,0,0,194,0,146,0,0,0,25,0,0,0,53,0,0,0,0,0,0,0,13,0,171,0,71,0,0,0,0,0,151,0,83,0,88,0,234,0,0,0,17,0,86,0,200,0,90,0,185,0,223,0,234,0,6,0,71,0,0,0,174,0,182,0,136,0,0,0,0,0,0,0,0,0,136,0,99,0,45,0,0,0,197,0,223,0,254,0,0,0,176,0,0,0,158,0,0,0,92,0,144,0,0,0,167,0,78,0,0,0,120,0,85,0,10,0,97,0,122,0,186,0,127,0,164,0,225,0,125,0,0,0,0,0,164,0,189,0,68,0,54,0,146,0,0,0,39,0,100,0,247,0,42,0,48,0,55,0,197,0,175,0,203,0,151,0,0,0,188,0,63,0,0,0,152,0,0,0,27,0,0,0,146,0,0,0,122,0,121,0,16,0,206,0,0,0,209,0,117,0,222,0,145,0,182,0,0,0,11,0,102,0,0,0,26,0,25,0,0,0,130,0,140,0,99,0,162,0,0,0,98,0,219,0,210,0,49,0,119,0,186,0,189,0,47,0);
signal scenario_full  : scenario_type := (18,31,31,31,165,31,248,31,248,30,248,29,46,31,52,31,197,31,145,31,150,31,51,31,90,31,103,31,187,31,158,31,216,31,137,31,26,31,10,31,56,31,56,30,56,29,244,31,208,31,71,31,94,31,51,31,51,30,169,31,33,31,212,31,212,30,23,31,10,31,143,31,117,31,95,31,186,31,252,31,252,30,200,31,49,31,49,30,97,31,8,31,97,31,97,30,180,31,180,30,205,31,107,31,142,31,156,31,167,31,39,31,126,31,32,31,32,30,32,29,172,31,172,30,208,31,146,31,146,30,146,29,247,31,176,31,197,31,175,31,197,31,197,30,97,31,95,31,218,31,218,30,218,29,9,31,16,31,2,31,142,31,221,31,98,31,120,31,208,31,82,31,18,31,235,31,235,30,65,31,65,30,253,31,160,31,106,31,122,31,122,30,251,31,37,31,145,31,162,31,189,31,189,30,133,31,225,31,83,31,238,31,46,31,2,31,116,31,137,31,137,30,126,31,210,31,140,31,223,31,160,31,160,30,205,31,212,31,191,31,170,31,150,31,76,31,123,31,193,31,138,31,185,31,102,31,43,31,43,30,123,31,123,30,198,31,8,31,119,31,119,30,154,31,23,31,23,30,153,31,228,31,228,30,3,31,57,31,33,31,19,31,234,31,185,31,83,31,24,31,4,31,95,31,12,31,46,31,244,31,124,31,7,31,138,31,117,31,70,31,70,30,58,31,107,31,150,31,150,30,60,31,230,31,230,30,157,31,175,31,51,31,169,31,169,30,7,31,180,31,13,31,78,31,120,31,120,30,203,31,203,30,216,31,169,31,169,30,169,29,144,31,167,31,58,31,113,31,113,30,125,31,216,31,191,31,18,31,65,31,215,31,215,30,101,31,75,31,88,31,158,31,158,30,167,31,136,31,133,31,57,31,57,30,110,31,110,30,49,31,158,31,158,30,233,31,198,31,23,31,1,31,211,31,110,31,40,31,147,31,171,31,181,31,123,31,167,31,167,30,167,29,76,31,88,31,237,31,221,31,79,31,132,31,36,31,32,31,32,30,1,31,52,31,82,31,82,30,214,31,227,31,182,31,112,31,224,31,142,31,48,31,48,30,164,31,48,31,156,31,174,31,58,31,58,30,238,31,225,31,175,31,117,31,29,31,29,30,35,31,231,31,5,31,77,31,77,30,77,29,39,31,50,31,118,31,72,31,201,31,90,31,128,31,122,31,104,31,195,31,71,31,70,31,70,30,196,31,166,31,143,31,169,31,220,31,250,31,250,30,14,31,14,30,71,31,221,31,32,31,179,31,119,31,119,30,104,31,35,31,138,31,244,31,199,31,58,31,241,31,55,31,55,30,55,29,50,31,137,31,201,31,201,30,201,29,201,28,62,31,94,31,217,31,179,31,14,31,191,31,244,31,222,31,144,31,15,31,131,31,131,30,109,31,109,30,152,31,196,31,52,31,52,30,228,31,194,31,34,31,80,31,105,31,105,30,243,31,20,31,61,31,224,31,135,31,185,31,59,31,79,31,79,30,213,31,149,31,241,31,223,31,120,31,97,31,200,31,233,31,233,30,227,31,236,31,28,31,74,31,108,31,63,31,71,31,107,31,69,31,69,30,56,31,217,31,81,31,86,31,51,31,138,31,172,31,213,31,183,31,206,31,22,31,93,31,140,31,29,31,108,31,148,31,157,31,157,30,211,31,182,31,222,31,80,31,251,31,34,31,108,31,33,31,79,31,203,31,240,31,12,31,27,31,188,31,94,31,143,31,47,31,140,31,161,31,79,31,23,31,167,31,167,30,195,31,5,31,24,31,33,31,45,31,217,31,194,31,138,31,236,31,109,31,201,31,7,31,187,31,187,30,98,31,98,30,90,31,145,31,145,30,47,31,210,31,161,31,13,31,210,31,210,30,116,31,156,31,114,31,177,31,201,31,62,31,204,31,16,31,78,31,78,30,56,31,42,31,42,30,48,31,64,31,112,31,87,31,155,31,155,30,191,31,216,31,192,31,192,30,75,31,184,31,83,31,205,31,44,31,94,31,171,31,33,31,17,31,17,30,109,31,99,31,237,31,191,31,237,31,52,31,194,31,194,30,194,29,194,28,195,31,32,31,67,31,67,30,67,29,114,31,144,31,21,31,60,31,216,31,255,31,60,31,60,30,60,29,30,31,30,30,30,29,128,31,223,31,143,31,143,30,23,31,229,31,92,31,161,31,215,31,253,31,253,30,191,31,54,31,54,30,194,31,146,31,146,30,25,31,25,30,53,31,53,30,53,29,53,28,13,31,171,31,71,31,71,30,71,29,151,31,83,31,88,31,234,31,234,30,17,31,86,31,200,31,90,31,185,31,223,31,234,31,6,31,71,31,71,30,174,31,182,31,136,31,136,30,136,29,136,28,136,27,136,31,99,31,45,31,45,30,197,31,223,31,254,31,254,30,176,31,176,30,158,31,158,30,92,31,144,31,144,30,167,31,78,31,78,30,120,31,85,31,10,31,97,31,122,31,186,31,127,31,164,31,225,31,125,31,125,30,125,29,164,31,189,31,68,31,54,31,146,31,146,30,39,31,100,31,247,31,42,31,48,31,55,31,197,31,175,31,203,31,151,31,151,30,188,31,63,31,63,30,152,31,152,30,27,31,27,30,146,31,146,30,122,31,121,31,16,31,206,31,206,30,209,31,117,31,222,31,145,31,182,31,182,30,11,31,102,31,102,30,26,31,25,31,25,30,130,31,140,31,99,31,162,31,162,30,98,31,219,31,210,31,49,31,119,31,186,31,189,31,47,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
