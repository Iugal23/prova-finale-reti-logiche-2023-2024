-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 954;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (93,0,0,0,0,0,46,0,104,0,47,0,0,0,63,0,11,0,210,0,225,0,163,0,150,0,203,0,156,0,234,0,0,0,159,0,54,0,187,0,0,0,223,0,226,0,193,0,201,0,177,0,233,0,119,0,56,0,87,0,178,0,124,0,189,0,206,0,149,0,118,0,0,0,170,0,249,0,218,0,0,0,210,0,0,0,0,0,133,0,0,0,150,0,0,0,71,0,57,0,236,0,93,0,129,0,127,0,205,0,78,0,99,0,0,0,81,0,203,0,229,0,201,0,148,0,0,0,36,0,75,0,156,0,0,0,255,0,87,0,1,0,186,0,14,0,175,0,45,0,47,0,169,0,234,0,0,0,161,0,234,0,129,0,120,0,0,0,13,0,177,0,30,0,236,0,29,0,0,0,24,0,141,0,0,0,0,0,0,0,186,0,121,0,0,0,143,0,0,0,189,0,18,0,226,0,0,0,0,0,37,0,12,0,187,0,246,0,74,0,209,0,100,0,206,0,61,0,99,0,13,0,0,0,153,0,15,0,0,0,81,0,18,0,146,0,28,0,0,0,0,0,12,0,52,0,39,0,237,0,238,0,37,0,152,0,21,0,38,0,41,0,0,0,0,0,44,0,140,0,129,0,242,0,152,0,83,0,89,0,115,0,169,0,65,0,223,0,0,0,255,0,245,0,205,0,136,0,0,0,0,0,102,0,68,0,30,0,130,0,95,0,29,0,137,0,16,0,173,0,247,0,193,0,0,0,9,0,241,0,166,0,0,0,154,0,144,0,149,0,185,0,177,0,0,0,6,0,130,0,243,0,0,0,243,0,0,0,0,0,134,0,209,0,85,0,202,0,149,0,0,0,240,0,60,0,161,0,121,0,4,0,16,0,138,0,78,0,0,0,252,0,83,0,117,0,130,0,0,0,0,0,230,0,0,0,252,0,137,0,198,0,9,0,13,0,179,0,0,0,82,0,88,0,0,0,85,0,235,0,109,0,80,0,209,0,0,0,3,0,132,0,7,0,46,0,43,0,69,0,214,0,109,0,238,0,24,0,10,0,165,0,41,0,167,0,0,0,211,0,35,0,62,0,185,0,50,0,129,0,31,0,105,0,151,0,101,0,222,0,146,0,168,0,0,0,70,0,75,0,102,0,0,0,16,0,0,0,124,0,5,0,190,0,224,0,6,0,223,0,217,0,227,0,144,0,0,0,0,0,12,0,10,0,233,0,88,0,18,0,2,0,94,0,109,0,86,0,230,0,158,0,39,0,205,0,98,0,0,0,70,0,0,0,0,0,29,0,88,0,0,0,114,0,0,0,227,0,0,0,236,0,21,0,40,0,28,0,8,0,134,0,94,0,218,0,227,0,11,0,159,0,121,0,224,0,197,0,0,0,0,0,109,0,0,0,232,0,242,0,148,0,0,0,68,0,157,0,230,0,177,0,0,0,253,0,71,0,83,0,120,0,146,0,23,0,44,0,97,0,146,0,0,0,242,0,144,0,119,0,190,0,102,0,182,0,197,0,228,0,35,0,162,0,163,0,251,0,24,0,0,0,22,0,241,0,0,0,252,0,9,0,186,0,193,0,190,0,195,0,77,0,218,0,206,0,76,0,34,0,201,0,0,0,73,0,175,0,45,0,158,0,0,0,78,0,249,0,73,0,169,0,141,0,70,0,91,0,231,0,0,0,0,0,168,0,125,0,139,0,182,0,6,0,37,0,93,0,78,0,0,0,0,0,159,0,40,0,221,0,130,0,170,0,190,0,194,0,200,0,212,0,232,0,124,0,0,0,177,0,226,0,0,0,0,0,116,0,0,0,115,0,0,0,33,0,126,0,115,0,209,0,77,0,217,0,59,0,185,0,0,0,88,0,0,0,0,0,95,0,0,0,111,0,92,0,71,0,43,0,42,0,0,0,173,0,84,0,164,0,118,0,0,0,38,0,243,0,249,0,0,0,0,0,101,0,30,0,0,0,161,0,202,0,0,0,56,0,169,0,127,0,155,0,173,0,78,0,36,0,87,0,66,0,129,0,39,0,0,0,77,0,21,0,202,0,0,0,64,0,49,0,98,0,159,0,0,0,56,0,30,0,88,0,182,0,109,0,173,0,207,0,60,0,150,0,197,0,142,0,200,0,135,0,173,0,171,0,0,0,0,0,127,0,108,0,158,0,97,0,0,0,0,0,227,0,21,0,240,0,73,0,0,0,96,0,140,0,0,0,0,0,0,0,0,0,65,0,0,0,0,0,255,0,129,0,126,0,222,0,166,0,161,0,22,0,25,0,2,0,75,0,55,0,231,0,86,0,7,0,0,0,128,0,105,0,203,0,205,0,1,0,100,0,44,0,0,0,37,0,43,0,42,0,108,0,176,0,95,0,61,0,1,0,91,0,161,0,16,0,4,0,210,0,252,0,0,0,107,0,74,0,50,0,250,0,109,0,0,0,0,0,0,0,92,0,106,0,99,0,112,0,0,0,0,0,115,0,0,0,33,0,140,0,64,0,97,0,60,0,0,0,22,0,172,0,56,0,118,0,14,0,11,0,111,0,30,0,0,0,98,0,201,0,181,0,0,0,76,0,95,0,113,0,214,0,150,0,0,0,156,0,192,0,229,0,5,0,112,0,211,0,133,0,77,0,0,0,231,0,214,0,82,0,0,0,53,0,166,0,0,0,86,0,253,0,25,0,108,0,170,0,130,0,58,0,102,0,134,0,0,0,49,0,0,0,237,0,190,0,86,0,39,0,173,0,67,0,41,0,136,0,117,0,237,0,175,0,100,0,92,0,183,0,0,0,0,0,132,0,67,0,0,0,213,0,78,0,0,0,32,0,0,0,33,0,0,0,194,0,176,0,0,0,137,0,0,0,158,0,0,0,80,0,0,0,43,0,0,0,190,0,214,0,74,0,0,0,137,0,0,0,0,0,235,0,162,0,184,0,254,0,0,0,197,0,142,0,99,0,132,0,119,0,54,0,239,0,226,0,9,0,25,0,165,0,79,0,221,0,248,0,23,0,0,0,66,0,9,0,253,0,0,0,193,0,0,0,190,0,0,0,29,0,112,0,0,0,73,0,122,0,169,0,197,0,0,0,0,0,187,0,133,0,63,0,174,0,108,0,181,0,130,0,224,0,251,0,190,0,0,0,127,0,35,0,0,0,232,0,105,0,0,0,250,0,131,0,159,0,79,0,253,0,186,0,0,0,121,0,77,0,90,0,89,0,63,0,184,0,112,0,37,0,244,0,154,0,0,0,243,0,111,0,89,0,0,0,0,0,100,0,0,0,221,0,212,0,240,0,221,0,230,0,0,0,248,0,141,0,194,0,234,0,82,0,0,0,0,0,116,0,59,0,0,0,160,0,11,0,18,0,22,0,27,0,108,0,0,0,166,0,45,0,187,0,146,0,91,0,16,0,53,0,26,0,13,0,89,0,43,0,4,0,226,0,19,0,104,0,0,0,4,0,225,0,0,0,107,0,74,0,0,0,213,0,0,0,66,0,203,0,108,0,48,0,0,0,157,0,9,0,26,0,0,0,0,0,181,0,249,0,3,0,0,0,204,0,231,0,0,0,91,0,230,0,112,0,173,0,0,0,31,0,232,0,25,0,0,0,40,0,0,0,98,0,34,0,88,0,4,0,138,0,53,0,0,0,172,0,211,0,76,0,142,0,132,0,196,0,184,0,184,0,0,0,86,0,0,0,164,0,1,0,77,0,131,0,218,0,170,0,57,0,90,0,82,0,163,0,173,0,102,0,179,0,135,0,225,0,91,0,70,0,116,0,250,0,91,0,25,0,252,0,0,0,31,0,0,0,0,0,148,0,17,0,34,0,101,0,214,0,102,0,146,0,0,0,73,0,0,0,0,0,28,0,222,0,0,0,109,0,64,0,98,0,207,0,253,0,41,0,68,0,162,0,0,0,137,0,10,0,183,0,130,0,161,0,184,0,126,0,117,0,107,0,174,0,134,0,109,0,248,0,136,0,144,0,115,0,159,0,97,0,80,0,0,0,198,0,129,0,184,0,36,0,242,0,184,0,79,0,0,0,103,0,0,0,1,0,107,0,0,0,75,0,42,0,0,0,26,0,180,0,125,0,12,0,54,0,218,0,0,0,0,0,155,0,0,0,148,0,163,0,44,0,107,0,0,0,0,0,238,0,146,0,77,0,180,0,90,0,201,0,0,0,59,0,7,0,218,0,0,0,0,0,253,0,101,0,195,0,64,0,130,0,0,0,0,0,0,0,203,0,253,0,114,0,0,0,192,0,0,0,63,0,0,0);
signal scenario_full  : scenario_type := (93,31,93,30,93,29,46,31,104,31,47,31,47,30,63,31,11,31,210,31,225,31,163,31,150,31,203,31,156,31,234,31,234,30,159,31,54,31,187,31,187,30,223,31,226,31,193,31,201,31,177,31,233,31,119,31,56,31,87,31,178,31,124,31,189,31,206,31,149,31,118,31,118,30,170,31,249,31,218,31,218,30,210,31,210,30,210,29,133,31,133,30,150,31,150,30,71,31,57,31,236,31,93,31,129,31,127,31,205,31,78,31,99,31,99,30,81,31,203,31,229,31,201,31,148,31,148,30,36,31,75,31,156,31,156,30,255,31,87,31,1,31,186,31,14,31,175,31,45,31,47,31,169,31,234,31,234,30,161,31,234,31,129,31,120,31,120,30,13,31,177,31,30,31,236,31,29,31,29,30,24,31,141,31,141,30,141,29,141,28,186,31,121,31,121,30,143,31,143,30,189,31,18,31,226,31,226,30,226,29,37,31,12,31,187,31,246,31,74,31,209,31,100,31,206,31,61,31,99,31,13,31,13,30,153,31,15,31,15,30,81,31,18,31,146,31,28,31,28,30,28,29,12,31,52,31,39,31,237,31,238,31,37,31,152,31,21,31,38,31,41,31,41,30,41,29,44,31,140,31,129,31,242,31,152,31,83,31,89,31,115,31,169,31,65,31,223,31,223,30,255,31,245,31,205,31,136,31,136,30,136,29,102,31,68,31,30,31,130,31,95,31,29,31,137,31,16,31,173,31,247,31,193,31,193,30,9,31,241,31,166,31,166,30,154,31,144,31,149,31,185,31,177,31,177,30,6,31,130,31,243,31,243,30,243,31,243,30,243,29,134,31,209,31,85,31,202,31,149,31,149,30,240,31,60,31,161,31,121,31,4,31,16,31,138,31,78,31,78,30,252,31,83,31,117,31,130,31,130,30,130,29,230,31,230,30,252,31,137,31,198,31,9,31,13,31,179,31,179,30,82,31,88,31,88,30,85,31,235,31,109,31,80,31,209,31,209,30,3,31,132,31,7,31,46,31,43,31,69,31,214,31,109,31,238,31,24,31,10,31,165,31,41,31,167,31,167,30,211,31,35,31,62,31,185,31,50,31,129,31,31,31,105,31,151,31,101,31,222,31,146,31,168,31,168,30,70,31,75,31,102,31,102,30,16,31,16,30,124,31,5,31,190,31,224,31,6,31,223,31,217,31,227,31,144,31,144,30,144,29,12,31,10,31,233,31,88,31,18,31,2,31,94,31,109,31,86,31,230,31,158,31,39,31,205,31,98,31,98,30,70,31,70,30,70,29,29,31,88,31,88,30,114,31,114,30,227,31,227,30,236,31,21,31,40,31,28,31,8,31,134,31,94,31,218,31,227,31,11,31,159,31,121,31,224,31,197,31,197,30,197,29,109,31,109,30,232,31,242,31,148,31,148,30,68,31,157,31,230,31,177,31,177,30,253,31,71,31,83,31,120,31,146,31,23,31,44,31,97,31,146,31,146,30,242,31,144,31,119,31,190,31,102,31,182,31,197,31,228,31,35,31,162,31,163,31,251,31,24,31,24,30,22,31,241,31,241,30,252,31,9,31,186,31,193,31,190,31,195,31,77,31,218,31,206,31,76,31,34,31,201,31,201,30,73,31,175,31,45,31,158,31,158,30,78,31,249,31,73,31,169,31,141,31,70,31,91,31,231,31,231,30,231,29,168,31,125,31,139,31,182,31,6,31,37,31,93,31,78,31,78,30,78,29,159,31,40,31,221,31,130,31,170,31,190,31,194,31,200,31,212,31,232,31,124,31,124,30,177,31,226,31,226,30,226,29,116,31,116,30,115,31,115,30,33,31,126,31,115,31,209,31,77,31,217,31,59,31,185,31,185,30,88,31,88,30,88,29,95,31,95,30,111,31,92,31,71,31,43,31,42,31,42,30,173,31,84,31,164,31,118,31,118,30,38,31,243,31,249,31,249,30,249,29,101,31,30,31,30,30,161,31,202,31,202,30,56,31,169,31,127,31,155,31,173,31,78,31,36,31,87,31,66,31,129,31,39,31,39,30,77,31,21,31,202,31,202,30,64,31,49,31,98,31,159,31,159,30,56,31,30,31,88,31,182,31,109,31,173,31,207,31,60,31,150,31,197,31,142,31,200,31,135,31,173,31,171,31,171,30,171,29,127,31,108,31,158,31,97,31,97,30,97,29,227,31,21,31,240,31,73,31,73,30,96,31,140,31,140,30,140,29,140,28,140,27,65,31,65,30,65,29,255,31,129,31,126,31,222,31,166,31,161,31,22,31,25,31,2,31,75,31,55,31,231,31,86,31,7,31,7,30,128,31,105,31,203,31,205,31,1,31,100,31,44,31,44,30,37,31,43,31,42,31,108,31,176,31,95,31,61,31,1,31,91,31,161,31,16,31,4,31,210,31,252,31,252,30,107,31,74,31,50,31,250,31,109,31,109,30,109,29,109,28,92,31,106,31,99,31,112,31,112,30,112,29,115,31,115,30,33,31,140,31,64,31,97,31,60,31,60,30,22,31,172,31,56,31,118,31,14,31,11,31,111,31,30,31,30,30,98,31,201,31,181,31,181,30,76,31,95,31,113,31,214,31,150,31,150,30,156,31,192,31,229,31,5,31,112,31,211,31,133,31,77,31,77,30,231,31,214,31,82,31,82,30,53,31,166,31,166,30,86,31,253,31,25,31,108,31,170,31,130,31,58,31,102,31,134,31,134,30,49,31,49,30,237,31,190,31,86,31,39,31,173,31,67,31,41,31,136,31,117,31,237,31,175,31,100,31,92,31,183,31,183,30,183,29,132,31,67,31,67,30,213,31,78,31,78,30,32,31,32,30,33,31,33,30,194,31,176,31,176,30,137,31,137,30,158,31,158,30,80,31,80,30,43,31,43,30,190,31,214,31,74,31,74,30,137,31,137,30,137,29,235,31,162,31,184,31,254,31,254,30,197,31,142,31,99,31,132,31,119,31,54,31,239,31,226,31,9,31,25,31,165,31,79,31,221,31,248,31,23,31,23,30,66,31,9,31,253,31,253,30,193,31,193,30,190,31,190,30,29,31,112,31,112,30,73,31,122,31,169,31,197,31,197,30,197,29,187,31,133,31,63,31,174,31,108,31,181,31,130,31,224,31,251,31,190,31,190,30,127,31,35,31,35,30,232,31,105,31,105,30,250,31,131,31,159,31,79,31,253,31,186,31,186,30,121,31,77,31,90,31,89,31,63,31,184,31,112,31,37,31,244,31,154,31,154,30,243,31,111,31,89,31,89,30,89,29,100,31,100,30,221,31,212,31,240,31,221,31,230,31,230,30,248,31,141,31,194,31,234,31,82,31,82,30,82,29,116,31,59,31,59,30,160,31,11,31,18,31,22,31,27,31,108,31,108,30,166,31,45,31,187,31,146,31,91,31,16,31,53,31,26,31,13,31,89,31,43,31,4,31,226,31,19,31,104,31,104,30,4,31,225,31,225,30,107,31,74,31,74,30,213,31,213,30,66,31,203,31,108,31,48,31,48,30,157,31,9,31,26,31,26,30,26,29,181,31,249,31,3,31,3,30,204,31,231,31,231,30,91,31,230,31,112,31,173,31,173,30,31,31,232,31,25,31,25,30,40,31,40,30,98,31,34,31,88,31,4,31,138,31,53,31,53,30,172,31,211,31,76,31,142,31,132,31,196,31,184,31,184,31,184,30,86,31,86,30,164,31,1,31,77,31,131,31,218,31,170,31,57,31,90,31,82,31,163,31,173,31,102,31,179,31,135,31,225,31,91,31,70,31,116,31,250,31,91,31,25,31,252,31,252,30,31,31,31,30,31,29,148,31,17,31,34,31,101,31,214,31,102,31,146,31,146,30,73,31,73,30,73,29,28,31,222,31,222,30,109,31,64,31,98,31,207,31,253,31,41,31,68,31,162,31,162,30,137,31,10,31,183,31,130,31,161,31,184,31,126,31,117,31,107,31,174,31,134,31,109,31,248,31,136,31,144,31,115,31,159,31,97,31,80,31,80,30,198,31,129,31,184,31,36,31,242,31,184,31,79,31,79,30,103,31,103,30,1,31,107,31,107,30,75,31,42,31,42,30,26,31,180,31,125,31,12,31,54,31,218,31,218,30,218,29,155,31,155,30,148,31,163,31,44,31,107,31,107,30,107,29,238,31,146,31,77,31,180,31,90,31,201,31,201,30,59,31,7,31,218,31,218,30,218,29,253,31,101,31,195,31,64,31,130,31,130,30,130,29,130,28,203,31,253,31,114,31,114,30,192,31,192,30,63,31,63,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
