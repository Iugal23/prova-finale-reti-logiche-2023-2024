-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_994 is
end project_tb_994;

architecture project_tb_arch_994 of project_tb_994 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 388;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (206,0,254,0,247,0,99,0,37,0,104,0,6,0,199,0,181,0,103,0,102,0,216,0,23,0,255,0,190,0,182,0,0,0,169,0,102,0,233,0,0,0,66,0,0,0,122,0,206,0,182,0,19,0,235,0,221,0,101,0,121,0,215,0,231,0,0,0,10,0,126,0,247,0,188,0,112,0,180,0,0,0,154,0,154,0,121,0,38,0,167,0,248,0,0,0,0,0,49,0,139,0,232,0,241,0,34,0,218,0,37,0,142,0,216,0,0,0,216,0,0,0,240,0,153,0,124,0,213,0,134,0,204,0,0,0,0,0,97,0,218,0,189,0,232,0,198,0,14,0,134,0,106,0,147,0,189,0,4,0,252,0,221,0,57,0,217,0,188,0,180,0,248,0,222,0,16,0,70,0,47,0,140,0,170,0,0,0,129,0,142,0,0,0,0,0,10,0,172,0,226,0,236,0,11,0,39,0,160,0,0,0,19,0,191,0,119,0,66,0,35,0,1,0,42,0,171,0,55,0,0,0,69,0,110,0,199,0,33,0,115,0,184,0,66,0,131,0,150,0,217,0,137,0,124,0,227,0,23,0,0,0,191,0,147,0,0,0,0,0,154,0,181,0,0,0,189,0,0,0,168,0,87,0,38,0,101,0,0,0,156,0,185,0,0,0,88,0,0,0,160,0,22,0,241,0,218,0,184,0,117,0,19,0,3,0,31,0,0,0,201,0,61,0,48,0,114,0,0,0,230,0,14,0,142,0,106,0,246,0,148,0,112,0,13,0,22,0,156,0,0,0,123,0,114,0,191,0,126,0,20,0,206,0,41,0,216,0,19,0,96,0,242,0,195,0,52,0,0,0,237,0,0,0,0,0,189,0,222,0,97,0,189,0,60,0,200,0,213,0,230,0,173,0,62,0,193,0,39,0,56,0,216,0,52,0,48,0,41,0,43,0,0,0,219,0,151,0,98,0,45,0,120,0,183,0,0,0,0,0,79,0,131,0,243,0,28,0,32,0,209,0,92,0,107,0,10,0,0,0,61,0,0,0,40,0,0,0,204,0,155,0,253,0,111,0,247,0,27,0,0,0,210,0,0,0,133,0,120,0,0,0,0,0,235,0,0,0,78,0,0,0,116,0,249,0,180,0,209,0,42,0,180,0,160,0,189,0,74,0,0,0,222,0,159,0,248,0,0,0,40,0,252,0,244,0,0,0,223,0,174,0,0,0,19,0,253,0,232,0,6,0,68,0,235,0,209,0,45,0,166,0,0,0,235,0,251,0,247,0,187,0,121,0,206,0,0,0,121,0,37,0,0,0,158,0,219,0,213,0,141,0,17,0,166,0,212,0,194,0,143,0,214,0,0,0,172,0,242,0,0,0,255,0,159,0,252,0,58,0,126,0,247,0,191,0,139,0,83,0,0,0,172,0,0,0,0,0,16,0,193,0,155,0,115,0,0,0,5,0,35,0,175,0,99,0,111,0,242,0,82,0,87,0,199,0,0,0,103,0,183,0,0,0,119,0,244,0,131,0,0,0,104,0,192,0,0,0,24,0,38,0,0,0,0,0,62,0,192,0,127,0,183,0,140,0,153,0,129,0,238,0,236,0,43,0,93,0,45,0,163,0,46,0,0,0,188,0,236,0,26,0,72,0,100,0,0,0,201,0,226,0,28,0,25,0,43,0,0,0,197,0,175,0,145,0,48,0,208,0,213,0,224,0,0,0,0,0,0,0,106,0,81,0,112,0);
signal scenario_full  : scenario_type := (206,31,254,31,247,31,99,31,37,31,104,31,6,31,199,31,181,31,103,31,102,31,216,31,23,31,255,31,190,31,182,31,182,30,169,31,102,31,233,31,233,30,66,31,66,30,122,31,206,31,182,31,19,31,235,31,221,31,101,31,121,31,215,31,231,31,231,30,10,31,126,31,247,31,188,31,112,31,180,31,180,30,154,31,154,31,121,31,38,31,167,31,248,31,248,30,248,29,49,31,139,31,232,31,241,31,34,31,218,31,37,31,142,31,216,31,216,30,216,31,216,30,240,31,153,31,124,31,213,31,134,31,204,31,204,30,204,29,97,31,218,31,189,31,232,31,198,31,14,31,134,31,106,31,147,31,189,31,4,31,252,31,221,31,57,31,217,31,188,31,180,31,248,31,222,31,16,31,70,31,47,31,140,31,170,31,170,30,129,31,142,31,142,30,142,29,10,31,172,31,226,31,236,31,11,31,39,31,160,31,160,30,19,31,191,31,119,31,66,31,35,31,1,31,42,31,171,31,55,31,55,30,69,31,110,31,199,31,33,31,115,31,184,31,66,31,131,31,150,31,217,31,137,31,124,31,227,31,23,31,23,30,191,31,147,31,147,30,147,29,154,31,181,31,181,30,189,31,189,30,168,31,87,31,38,31,101,31,101,30,156,31,185,31,185,30,88,31,88,30,160,31,22,31,241,31,218,31,184,31,117,31,19,31,3,31,31,31,31,30,201,31,61,31,48,31,114,31,114,30,230,31,14,31,142,31,106,31,246,31,148,31,112,31,13,31,22,31,156,31,156,30,123,31,114,31,191,31,126,31,20,31,206,31,41,31,216,31,19,31,96,31,242,31,195,31,52,31,52,30,237,31,237,30,237,29,189,31,222,31,97,31,189,31,60,31,200,31,213,31,230,31,173,31,62,31,193,31,39,31,56,31,216,31,52,31,48,31,41,31,43,31,43,30,219,31,151,31,98,31,45,31,120,31,183,31,183,30,183,29,79,31,131,31,243,31,28,31,32,31,209,31,92,31,107,31,10,31,10,30,61,31,61,30,40,31,40,30,204,31,155,31,253,31,111,31,247,31,27,31,27,30,210,31,210,30,133,31,120,31,120,30,120,29,235,31,235,30,78,31,78,30,116,31,249,31,180,31,209,31,42,31,180,31,160,31,189,31,74,31,74,30,222,31,159,31,248,31,248,30,40,31,252,31,244,31,244,30,223,31,174,31,174,30,19,31,253,31,232,31,6,31,68,31,235,31,209,31,45,31,166,31,166,30,235,31,251,31,247,31,187,31,121,31,206,31,206,30,121,31,37,31,37,30,158,31,219,31,213,31,141,31,17,31,166,31,212,31,194,31,143,31,214,31,214,30,172,31,242,31,242,30,255,31,159,31,252,31,58,31,126,31,247,31,191,31,139,31,83,31,83,30,172,31,172,30,172,29,16,31,193,31,155,31,115,31,115,30,5,31,35,31,175,31,99,31,111,31,242,31,82,31,87,31,199,31,199,30,103,31,183,31,183,30,119,31,244,31,131,31,131,30,104,31,192,31,192,30,24,31,38,31,38,30,38,29,62,31,192,31,127,31,183,31,140,31,153,31,129,31,238,31,236,31,43,31,93,31,45,31,163,31,46,31,46,30,188,31,236,31,26,31,72,31,100,31,100,30,201,31,226,31,28,31,25,31,43,31,43,30,197,31,175,31,145,31,48,31,208,31,213,31,224,31,224,30,224,29,224,28,106,31,81,31,112,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
