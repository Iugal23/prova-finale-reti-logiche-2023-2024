-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_687 is
end project_tb_687;

architecture project_tb_arch_687 of project_tb_687 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 650;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (189,0,193,0,176,0,0,0,239,0,209,0,0,0,0,0,0,0,25,0,24,0,230,0,254,0,0,0,148,0,174,0,0,0,6,0,0,0,230,0,202,0,222,0,0,0,159,0,0,0,0,0,146,0,30,0,238,0,27,0,172,0,140,0,174,0,0,0,247,0,203,0,193,0,0,0,52,0,32,0,54,0,162,0,45,0,48,0,155,0,0,0,0,0,86,0,155,0,17,0,208,0,155,0,168,0,227,0,0,0,94,0,33,0,146,0,178,0,242,0,122,0,200,0,122,0,120,0,16,0,0,0,78,0,239,0,175,0,58,0,214,0,54,0,85,0,12,0,94,0,136,0,222,0,198,0,4,0,214,0,0,0,226,0,241,0,234,0,0,0,0,0,165,0,238,0,0,0,0,0,8,0,196,0,123,0,177,0,12,0,96,0,106,0,140,0,38,0,0,0,55,0,2,0,134,0,59,0,206,0,67,0,169,0,211,0,0,0,170,0,110,0,110,0,92,0,0,0,246,0,97,0,87,0,177,0,62,0,178,0,6,0,73,0,108,0,58,0,98,0,209,0,10,0,89,0,37,0,0,0,0,0,90,0,46,0,0,0,143,0,125,0,0,0,0,0,84,0,233,0,93,0,98,0,132,0,178,0,168,0,233,0,0,0,30,0,14,0,44,0,238,0,0,0,149,0,230,0,228,0,128,0,167,0,137,0,218,0,50,0,222,0,89,0,219,0,0,0,7,0,31,0,0,0,7,0,124,0,227,0,79,0,182,0,154,0,104,0,208,0,74,0,68,0,118,0,45,0,216,0,167,0,9,0,23,0,158,0,229,0,88,0,138,0,110,0,118,0,0,0,206,0,54,0,124,0,154,0,232,0,0,0,103,0,215,0,140,0,125,0,30,0,223,0,17,0,61,0,0,0,152,0,0,0,225,0,88,0,53,0,54,0,0,0,135,0,92,0,0,0,0,0,211,0,111,0,110,0,205,0,143,0,30,0,122,0,19,0,73,0,217,0,0,0,51,0,171,0,218,0,159,0,192,0,0,0,211,0,0,0,63,0,0,0,13,0,70,0,135,0,179,0,232,0,253,0,6,0,188,0,198,0,249,0,105,0,25,0,27,0,164,0,98,0,7,0,205,0,60,0,23,0,5,0,63,0,0,0,206,0,221,0,65,0,30,0,244,0,85,0,229,0,73,0,203,0,32,0,138,0,182,0,106,0,168,0,74,0,162,0,11,0,91,0,181,0,0,0,154,0,0,0,2,0,139,0,42,0,130,0,0,0,147,0,0,0,0,0,105,0,25,0,78,0,100,0,15,0,0,0,156,0,74,0,0,0,242,0,106,0,172,0,121,0,126,0,165,0,61,0,131,0,173,0,171,0,0,0,0,0,236,0,88,0,167,0,188,0,211,0,40,0,0,0,252,0,123,0,0,0,0,0,145,0,65,0,0,0,249,0,0,0,0,0,128,0,143,0,221,0,0,0,156,0,60,0,130,0,0,0,14,0,181,0,207,0,142,0,84,0,14,0,61,0,127,0,89,0,179,0,219,0,99,0,187,0,162,0,0,0,144,0,82,0,179,0,164,0,245,0,210,0,0,0,233,0,109,0,0,0,33,0,19,0,240,0,122,0,0,0,208,0,49,0,97,0,0,0,0,0,194,0,50,0,195,0,214,0,134,0,239,0,57,0,234,0,241,0,0,0,23,0,11,0,72,0,0,0,0,0,249,0,106,0,54,0,236,0,176,0,37,0,0,0,148,0,0,0,69,0,255,0,44,0,174,0,110,0,11,0,253,0,86,0,0,0,0,0,0,0,53,0,228,0,160,0,80,0,99,0,0,0,110,0,150,0,86,0,0,0,139,0,28,0,0,0,209,0,48,0,95,0,242,0,204,0,5,0,127,0,124,0,64,0,209,0,231,0,17,0,250,0,234,0,28,0,154,0,163,0,172,0,150,0,214,0,228,0,159,0,117,0,5,0,61,0,182,0,246,0,243,0,166,0,0,0,0,0,255,0,25,0,0,0,0,0,196,0,27,0,68,0,73,0,113,0,0,0,19,0,189,0,0,0,20,0,239,0,0,0,143,0,0,0,248,0,167,0,0,0,10,0,0,0,33,0,197,0,0,0,75,0,208,0,61,0,70,0,0,0,0,0,0,0,224,0,126,0,104,0,59,0,151,0,0,0,0,0,0,0,74,0,42,0,116,0,17,0,0,0,209,0,155,0,123,0,190,0,25,0,154,0,0,0,195,0,100,0,56,0,0,0,176,0,82,0,226,0,162,0,150,0,252,0,77,0,167,0,15,0,242,0,6,0,98,0,26,0,48,0,0,0,64,0,0,0,244,0,206,0,117,0,0,0,237,0,0,0,7,0,1,0,20,0,95,0,145,0,158,0,0,0,200,0,52,0,251,0,115,0,36,0,177,0,43,0,43,0,234,0,218,0,243,0,92,0,113,0,120,0,0,0,223,0,188,0,0,0,100,0,221,0,162,0,52,0,90,0,248,0,226,0,217,0,187,0,157,0,167,0,0,0,242,0,22,0,0,0,197,0,42,0,166,0,70,0,102,0,0,0,6,0,0,0,29,0,0,0,36,0,110,0,216,0,246,0,144,0,74,0,236,0,138,0,0,0,104,0,122,0,0,0,37,0,0,0,8,0,231,0,246,0,217,0,0,0,0,0,0,0,84,0,204,0,98,0,179,0,223,0,67,0,117,0,245,0,248,0,0,0,47,0,188,0,0,0,36,0,0,0,62,0,0,0,60,0,0,0,29,0,89,0,228,0,147,0,0,0,36,0,159,0,200,0,105,0,217,0,110,0,60,0,158,0,0,0,232,0,162,0,68,0,92,0,83,0,175,0,0,0,123,0,156,0,25,0,28,0,124,0,219,0,112,0,215,0,0,0,35,0);
signal scenario_full  : scenario_type := (189,31,193,31,176,31,176,30,239,31,209,31,209,30,209,29,209,28,25,31,24,31,230,31,254,31,254,30,148,31,174,31,174,30,6,31,6,30,230,31,202,31,222,31,222,30,159,31,159,30,159,29,146,31,30,31,238,31,27,31,172,31,140,31,174,31,174,30,247,31,203,31,193,31,193,30,52,31,32,31,54,31,162,31,45,31,48,31,155,31,155,30,155,29,86,31,155,31,17,31,208,31,155,31,168,31,227,31,227,30,94,31,33,31,146,31,178,31,242,31,122,31,200,31,122,31,120,31,16,31,16,30,78,31,239,31,175,31,58,31,214,31,54,31,85,31,12,31,94,31,136,31,222,31,198,31,4,31,214,31,214,30,226,31,241,31,234,31,234,30,234,29,165,31,238,31,238,30,238,29,8,31,196,31,123,31,177,31,12,31,96,31,106,31,140,31,38,31,38,30,55,31,2,31,134,31,59,31,206,31,67,31,169,31,211,31,211,30,170,31,110,31,110,31,92,31,92,30,246,31,97,31,87,31,177,31,62,31,178,31,6,31,73,31,108,31,58,31,98,31,209,31,10,31,89,31,37,31,37,30,37,29,90,31,46,31,46,30,143,31,125,31,125,30,125,29,84,31,233,31,93,31,98,31,132,31,178,31,168,31,233,31,233,30,30,31,14,31,44,31,238,31,238,30,149,31,230,31,228,31,128,31,167,31,137,31,218,31,50,31,222,31,89,31,219,31,219,30,7,31,31,31,31,30,7,31,124,31,227,31,79,31,182,31,154,31,104,31,208,31,74,31,68,31,118,31,45,31,216,31,167,31,9,31,23,31,158,31,229,31,88,31,138,31,110,31,118,31,118,30,206,31,54,31,124,31,154,31,232,31,232,30,103,31,215,31,140,31,125,31,30,31,223,31,17,31,61,31,61,30,152,31,152,30,225,31,88,31,53,31,54,31,54,30,135,31,92,31,92,30,92,29,211,31,111,31,110,31,205,31,143,31,30,31,122,31,19,31,73,31,217,31,217,30,51,31,171,31,218,31,159,31,192,31,192,30,211,31,211,30,63,31,63,30,13,31,70,31,135,31,179,31,232,31,253,31,6,31,188,31,198,31,249,31,105,31,25,31,27,31,164,31,98,31,7,31,205,31,60,31,23,31,5,31,63,31,63,30,206,31,221,31,65,31,30,31,244,31,85,31,229,31,73,31,203,31,32,31,138,31,182,31,106,31,168,31,74,31,162,31,11,31,91,31,181,31,181,30,154,31,154,30,2,31,139,31,42,31,130,31,130,30,147,31,147,30,147,29,105,31,25,31,78,31,100,31,15,31,15,30,156,31,74,31,74,30,242,31,106,31,172,31,121,31,126,31,165,31,61,31,131,31,173,31,171,31,171,30,171,29,236,31,88,31,167,31,188,31,211,31,40,31,40,30,252,31,123,31,123,30,123,29,145,31,65,31,65,30,249,31,249,30,249,29,128,31,143,31,221,31,221,30,156,31,60,31,130,31,130,30,14,31,181,31,207,31,142,31,84,31,14,31,61,31,127,31,89,31,179,31,219,31,99,31,187,31,162,31,162,30,144,31,82,31,179,31,164,31,245,31,210,31,210,30,233,31,109,31,109,30,33,31,19,31,240,31,122,31,122,30,208,31,49,31,97,31,97,30,97,29,194,31,50,31,195,31,214,31,134,31,239,31,57,31,234,31,241,31,241,30,23,31,11,31,72,31,72,30,72,29,249,31,106,31,54,31,236,31,176,31,37,31,37,30,148,31,148,30,69,31,255,31,44,31,174,31,110,31,11,31,253,31,86,31,86,30,86,29,86,28,53,31,228,31,160,31,80,31,99,31,99,30,110,31,150,31,86,31,86,30,139,31,28,31,28,30,209,31,48,31,95,31,242,31,204,31,5,31,127,31,124,31,64,31,209,31,231,31,17,31,250,31,234,31,28,31,154,31,163,31,172,31,150,31,214,31,228,31,159,31,117,31,5,31,61,31,182,31,246,31,243,31,166,31,166,30,166,29,255,31,25,31,25,30,25,29,196,31,27,31,68,31,73,31,113,31,113,30,19,31,189,31,189,30,20,31,239,31,239,30,143,31,143,30,248,31,167,31,167,30,10,31,10,30,33,31,197,31,197,30,75,31,208,31,61,31,70,31,70,30,70,29,70,28,224,31,126,31,104,31,59,31,151,31,151,30,151,29,151,28,74,31,42,31,116,31,17,31,17,30,209,31,155,31,123,31,190,31,25,31,154,31,154,30,195,31,100,31,56,31,56,30,176,31,82,31,226,31,162,31,150,31,252,31,77,31,167,31,15,31,242,31,6,31,98,31,26,31,48,31,48,30,64,31,64,30,244,31,206,31,117,31,117,30,237,31,237,30,7,31,1,31,20,31,95,31,145,31,158,31,158,30,200,31,52,31,251,31,115,31,36,31,177,31,43,31,43,31,234,31,218,31,243,31,92,31,113,31,120,31,120,30,223,31,188,31,188,30,100,31,221,31,162,31,52,31,90,31,248,31,226,31,217,31,187,31,157,31,167,31,167,30,242,31,22,31,22,30,197,31,42,31,166,31,70,31,102,31,102,30,6,31,6,30,29,31,29,30,36,31,110,31,216,31,246,31,144,31,74,31,236,31,138,31,138,30,104,31,122,31,122,30,37,31,37,30,8,31,231,31,246,31,217,31,217,30,217,29,217,28,84,31,204,31,98,31,179,31,223,31,67,31,117,31,245,31,248,31,248,30,47,31,188,31,188,30,36,31,36,30,62,31,62,30,60,31,60,30,29,31,89,31,228,31,147,31,147,30,36,31,159,31,200,31,105,31,217,31,110,31,60,31,158,31,158,30,232,31,162,31,68,31,92,31,83,31,175,31,175,30,123,31,156,31,25,31,28,31,124,31,219,31,112,31,215,31,215,30,35,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
