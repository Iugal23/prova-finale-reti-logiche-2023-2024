-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_250 is
end project_tb_250;

architecture project_tb_arch_250 of project_tb_250 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 467;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (179,0,62,0,133,0,246,0,48,0,191,0,9,0,178,0,0,0,80,0,0,0,180,0,0,0,252,0,30,0,0,0,14,0,0,0,67,0,35,0,65,0,0,0,181,0,36,0,44,0,112,0,230,0,61,0,113,0,0,0,0,0,99,0,118,0,0,0,0,0,171,0,198,0,70,0,0,0,0,0,0,0,251,0,68,0,207,0,204,0,176,0,220,0,53,0,0,0,250,0,34,0,0,0,0,0,211,0,209,0,127,0,115,0,0,0,140,0,157,0,90,0,7,0,234,0,30,0,23,0,28,0,41,0,0,0,34,0,39,0,44,0,28,0,101,0,0,0,69,0,213,0,0,0,0,0,244,0,207,0,189,0,186,0,190,0,82,0,73,0,0,0,239,0,99,0,222,0,0,0,229,0,205,0,0,0,225,0,220,0,98,0,0,0,161,0,44,0,153,0,191,0,210,0,20,0,67,0,215,0,96,0,19,0,248,0,14,0,214,0,167,0,59,0,117,0,195,0,93,0,101,0,124,0,241,0,128,0,37,0,123,0,208,0,220,0,0,0,0,0,3,0,0,0,173,0,69,0,129,0,177,0,0,0,0,0,16,0,247,0,118,0,0,0,133,0,0,0,123,0,42,0,171,0,49,0,1,0,136,0,0,0,169,0,0,0,186,0,227,0,0,0,229,0,0,0,173,0,88,0,214,0,130,0,54,0,87,0,6,0,71,0,204,0,165,0,63,0,220,0,43,0,0,0,167,0,254,0,85,0,194,0,12,0,17,0,27,0,0,0,201,0,0,0,249,0,85,0,214,0,38,0,0,0,164,0,0,0,0,0,0,0,0,0,143,0,0,0,93,0,0,0,212,0,206,0,127,0,22,0,184,0,70,0,68,0,86,0,235,0,21,0,0,0,59,0,198,0,63,0,189,0,196,0,130,0,112,0,170,0,152,0,0,0,234,0,238,0,239,0,174,0,87,0,51,0,0,0,45,0,0,0,48,0,0,0,205,0,40,0,0,0,180,0,33,0,90,0,33,0,191,0,206,0,29,0,0,0,214,0,103,0,95,0,2,0,0,0,100,0,117,0,169,0,100,0,0,0,0,0,0,0,72,0,0,0,0,0,116,0,0,0,0,0,75,0,78,0,74,0,49,0,22,0,27,0,201,0,228,0,33,0,113,0,121,0,9,0,39,0,193,0,92,0,71,0,0,0,0,0,103,0,249,0,114,0,200,0,0,0,0,0,204,0,14,0,98,0,16,0,83,0,0,0,145,0,0,0,163,0,203,0,119,0,126,0,66,0,0,0,0,0,184,0,89,0,72,0,23,0,45,0,231,0,0,0,165,0,122,0,187,0,3,0,146,0,0,0,242,0,151,0,238,0,0,0,0,0,12,0,0,0,59,0,0,0,50,0,131,0,60,0,219,0,226,0,67,0,195,0,121,0,252,0,50,0,102,0,233,0,188,0,0,0,0,0,86,0,16,0,8,0,0,0,0,0,120,0,0,0,107,0,154,0,127,0,228,0,170,0,55,0,80,0,137,0,5,0,216,0,186,0,235,0,112,0,51,0,185,0,84,0,35,0,0,0,82,0,242,0,0,0,44,0,180,0,84,0,129,0,3,0,123,0,0,0,0,0,6,0,0,0,14,0,41,0,202,0,174,0,12,0,18,0,203,0,65,0,39,0,98,0,172,0,113,0,183,0,0,0,0,0,111,0,110,0,196,0,0,0,220,0,166,0,0,0,40,0,44,0,142,0,54,0,22,0,205,0,41,0,0,0,85,0,230,0,0,0,91,0,56,0,0,0,0,0,0,0,242,0,146,0,181,0,155,0,212,0,158,0,191,0,5,0,0,0,35,0,246,0,47,0,49,0,193,0,222,0,111,0,133,0,6,0,31,0,229,0,88,0,225,0,0,0,68,0,0,0,44,0,0,0,92,0,4,0,47,0,159,0,12,0,167,0,81,0,125,0,41,0,93,0,30,0,106,0,0,0,7,0,213,0,105,0,0,0,11,0,219,0,5,0,229,0,13,0,83,0,0,0,67,0,169,0,25,0,0,0,137,0,230,0,0,0,51,0,177,0,236,0,0,0,0,0);
signal scenario_full  : scenario_type := (179,31,62,31,133,31,246,31,48,31,191,31,9,31,178,31,178,30,80,31,80,30,180,31,180,30,252,31,30,31,30,30,14,31,14,30,67,31,35,31,65,31,65,30,181,31,36,31,44,31,112,31,230,31,61,31,113,31,113,30,113,29,99,31,118,31,118,30,118,29,171,31,198,31,70,31,70,30,70,29,70,28,251,31,68,31,207,31,204,31,176,31,220,31,53,31,53,30,250,31,34,31,34,30,34,29,211,31,209,31,127,31,115,31,115,30,140,31,157,31,90,31,7,31,234,31,30,31,23,31,28,31,41,31,41,30,34,31,39,31,44,31,28,31,101,31,101,30,69,31,213,31,213,30,213,29,244,31,207,31,189,31,186,31,190,31,82,31,73,31,73,30,239,31,99,31,222,31,222,30,229,31,205,31,205,30,225,31,220,31,98,31,98,30,161,31,44,31,153,31,191,31,210,31,20,31,67,31,215,31,96,31,19,31,248,31,14,31,214,31,167,31,59,31,117,31,195,31,93,31,101,31,124,31,241,31,128,31,37,31,123,31,208,31,220,31,220,30,220,29,3,31,3,30,173,31,69,31,129,31,177,31,177,30,177,29,16,31,247,31,118,31,118,30,133,31,133,30,123,31,42,31,171,31,49,31,1,31,136,31,136,30,169,31,169,30,186,31,227,31,227,30,229,31,229,30,173,31,88,31,214,31,130,31,54,31,87,31,6,31,71,31,204,31,165,31,63,31,220,31,43,31,43,30,167,31,254,31,85,31,194,31,12,31,17,31,27,31,27,30,201,31,201,30,249,31,85,31,214,31,38,31,38,30,164,31,164,30,164,29,164,28,164,27,143,31,143,30,93,31,93,30,212,31,206,31,127,31,22,31,184,31,70,31,68,31,86,31,235,31,21,31,21,30,59,31,198,31,63,31,189,31,196,31,130,31,112,31,170,31,152,31,152,30,234,31,238,31,239,31,174,31,87,31,51,31,51,30,45,31,45,30,48,31,48,30,205,31,40,31,40,30,180,31,33,31,90,31,33,31,191,31,206,31,29,31,29,30,214,31,103,31,95,31,2,31,2,30,100,31,117,31,169,31,100,31,100,30,100,29,100,28,72,31,72,30,72,29,116,31,116,30,116,29,75,31,78,31,74,31,49,31,22,31,27,31,201,31,228,31,33,31,113,31,121,31,9,31,39,31,193,31,92,31,71,31,71,30,71,29,103,31,249,31,114,31,200,31,200,30,200,29,204,31,14,31,98,31,16,31,83,31,83,30,145,31,145,30,163,31,203,31,119,31,126,31,66,31,66,30,66,29,184,31,89,31,72,31,23,31,45,31,231,31,231,30,165,31,122,31,187,31,3,31,146,31,146,30,242,31,151,31,238,31,238,30,238,29,12,31,12,30,59,31,59,30,50,31,131,31,60,31,219,31,226,31,67,31,195,31,121,31,252,31,50,31,102,31,233,31,188,31,188,30,188,29,86,31,16,31,8,31,8,30,8,29,120,31,120,30,107,31,154,31,127,31,228,31,170,31,55,31,80,31,137,31,5,31,216,31,186,31,235,31,112,31,51,31,185,31,84,31,35,31,35,30,82,31,242,31,242,30,44,31,180,31,84,31,129,31,3,31,123,31,123,30,123,29,6,31,6,30,14,31,41,31,202,31,174,31,12,31,18,31,203,31,65,31,39,31,98,31,172,31,113,31,183,31,183,30,183,29,111,31,110,31,196,31,196,30,220,31,166,31,166,30,40,31,44,31,142,31,54,31,22,31,205,31,41,31,41,30,85,31,230,31,230,30,91,31,56,31,56,30,56,29,56,28,242,31,146,31,181,31,155,31,212,31,158,31,191,31,5,31,5,30,35,31,246,31,47,31,49,31,193,31,222,31,111,31,133,31,6,31,31,31,229,31,88,31,225,31,225,30,68,31,68,30,44,31,44,30,92,31,4,31,47,31,159,31,12,31,167,31,81,31,125,31,41,31,93,31,30,31,106,31,106,30,7,31,213,31,105,31,105,30,11,31,219,31,5,31,229,31,13,31,83,31,83,30,67,31,169,31,25,31,25,30,137,31,230,31,230,30,51,31,177,31,236,31,236,30,236,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
