-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 682;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (68,0,84,0,41,0,233,0,23,0,0,0,128,0,189,0,151,0,26,0,0,0,0,0,72,0,111,0,10,0,122,0,130,0,140,0,85,0,19,0,172,0,237,0,47,0,0,0,121,0,138,0,225,0,192,0,172,0,89,0,176,0,0,0,0,0,0,0,130,0,118,0,104,0,139,0,146,0,33,0,8,0,177,0,253,0,31,0,242,0,237,0,247,0,0,0,52,0,143,0,60,0,241,0,188,0,108,0,0,0,96,0,181,0,0,0,244,0,65,0,165,0,212,0,247,0,135,0,3,0,143,0,110,0,175,0,54,0,140,0,0,0,74,0,0,0,0,0,67,0,98,0,109,0,215,0,199,0,0,0,0,0,0,0,162,0,25,0,0,0,112,0,0,0,225,0,192,0,87,0,253,0,0,0,0,0,153,0,83,0,166,0,251,0,113,0,44,0,85,0,76,0,24,0,55,0,54,0,76,0,32,0,0,0,135,0,87,0,0,0,249,0,62,0,168,0,214,0,88,0,53,0,0,0,37,0,127,0,10,0,14,0,198,0,38,0,83,0,189,0,0,0,41,0,197,0,27,0,194,0,0,0,7,0,31,0,0,0,0,0,27,0,243,0,173,0,202,0,87,0,31,0,0,0,125,0,51,0,212,0,229,0,92,0,126,0,190,0,71,0,29,0,230,0,124,0,152,0,154,0,0,0,250,0,231,0,59,0,34,0,128,0,64,0,20,0,152,0,105,0,105,0,54,0,22,0,0,0,252,0,163,0,9,0,40,0,3,0,0,0,139,0,0,0,167,0,176,0,162,0,87,0,0,0,0,0,77,0,0,0,0,0,96,0,73,0,36,0,104,0,104,0,176,0,119,0,87,0,28,0,198,0,60,0,167,0,0,0,56,0,26,0,66,0,28,0,124,0,193,0,12,0,0,0,249,0,223,0,142,0,0,0,75,0,10,0,235,0,37,0,0,0,144,0,200,0,0,0,0,0,17,0,0,0,36,0,82,0,33,0,194,0,0,0,118,0,83,0,198,0,37,0,96,0,228,0,0,0,143,0,0,0,0,0,133,0,0,0,246,0,183,0,109,0,0,0,0,0,22,0,78,0,167,0,252,0,152,0,0,0,104,0,77,0,255,0,6,0,148,0,194,0,56,0,0,0,0,0,12,0,208,0,203,0,0,0,174,0,0,0,166,0,127,0,157,0,215,0,151,0,82,0,132,0,0,0,46,0,15,0,0,0,40,0,249,0,78,0,248,0,22,0,0,0,241,0,118,0,170,0,52,0,244,0,143,0,30,0,95,0,0,0,221,0,0,0,117,0,7,0,4,0,95,0,195,0,180,0,63,0,210,0,0,0,178,0,207,0,236,0,150,0,0,0,0,0,0,0,0,0,201,0,0,0,179,0,201,0,25,0,6,0,123,0,0,0,202,0,124,0,80,0,61,0,174,0,137,0,48,0,65,0,148,0,105,0,0,0,11,0,58,0,176,0,255,0,38,0,99,0,20,0,148,0,146,0,28,0,110,0,66,0,163,0,205,0,205,0,120,0,211,0,101,0,132,0,175,0,52,0,199,0,228,0,219,0,38,0,65,0,207,0,6,0,50,0,0,0,105,0,236,0,0,0,0,0,191,0,187,0,18,0,17,0,117,0,17,0,81,0,74,0,103,0,2,0,59,0,120,0,0,0,0,0,5,0,139,0,0,0,95,0,153,0,215,0,218,0,169,0,155,0,108,0,228,0,236,0,0,0,236,0,181,0,213,0,58,0,207,0,195,0,225,0,117,0,0,0,218,0,36,0,101,0,164,0,246,0,238,0,132,0,233,0,0,0,0,0,5,0,207,0,227,0,0,0,170,0,131,0,0,0,0,0,124,0,152,0,239,0,46,0,152,0,38,0,244,0,41,0,120,0,237,0,149,0,13,0,192,0,196,0,67,0,80,0,234,0,216,0,2,0,9,0,32,0,0,0,62,0,25,0,14,0,0,0,226,0,12,0,168,0,131,0,211,0,157,0,4,0,109,0,92,0,193,0,227,0,226,0,211,0,63,0,27,0,221,0,160,0,216,0,108,0,239,0,47,0,220,0,0,0,170,0,0,0,228,0,49,0,0,0,93,0,131,0,157,0,30,0,28,0,0,0,96,0,167,0,10,0,54,0,57,0,116,0,0,0,0,0,181,0,38,0,73,0,241,0,248,0,38,0,0,0,132,0,80,0,26,0,218,0,0,0,0,0,134,0,72,0,31,0,163,0,209,0,170,0,0,0,0,0,70,0,172,0,188,0,66,0,105,0,53,0,34,0,0,0,16,0,10,0,241,0,116,0,192,0,0,0,0,0,231,0,184,0,156,0,184,0,0,0,193,0,147,0,144,0,0,0,213,0,82,0,78,0,220,0,93,0,0,0,97,0,0,0,0,0,61,0,12,0,173,0,21,0,190,0,0,0,229,0,2,0,0,0,126,0,235,0,49,0,117,0,93,0,0,0,27,0,0,0,55,0,36,0,0,0,90,0,220,0,0,0,0,0,104,0,197,0,9,0,107,0,232,0,46,0,146,0,0,0,9,0,145,0,114,0,45,0,149,0,132,0,251,0,0,0,165,0,196,0,28,0,233,0,0,0,0,0,0,0,237,0,0,0,86,0,143,0,0,0,79,0,202,0,241,0,20,0,244,0,102,0,0,0,255,0,0,0,0,0,170,0,141,0,197,0,9,0,1,0,227,0,0,0,0,0,83,0,142,0,122,0,171,0,118,0,23,0,14,0,105,0,209,0,220,0,4,0,74,0,116,0,0,0,0,0,162,0,146,0,126,0,130,0,177,0,219,0,24,0,122,0,18,0,0,0,151,0,0,0,78,0,188,0,209,0,130,0,131,0,106,0,0,0,51,0,25,0,149,0,135,0,146,0,186,0,49,0,26,0,191,0,141,0,241,0,254,0,72,0,49,0,212,0,11,0,157,0,173,0,33,0,104,0,173,0,0,0,153,0,119,0,64,0,53,0,0,0,0,0,16,0,35,0,219,0,0,0,27,0,225,0,246,0,0,0,54,0,61,0,0,0);
signal scenario_full  : scenario_type := (68,31,84,31,41,31,233,31,23,31,23,30,128,31,189,31,151,31,26,31,26,30,26,29,72,31,111,31,10,31,122,31,130,31,140,31,85,31,19,31,172,31,237,31,47,31,47,30,121,31,138,31,225,31,192,31,172,31,89,31,176,31,176,30,176,29,176,28,130,31,118,31,104,31,139,31,146,31,33,31,8,31,177,31,253,31,31,31,242,31,237,31,247,31,247,30,52,31,143,31,60,31,241,31,188,31,108,31,108,30,96,31,181,31,181,30,244,31,65,31,165,31,212,31,247,31,135,31,3,31,143,31,110,31,175,31,54,31,140,31,140,30,74,31,74,30,74,29,67,31,98,31,109,31,215,31,199,31,199,30,199,29,199,28,162,31,25,31,25,30,112,31,112,30,225,31,192,31,87,31,253,31,253,30,253,29,153,31,83,31,166,31,251,31,113,31,44,31,85,31,76,31,24,31,55,31,54,31,76,31,32,31,32,30,135,31,87,31,87,30,249,31,62,31,168,31,214,31,88,31,53,31,53,30,37,31,127,31,10,31,14,31,198,31,38,31,83,31,189,31,189,30,41,31,197,31,27,31,194,31,194,30,7,31,31,31,31,30,31,29,27,31,243,31,173,31,202,31,87,31,31,31,31,30,125,31,51,31,212,31,229,31,92,31,126,31,190,31,71,31,29,31,230,31,124,31,152,31,154,31,154,30,250,31,231,31,59,31,34,31,128,31,64,31,20,31,152,31,105,31,105,31,54,31,22,31,22,30,252,31,163,31,9,31,40,31,3,31,3,30,139,31,139,30,167,31,176,31,162,31,87,31,87,30,87,29,77,31,77,30,77,29,96,31,73,31,36,31,104,31,104,31,176,31,119,31,87,31,28,31,198,31,60,31,167,31,167,30,56,31,26,31,66,31,28,31,124,31,193,31,12,31,12,30,249,31,223,31,142,31,142,30,75,31,10,31,235,31,37,31,37,30,144,31,200,31,200,30,200,29,17,31,17,30,36,31,82,31,33,31,194,31,194,30,118,31,83,31,198,31,37,31,96,31,228,31,228,30,143,31,143,30,143,29,133,31,133,30,246,31,183,31,109,31,109,30,109,29,22,31,78,31,167,31,252,31,152,31,152,30,104,31,77,31,255,31,6,31,148,31,194,31,56,31,56,30,56,29,12,31,208,31,203,31,203,30,174,31,174,30,166,31,127,31,157,31,215,31,151,31,82,31,132,31,132,30,46,31,15,31,15,30,40,31,249,31,78,31,248,31,22,31,22,30,241,31,118,31,170,31,52,31,244,31,143,31,30,31,95,31,95,30,221,31,221,30,117,31,7,31,4,31,95,31,195,31,180,31,63,31,210,31,210,30,178,31,207,31,236,31,150,31,150,30,150,29,150,28,150,27,201,31,201,30,179,31,201,31,25,31,6,31,123,31,123,30,202,31,124,31,80,31,61,31,174,31,137,31,48,31,65,31,148,31,105,31,105,30,11,31,58,31,176,31,255,31,38,31,99,31,20,31,148,31,146,31,28,31,110,31,66,31,163,31,205,31,205,31,120,31,211,31,101,31,132,31,175,31,52,31,199,31,228,31,219,31,38,31,65,31,207,31,6,31,50,31,50,30,105,31,236,31,236,30,236,29,191,31,187,31,18,31,17,31,117,31,17,31,81,31,74,31,103,31,2,31,59,31,120,31,120,30,120,29,5,31,139,31,139,30,95,31,153,31,215,31,218,31,169,31,155,31,108,31,228,31,236,31,236,30,236,31,181,31,213,31,58,31,207,31,195,31,225,31,117,31,117,30,218,31,36,31,101,31,164,31,246,31,238,31,132,31,233,31,233,30,233,29,5,31,207,31,227,31,227,30,170,31,131,31,131,30,131,29,124,31,152,31,239,31,46,31,152,31,38,31,244,31,41,31,120,31,237,31,149,31,13,31,192,31,196,31,67,31,80,31,234,31,216,31,2,31,9,31,32,31,32,30,62,31,25,31,14,31,14,30,226,31,12,31,168,31,131,31,211,31,157,31,4,31,109,31,92,31,193,31,227,31,226,31,211,31,63,31,27,31,221,31,160,31,216,31,108,31,239,31,47,31,220,31,220,30,170,31,170,30,228,31,49,31,49,30,93,31,131,31,157,31,30,31,28,31,28,30,96,31,167,31,10,31,54,31,57,31,116,31,116,30,116,29,181,31,38,31,73,31,241,31,248,31,38,31,38,30,132,31,80,31,26,31,218,31,218,30,218,29,134,31,72,31,31,31,163,31,209,31,170,31,170,30,170,29,70,31,172,31,188,31,66,31,105,31,53,31,34,31,34,30,16,31,10,31,241,31,116,31,192,31,192,30,192,29,231,31,184,31,156,31,184,31,184,30,193,31,147,31,144,31,144,30,213,31,82,31,78,31,220,31,93,31,93,30,97,31,97,30,97,29,61,31,12,31,173,31,21,31,190,31,190,30,229,31,2,31,2,30,126,31,235,31,49,31,117,31,93,31,93,30,27,31,27,30,55,31,36,31,36,30,90,31,220,31,220,30,220,29,104,31,197,31,9,31,107,31,232,31,46,31,146,31,146,30,9,31,145,31,114,31,45,31,149,31,132,31,251,31,251,30,165,31,196,31,28,31,233,31,233,30,233,29,233,28,237,31,237,30,86,31,143,31,143,30,79,31,202,31,241,31,20,31,244,31,102,31,102,30,255,31,255,30,255,29,170,31,141,31,197,31,9,31,1,31,227,31,227,30,227,29,83,31,142,31,122,31,171,31,118,31,23,31,14,31,105,31,209,31,220,31,4,31,74,31,116,31,116,30,116,29,162,31,146,31,126,31,130,31,177,31,219,31,24,31,122,31,18,31,18,30,151,31,151,30,78,31,188,31,209,31,130,31,131,31,106,31,106,30,51,31,25,31,149,31,135,31,146,31,186,31,49,31,26,31,191,31,141,31,241,31,254,31,72,31,49,31,212,31,11,31,157,31,173,31,33,31,104,31,173,31,173,30,153,31,119,31,64,31,53,31,53,30,53,29,16,31,35,31,219,31,219,30,27,31,225,31,246,31,246,30,54,31,61,31,61,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
