-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 680;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (11,0,174,0,124,0,0,0,177,0,0,0,0,0,123,0,152,0,221,0,98,0,188,0,0,0,5,0,72,0,11,0,138,0,212,0,12,0,48,0,27,0,58,0,198,0,95,0,0,0,198,0,151,0,246,0,221,0,0,0,219,0,71,0,127,0,0,0,127,0,230,0,114,0,152,0,205,0,153,0,139,0,4,0,182,0,254,0,255,0,26,0,114,0,215,0,83,0,137,0,102,0,0,0,37,0,106,0,72,0,66,0,52,0,92,0,132,0,0,0,0,0,153,0,98,0,235,0,167,0,52,0,183,0,118,0,24,0,49,0,246,0,136,0,240,0,84,0,225,0,64,0,27,0,179,0,147,0,38,0,202,0,104,0,156,0,0,0,161,0,0,0,83,0,57,0,126,0,187,0,225,0,199,0,165,0,126,0,0,0,186,0,82,0,0,0,187,0,115,0,144,0,40,0,240,0,250,0,209,0,3,0,3,0,129,0,20,0,0,0,143,0,33,0,242,0,244,0,161,0,120,0,0,0,79,0,6,0,106,0,46,0,214,0,31,0,237,0,0,0,34,0,83,0,164,0,0,0,13,0,67,0,246,0,120,0,17,0,0,0,163,0,181,0,109,0,0,0,78,0,67,0,0,0,187,0,15,0,0,0,39,0,169,0,0,0,8,0,36,0,18,0,118,0,0,0,66,0,202,0,107,0,26,0,109,0,41,0,199,0,8,0,0,0,156,0,252,0,0,0,0,0,95,0,84,0,4,0,111,0,0,0,181,0,203,0,13,0,120,0,182,0,0,0,35,0,4,0,0,0,190,0,160,0,200,0,0,0,227,0,19,0,0,0,4,0,174,0,0,0,53,0,0,0,60,0,150,0,0,0,0,0,10,0,0,0,0,0,0,0,58,0,165,0,62,0,220,0,247,0,0,0,21,0,223,0,0,0,76,0,0,0,105,0,9,0,66,0,0,0,0,0,43,0,49,0,0,0,76,0,0,0,168,0,146,0,111,0,0,0,0,0,0,0,14,0,161,0,50,0,114,0,200,0,235,0,119,0,12,0,7,0,0,0,16,0,150,0,0,0,0,0,0,0,94,0,69,0,164,0,35,0,0,0,244,0,176,0,92,0,182,0,93,0,35,0,133,0,175,0,245,0,0,0,0,0,211,0,0,0,208,0,176,0,237,0,0,0,34,0,47,0,0,0,29,0,240,0,75,0,81,0,0,0,0,0,2,0,192,0,187,0,0,0,34,0,165,0,175,0,239,0,163,0,135,0,244,0,170,0,0,0,130,0,230,0,0,0,207,0,133,0,59,0,56,0,232,0,247,0,45,0,136,0,41,0,255,0,0,0,146,0,109,0,159,0,1,0,240,0,37,0,208,0,84,0,147,0,227,0,0,0,182,0,0,0,182,0,0,0,229,0,36,0,249,0,173,0,54,0,0,0,120,0,147,0,166,0,38,0,101,0,254,0,30,0,20,0,239,0,66,0,19,0,139,0,126,0,20,0,0,0,59,0,240,0,217,0,174,0,226,0,171,0,167,0,200,0,0,0,255,0,63,0,96,0,221,0,44,0,84,0,237,0,0,0,205,0,0,0,0,0,96,0,0,0,179,0,198,0,102,0,198,0,15,0,0,0,0,0,98,0,16,0,251,0,40,0,29,0,0,0,33,0,173,0,33,0,92,0,0,0,24,0,200,0,89,0,37,0,117,0,223,0,180,0,33,0,145,0,71,0,176,0,209,0,4,0,0,0,85,0,153,0,0,0,0,0,54,0,178,0,96,0,2,0,246,0,173,0,21,0,10,0,43,0,248,0,160,0,90,0,158,0,204,0,56,0,15,0,120,0,0,0,74,0,57,0,0,0,121,0,186,0,251,0,92,0,70,0,0,0,20,0,215,0,0,0,0,0,248,0,30,0,153,0,0,0,37,0,0,0,0,0,252,0,128,0,128,0,34,0,26,0,64,0,18,0,184,0,176,0,53,0,22,0,0,0,143,0,16,0,0,0,124,0,113,0,89,0,168,0,25,0,49,0,136,0,168,0,227,0,105,0,200,0,11,0,0,0,11,0,160,0,186,0,248,0,0,0,135,0,238,0,244,0,66,0,163,0,113,0,12,0,250,0,0,0,0,0,7,0,39,0,6,0,43,0,114,0,223,0,179,0,106,0,200,0,138,0,0,0,33,0,9,0,209,0,174,0,176,0,16,0,36,0,121,0,224,0,149,0,213,0,181,0,78,0,197,0,0,0,42,0,7,0,252,0,164,0,115,0,0,0,154,0,177,0,133,0,0,0,204,0,192,0,0,0,221,0,225,0,48,0,0,0,192,0,0,0,137,0,55,0,218,0,254,0,182,0,25,0,229,0,233,0,175,0,99,0,97,0,217,0,36,0,116,0,42,0,53,0,153,0,134,0,0,0,249,0,145,0,0,0,184,0,99,0,120,0,19,0,239,0,47,0,75,0,0,0,140,0,90,0,81,0,121,0,66,0,161,0,158,0,0,0,0,0,173,0,0,0,248,0,244,0,196,0,19,0,0,0,51,0,0,0,0,0,24,0,0,0,248,0,104,0,107,0,63,0,71,0,21,0,0,0,52,0,177,0,67,0,0,0,232,0,146,0,53,0,2,0,191,0,114,0,0,0,0,0,13,0,31,0,233,0,19,0,147,0,174,0,86,0,28,0,242,0,223,0,221,0,166,0,254,0,0,0,59,0,0,0,171,0,175,0,145,0,130,0,65,0,1,0,178,0,239,0,0,0,145,0,153,0,243,0,0,0,158,0,145,0,192,0,5,0,157,0,160,0,0,0,132,0,27,0,113,0,102,0,113,0,11,0,0,0,44,0,0,0,0,0,0,0,82,0,69,0,225,0,136,0,160,0,0,0,63,0,196,0,137,0,48,0,66,0,135,0,22,0,0,0,0,0,51,0,0,0,125,0,209,0,33,0,0,0,65,0,175,0,120,0,164,0,10,0,202,0,0,0,27,0,225,0,190,0,65,0,0,0,91,0,167,0,127,0,4,0,92,0,154,0,41,0,194,0,178,0,209,0);
signal scenario_full  : scenario_type := (11,31,174,31,124,31,124,30,177,31,177,30,177,29,123,31,152,31,221,31,98,31,188,31,188,30,5,31,72,31,11,31,138,31,212,31,12,31,48,31,27,31,58,31,198,31,95,31,95,30,198,31,151,31,246,31,221,31,221,30,219,31,71,31,127,31,127,30,127,31,230,31,114,31,152,31,205,31,153,31,139,31,4,31,182,31,254,31,255,31,26,31,114,31,215,31,83,31,137,31,102,31,102,30,37,31,106,31,72,31,66,31,52,31,92,31,132,31,132,30,132,29,153,31,98,31,235,31,167,31,52,31,183,31,118,31,24,31,49,31,246,31,136,31,240,31,84,31,225,31,64,31,27,31,179,31,147,31,38,31,202,31,104,31,156,31,156,30,161,31,161,30,83,31,57,31,126,31,187,31,225,31,199,31,165,31,126,31,126,30,186,31,82,31,82,30,187,31,115,31,144,31,40,31,240,31,250,31,209,31,3,31,3,31,129,31,20,31,20,30,143,31,33,31,242,31,244,31,161,31,120,31,120,30,79,31,6,31,106,31,46,31,214,31,31,31,237,31,237,30,34,31,83,31,164,31,164,30,13,31,67,31,246,31,120,31,17,31,17,30,163,31,181,31,109,31,109,30,78,31,67,31,67,30,187,31,15,31,15,30,39,31,169,31,169,30,8,31,36,31,18,31,118,31,118,30,66,31,202,31,107,31,26,31,109,31,41,31,199,31,8,31,8,30,156,31,252,31,252,30,252,29,95,31,84,31,4,31,111,31,111,30,181,31,203,31,13,31,120,31,182,31,182,30,35,31,4,31,4,30,190,31,160,31,200,31,200,30,227,31,19,31,19,30,4,31,174,31,174,30,53,31,53,30,60,31,150,31,150,30,150,29,10,31,10,30,10,29,10,28,58,31,165,31,62,31,220,31,247,31,247,30,21,31,223,31,223,30,76,31,76,30,105,31,9,31,66,31,66,30,66,29,43,31,49,31,49,30,76,31,76,30,168,31,146,31,111,31,111,30,111,29,111,28,14,31,161,31,50,31,114,31,200,31,235,31,119,31,12,31,7,31,7,30,16,31,150,31,150,30,150,29,150,28,94,31,69,31,164,31,35,31,35,30,244,31,176,31,92,31,182,31,93,31,35,31,133,31,175,31,245,31,245,30,245,29,211,31,211,30,208,31,176,31,237,31,237,30,34,31,47,31,47,30,29,31,240,31,75,31,81,31,81,30,81,29,2,31,192,31,187,31,187,30,34,31,165,31,175,31,239,31,163,31,135,31,244,31,170,31,170,30,130,31,230,31,230,30,207,31,133,31,59,31,56,31,232,31,247,31,45,31,136,31,41,31,255,31,255,30,146,31,109,31,159,31,1,31,240,31,37,31,208,31,84,31,147,31,227,31,227,30,182,31,182,30,182,31,182,30,229,31,36,31,249,31,173,31,54,31,54,30,120,31,147,31,166,31,38,31,101,31,254,31,30,31,20,31,239,31,66,31,19,31,139,31,126,31,20,31,20,30,59,31,240,31,217,31,174,31,226,31,171,31,167,31,200,31,200,30,255,31,63,31,96,31,221,31,44,31,84,31,237,31,237,30,205,31,205,30,205,29,96,31,96,30,179,31,198,31,102,31,198,31,15,31,15,30,15,29,98,31,16,31,251,31,40,31,29,31,29,30,33,31,173,31,33,31,92,31,92,30,24,31,200,31,89,31,37,31,117,31,223,31,180,31,33,31,145,31,71,31,176,31,209,31,4,31,4,30,85,31,153,31,153,30,153,29,54,31,178,31,96,31,2,31,246,31,173,31,21,31,10,31,43,31,248,31,160,31,90,31,158,31,204,31,56,31,15,31,120,31,120,30,74,31,57,31,57,30,121,31,186,31,251,31,92,31,70,31,70,30,20,31,215,31,215,30,215,29,248,31,30,31,153,31,153,30,37,31,37,30,37,29,252,31,128,31,128,31,34,31,26,31,64,31,18,31,184,31,176,31,53,31,22,31,22,30,143,31,16,31,16,30,124,31,113,31,89,31,168,31,25,31,49,31,136,31,168,31,227,31,105,31,200,31,11,31,11,30,11,31,160,31,186,31,248,31,248,30,135,31,238,31,244,31,66,31,163,31,113,31,12,31,250,31,250,30,250,29,7,31,39,31,6,31,43,31,114,31,223,31,179,31,106,31,200,31,138,31,138,30,33,31,9,31,209,31,174,31,176,31,16,31,36,31,121,31,224,31,149,31,213,31,181,31,78,31,197,31,197,30,42,31,7,31,252,31,164,31,115,31,115,30,154,31,177,31,133,31,133,30,204,31,192,31,192,30,221,31,225,31,48,31,48,30,192,31,192,30,137,31,55,31,218,31,254,31,182,31,25,31,229,31,233,31,175,31,99,31,97,31,217,31,36,31,116,31,42,31,53,31,153,31,134,31,134,30,249,31,145,31,145,30,184,31,99,31,120,31,19,31,239,31,47,31,75,31,75,30,140,31,90,31,81,31,121,31,66,31,161,31,158,31,158,30,158,29,173,31,173,30,248,31,244,31,196,31,19,31,19,30,51,31,51,30,51,29,24,31,24,30,248,31,104,31,107,31,63,31,71,31,21,31,21,30,52,31,177,31,67,31,67,30,232,31,146,31,53,31,2,31,191,31,114,31,114,30,114,29,13,31,31,31,233,31,19,31,147,31,174,31,86,31,28,31,242,31,223,31,221,31,166,31,254,31,254,30,59,31,59,30,171,31,175,31,145,31,130,31,65,31,1,31,178,31,239,31,239,30,145,31,153,31,243,31,243,30,158,31,145,31,192,31,5,31,157,31,160,31,160,30,132,31,27,31,113,31,102,31,113,31,11,31,11,30,44,31,44,30,44,29,44,28,82,31,69,31,225,31,136,31,160,31,160,30,63,31,196,31,137,31,48,31,66,31,135,31,22,31,22,30,22,29,51,31,51,30,125,31,209,31,33,31,33,30,65,31,175,31,120,31,164,31,10,31,202,31,202,30,27,31,225,31,190,31,65,31,65,30,91,31,167,31,127,31,4,31,92,31,154,31,41,31,194,31,178,31,209,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
