-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 969;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (90,0,103,0,0,0,0,0,0,0,74,0,151,0,21,0,14,0,152,0,0,0,104,0,0,0,97,0,182,0,0,0,0,0,18,0,178,0,0,0,0,0,68,0,17,0,245,0,0,0,10,0,48,0,177,0,10,0,184,0,132,0,242,0,192,0,0,0,55,0,193,0,231,0,0,0,108,0,39,0,97,0,198,0,0,0,222,0,75,0,67,0,179,0,0,0,0,0,140,0,140,0,12,0,212,0,213,0,0,0,0,0,227,0,41,0,102,0,18,0,0,0,0,0,45,0,73,0,0,0,42,0,51,0,0,0,145,0,182,0,138,0,151,0,120,0,237,0,67,0,1,0,157,0,0,0,204,0,145,0,90,0,83,0,4,0,149,0,134,0,252,0,106,0,155,0,0,0,0,0,0,0,251,0,0,0,1,0,0,0,103,0,0,0,2,0,243,0,161,0,111,0,46,0,73,0,72,0,121,0,69,0,255,0,146,0,13,0,220,0,224,0,0,0,76,0,212,0,223,0,152,0,0,0,37,0,0,0,191,0,0,0,158,0,154,0,124,0,26,0,169,0,23,0,52,0,129,0,73,0,32,0,236,0,0,0,92,0,240,0,228,0,194,0,182,0,98,0,0,0,0,0,0,0,124,0,235,0,0,0,175,0,190,0,163,0,236,0,174,0,141,0,38,0,11,0,0,0,154,0,204,0,0,0,254,0,0,0,25,0,229,0,0,0,146,0,0,0,131,0,165,0,142,0,227,0,242,0,81,0,31,0,255,0,246,0,148,0,77,0,68,0,133,0,37,0,116,0,91,0,0,0,0,0,193,0,92,0,220,0,237,0,0,0,89,0,74,0,233,0,142,0,204,0,205,0,0,0,26,0,148,0,129,0,117,0,27,0,34,0,206,0,175,0,139,0,98,0,231,0,145,0,152,0,230,0,75,0,130,0,135,0,0,0,0,0,67,0,185,0,1,0,0,0,13,0,0,0,58,0,235,0,33,0,131,0,62,0,137,0,247,0,144,0,0,0,143,0,88,0,211,0,253,0,0,0,166,0,180,0,160,0,192,0,230,0,0,0,0,0,0,0,54,0,55,0,75,0,125,0,135,0,0,0,168,0,221,0,177,0,180,0,167,0,249,0,97,0,0,0,0,0,162,0,14,0,80,0,126,0,0,0,237,0,143,0,87,0,215,0,0,0,47,0,24,0,0,0,46,0,138,0,5,0,99,0,139,0,0,0,141,0,83,0,181,0,88,0,218,0,0,0,172,0,57,0,136,0,224,0,0,0,2,0,0,0,150,0,243,0,0,0,0,0,151,0,84,0,0,0,201,0,169,0,246,0,121,0,85,0,147,0,27,0,176,0,0,0,23,0,0,0,209,0,248,0,0,0,0,0,41,0,205,0,220,0,101,0,116,0,119,0,49,0,98,0,93,0,95,0,0,0,114,0,225,0,7,0,131,0,245,0,243,0,0,0,189,0,222,0,69,0,148,0,97,0,168,0,67,0,112,0,56,0,160,0,106,0,208,0,123,0,209,0,169,0,211,0,144,0,6,0,0,0,228,0,167,0,0,0,228,0,93,0,166,0,58,0,145,0,137,0,23,0,34,0,197,0,0,0,177,0,226,0,219,0,234,0,99,0,0,0,0,0,215,0,111,0,28,0,242,0,13,0,96,0,109,0,36,0,230,0,191,0,136,0,120,0,73,0,209,0,160,0,113,0,174,0,0,0,54,0,142,0,50,0,157,0,174,0,13,0,247,0,97,0,199,0,111,0,117,0,231,0,0,0,5,0,169,0,63,0,143,0,253,0,169,0,93,0,218,0,169,0,92,0,0,0,129,0,200,0,220,0,0,0,183,0,42,0,192,0,0,0,81,0,0,0,11,0,214,0,156,0,79,0,137,0,16,0,108,0,255,0,0,0,9,0,181,0,1,0,59,0,45,0,1,0,175,0,189,0,229,0,10,0,131,0,0,0,172,0,148,0,199,0,0,0,87,0,140,0,193,0,136,0,250,0,180,0,238,0,75,0,211,0,0,0,210,0,255,0,200,0,172,0,174,0,196,0,78,0,36,0,39,0,0,0,140,0,187,0,0,0,7,0,136,0,140,0,107,0,145,0,156,0,156,0,81,0,181,0,252,0,0,0,208,0,0,0,0,0,214,0,50,0,126,0,228,0,177,0,243,0,242,0,137,0,143,0,96,0,14,0,15,0,254,0,60,0,0,0,0,0,200,0,146,0,8,0,90,0,121,0,26,0,221,0,175,0,151,0,142,0,214,0,0,0,111,0,222,0,0,0,234,0,253,0,0,0,0,0,0,0,0,0,110,0,47,0,116,0,89,0,117,0,0,0,166,0,218,0,234,0,246,0,11,0,0,0,100,0,98,0,14,0,217,0,0,0,82,0,0,0,228,0,109,0,129,0,0,0,0,0,239,0,208,0,170,0,0,0,131,0,236,0,217,0,178,0,86,0,7,0,69,0,11,0,99,0,165,0,126,0,191,0,183,0,3,0,48,0,1,0,90,0,85,0,35,0,0,0,215,0,0,0,0,0,18,0,34,0,225,0,218,0,129,0,104,0,151,0,174,0,99,0,78,0,0,0,188,0,186,0,191,0,117,0,171,0,0,0,241,0,207,0,198,0,187,0,140,0,6,0,0,0,108,0,173,0,78,0,147,0,163,0,83,0,3,0,222,0,133,0,95,0,238,0,0,0,0,0,138,0,142,0,140,0,0,0,237,0,106,0,48,0,203,0,118,0,239,0,50,0,104,0,151,0,14,0,181,0,112,0,194,0,147,0,0,0,0,0,20,0,244,0,153,0,209,0,179,0,135,0,0,0,0,0,60,0,88,0,160,0,209,0,87,0,187,0,153,0,78,0,252,0,0,0,115,0,163,0,0,0,165,0,30,0,57,0,215,0,189,0,61,0,0,0,195,0,56,0,0,0,155,0,124,0,0,0,149,0,93,0,142,0,254,0,105,0,217,0,0,0,204,0,200,0,158,0,93,0,248,0,0,0,247,0,244,0,197,0,236,0,71,0,0,0,0,0,39,0,200,0,131,0,0,0,67,0,74,0,115,0,76,0,122,0,215,0,0,0,150,0,40,0,0,0,31,0,152,0,250,0,77,0,181,0,102,0,215,0,111,0,211,0,0,0,0,0,181,0,162,0,70,0,217,0,233,0,51,0,100,0,4,0,155,0,103,0,7,0,67,0,0,0,135,0,125,0,0,0,30,0,141,0,66,0,220,0,58,0,119,0,122,0,8,0,27,0,155,0,96,0,17,0,111,0,199,0,164,0,248,0,0,0,124,0,153,0,83,0,191,0,67,0,35,0,0,0,0,0,140,0,0,0,62,0,0,0,0,0,172,0,240,0,12,0,86,0,211,0,207,0,81,0,54,0,100,0,19,0,0,0,243,0,224,0,254,0,136,0,69,0,154,0,12,0,28,0,147,0,119,0,152,0,158,0,0,0,0,0,0,0,240,0,133,0,194,0,132,0,45,0,0,0,181,0,249,0,26,0,112,0,0,0,27,0,53,0,0,0,0,0,106,0,238,0,0,0,134,0,0,0,159,0,235,0,0,0,188,0,18,0,142,0,9,0,57,0,0,0,20,0,231,0,181,0,207,0,177,0,150,0,83,0,77,0,255,0,162,0,94,0,202,0,18,0,122,0,80,0,163,0,0,0,79,0,62,0,0,0,13,0,0,0,94,0,88,0,83,0,101,0,0,0,190,0,217,0,145,0,244,0,38,0,169,0,45,0,49,0,217,0,0,0,144,0,70,0,62,0,22,0,230,0,105,0,62,0,0,0,47,0,228,0,130,0,141,0,204,0,174,0,215,0,102,0,64,0,124,0,98,0,72,0,166,0,33,0,78,0,232,0,0,0,167,0,98,0,136,0,47,0,135,0,0,0,103,0,81,0,45,0,8,0,6,0,23,0,93,0,0,0,128,0,238,0,181,0,0,0,0,0,16,0,215,0,122,0,62,0,0,0,57,0,198,0,0,0,55,0,0,0,2,0,101,0,47,0,1,0,198,0,0,0,0,0,0,0,138,0,163,0,0,0,0,0,202,0,163,0,0,0,71,0,81,0,4,0,13,0,0,0,94,0,129,0,74,0,7,0,101,0,178,0,37,0,82,0,115,0,12,0,11,0,207,0,0,0,0,0,192,0,217,0,206,0,253,0,130,0,34,0,206,0,137,0,0,0,120,0,139,0,0,0,187,0,147,0,230,0,107,0,162,0,0,0,91,0,0,0,215,0,208,0,187,0,34,0,72,0,0,0,221,0,66,0,121,0,0,0,18,0,206,0,0,0,103,0,208,0,84,0,20,0,174,0);
signal scenario_full  : scenario_type := (90,31,103,31,103,30,103,29,103,28,74,31,151,31,21,31,14,31,152,31,152,30,104,31,104,30,97,31,182,31,182,30,182,29,18,31,178,31,178,30,178,29,68,31,17,31,245,31,245,30,10,31,48,31,177,31,10,31,184,31,132,31,242,31,192,31,192,30,55,31,193,31,231,31,231,30,108,31,39,31,97,31,198,31,198,30,222,31,75,31,67,31,179,31,179,30,179,29,140,31,140,31,12,31,212,31,213,31,213,30,213,29,227,31,41,31,102,31,18,31,18,30,18,29,45,31,73,31,73,30,42,31,51,31,51,30,145,31,182,31,138,31,151,31,120,31,237,31,67,31,1,31,157,31,157,30,204,31,145,31,90,31,83,31,4,31,149,31,134,31,252,31,106,31,155,31,155,30,155,29,155,28,251,31,251,30,1,31,1,30,103,31,103,30,2,31,243,31,161,31,111,31,46,31,73,31,72,31,121,31,69,31,255,31,146,31,13,31,220,31,224,31,224,30,76,31,212,31,223,31,152,31,152,30,37,31,37,30,191,31,191,30,158,31,154,31,124,31,26,31,169,31,23,31,52,31,129,31,73,31,32,31,236,31,236,30,92,31,240,31,228,31,194,31,182,31,98,31,98,30,98,29,98,28,124,31,235,31,235,30,175,31,190,31,163,31,236,31,174,31,141,31,38,31,11,31,11,30,154,31,204,31,204,30,254,31,254,30,25,31,229,31,229,30,146,31,146,30,131,31,165,31,142,31,227,31,242,31,81,31,31,31,255,31,246,31,148,31,77,31,68,31,133,31,37,31,116,31,91,31,91,30,91,29,193,31,92,31,220,31,237,31,237,30,89,31,74,31,233,31,142,31,204,31,205,31,205,30,26,31,148,31,129,31,117,31,27,31,34,31,206,31,175,31,139,31,98,31,231,31,145,31,152,31,230,31,75,31,130,31,135,31,135,30,135,29,67,31,185,31,1,31,1,30,13,31,13,30,58,31,235,31,33,31,131,31,62,31,137,31,247,31,144,31,144,30,143,31,88,31,211,31,253,31,253,30,166,31,180,31,160,31,192,31,230,31,230,30,230,29,230,28,54,31,55,31,75,31,125,31,135,31,135,30,168,31,221,31,177,31,180,31,167,31,249,31,97,31,97,30,97,29,162,31,14,31,80,31,126,31,126,30,237,31,143,31,87,31,215,31,215,30,47,31,24,31,24,30,46,31,138,31,5,31,99,31,139,31,139,30,141,31,83,31,181,31,88,31,218,31,218,30,172,31,57,31,136,31,224,31,224,30,2,31,2,30,150,31,243,31,243,30,243,29,151,31,84,31,84,30,201,31,169,31,246,31,121,31,85,31,147,31,27,31,176,31,176,30,23,31,23,30,209,31,248,31,248,30,248,29,41,31,205,31,220,31,101,31,116,31,119,31,49,31,98,31,93,31,95,31,95,30,114,31,225,31,7,31,131,31,245,31,243,31,243,30,189,31,222,31,69,31,148,31,97,31,168,31,67,31,112,31,56,31,160,31,106,31,208,31,123,31,209,31,169,31,211,31,144,31,6,31,6,30,228,31,167,31,167,30,228,31,93,31,166,31,58,31,145,31,137,31,23,31,34,31,197,31,197,30,177,31,226,31,219,31,234,31,99,31,99,30,99,29,215,31,111,31,28,31,242,31,13,31,96,31,109,31,36,31,230,31,191,31,136,31,120,31,73,31,209,31,160,31,113,31,174,31,174,30,54,31,142,31,50,31,157,31,174,31,13,31,247,31,97,31,199,31,111,31,117,31,231,31,231,30,5,31,169,31,63,31,143,31,253,31,169,31,93,31,218,31,169,31,92,31,92,30,129,31,200,31,220,31,220,30,183,31,42,31,192,31,192,30,81,31,81,30,11,31,214,31,156,31,79,31,137,31,16,31,108,31,255,31,255,30,9,31,181,31,1,31,59,31,45,31,1,31,175,31,189,31,229,31,10,31,131,31,131,30,172,31,148,31,199,31,199,30,87,31,140,31,193,31,136,31,250,31,180,31,238,31,75,31,211,31,211,30,210,31,255,31,200,31,172,31,174,31,196,31,78,31,36,31,39,31,39,30,140,31,187,31,187,30,7,31,136,31,140,31,107,31,145,31,156,31,156,31,81,31,181,31,252,31,252,30,208,31,208,30,208,29,214,31,50,31,126,31,228,31,177,31,243,31,242,31,137,31,143,31,96,31,14,31,15,31,254,31,60,31,60,30,60,29,200,31,146,31,8,31,90,31,121,31,26,31,221,31,175,31,151,31,142,31,214,31,214,30,111,31,222,31,222,30,234,31,253,31,253,30,253,29,253,28,253,27,110,31,47,31,116,31,89,31,117,31,117,30,166,31,218,31,234,31,246,31,11,31,11,30,100,31,98,31,14,31,217,31,217,30,82,31,82,30,228,31,109,31,129,31,129,30,129,29,239,31,208,31,170,31,170,30,131,31,236,31,217,31,178,31,86,31,7,31,69,31,11,31,99,31,165,31,126,31,191,31,183,31,3,31,48,31,1,31,90,31,85,31,35,31,35,30,215,31,215,30,215,29,18,31,34,31,225,31,218,31,129,31,104,31,151,31,174,31,99,31,78,31,78,30,188,31,186,31,191,31,117,31,171,31,171,30,241,31,207,31,198,31,187,31,140,31,6,31,6,30,108,31,173,31,78,31,147,31,163,31,83,31,3,31,222,31,133,31,95,31,238,31,238,30,238,29,138,31,142,31,140,31,140,30,237,31,106,31,48,31,203,31,118,31,239,31,50,31,104,31,151,31,14,31,181,31,112,31,194,31,147,31,147,30,147,29,20,31,244,31,153,31,209,31,179,31,135,31,135,30,135,29,60,31,88,31,160,31,209,31,87,31,187,31,153,31,78,31,252,31,252,30,115,31,163,31,163,30,165,31,30,31,57,31,215,31,189,31,61,31,61,30,195,31,56,31,56,30,155,31,124,31,124,30,149,31,93,31,142,31,254,31,105,31,217,31,217,30,204,31,200,31,158,31,93,31,248,31,248,30,247,31,244,31,197,31,236,31,71,31,71,30,71,29,39,31,200,31,131,31,131,30,67,31,74,31,115,31,76,31,122,31,215,31,215,30,150,31,40,31,40,30,31,31,152,31,250,31,77,31,181,31,102,31,215,31,111,31,211,31,211,30,211,29,181,31,162,31,70,31,217,31,233,31,51,31,100,31,4,31,155,31,103,31,7,31,67,31,67,30,135,31,125,31,125,30,30,31,141,31,66,31,220,31,58,31,119,31,122,31,8,31,27,31,155,31,96,31,17,31,111,31,199,31,164,31,248,31,248,30,124,31,153,31,83,31,191,31,67,31,35,31,35,30,35,29,140,31,140,30,62,31,62,30,62,29,172,31,240,31,12,31,86,31,211,31,207,31,81,31,54,31,100,31,19,31,19,30,243,31,224,31,254,31,136,31,69,31,154,31,12,31,28,31,147,31,119,31,152,31,158,31,158,30,158,29,158,28,240,31,133,31,194,31,132,31,45,31,45,30,181,31,249,31,26,31,112,31,112,30,27,31,53,31,53,30,53,29,106,31,238,31,238,30,134,31,134,30,159,31,235,31,235,30,188,31,18,31,142,31,9,31,57,31,57,30,20,31,231,31,181,31,207,31,177,31,150,31,83,31,77,31,255,31,162,31,94,31,202,31,18,31,122,31,80,31,163,31,163,30,79,31,62,31,62,30,13,31,13,30,94,31,88,31,83,31,101,31,101,30,190,31,217,31,145,31,244,31,38,31,169,31,45,31,49,31,217,31,217,30,144,31,70,31,62,31,22,31,230,31,105,31,62,31,62,30,47,31,228,31,130,31,141,31,204,31,174,31,215,31,102,31,64,31,124,31,98,31,72,31,166,31,33,31,78,31,232,31,232,30,167,31,98,31,136,31,47,31,135,31,135,30,103,31,81,31,45,31,8,31,6,31,23,31,93,31,93,30,128,31,238,31,181,31,181,30,181,29,16,31,215,31,122,31,62,31,62,30,57,31,198,31,198,30,55,31,55,30,2,31,101,31,47,31,1,31,198,31,198,30,198,29,198,28,138,31,163,31,163,30,163,29,202,31,163,31,163,30,71,31,81,31,4,31,13,31,13,30,94,31,129,31,74,31,7,31,101,31,178,31,37,31,82,31,115,31,12,31,11,31,207,31,207,30,207,29,192,31,217,31,206,31,253,31,130,31,34,31,206,31,137,31,137,30,120,31,139,31,139,30,187,31,147,31,230,31,107,31,162,31,162,30,91,31,91,30,215,31,208,31,187,31,34,31,72,31,72,30,221,31,66,31,121,31,121,30,18,31,206,31,206,30,103,31,208,31,84,31,20,31,174,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
