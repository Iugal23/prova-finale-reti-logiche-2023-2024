-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 194;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (36,0,149,0,0,0,134,0,191,0,182,0,249,0,90,0,183,0,92,0,131,0,148,0,99,0,138,0,47,0,209,0,198,0,45,0,58,0,0,0,206,0,71,0,3,0,156,0,162,0,179,0,212,0,84,0,174,0,9,0,0,0,67,0,102,0,52,0,0,0,220,0,206,0,120,0,106,0,0,0,47,0,217,0,180,0,0,0,45,0,241,0,0,0,228,0,156,0,207,0,146,0,17,0,0,0,59,0,140,0,0,0,217,0,129,0,237,0,62,0,68,0,141,0,17,0,94,0,120,0,154,0,0,0,108,0,166,0,127,0,246,0,0,0,191,0,30,0,88,0,232,0,158,0,235,0,245,0,26,0,51,0,36,0,75,0,154,0,205,0,189,0,0,0,229,0,8,0,51,0,217,0,15,0,98,0,145,0,35,0,64,0,77,0,78,0,78,0,30,0,209,0,0,0,0,0,19,0,193,0,6,0,108,0,214,0,242,0,234,0,51,0,17,0,96,0,221,0,7,0,252,0,0,0,102,0,137,0,239,0,2,0,167,0,144,0,0,0,94,0,0,0,145,0,233,0,121,0,232,0,178,0,0,0,243,0,113,0,13,0,189,0,27,0,239,0,187,0,163,0,0,0,0,0,0,0,244,0,171,0,83,0,0,0,61,0,143,0,154,0,0,0,23,0,0,0,0,0,233,0,87,0,228,0,240,0,11,0,70,0,0,0,235,0,217,0,140,0,222,0,111,0,0,0,215,0,165,0,0,0,83,0,130,0,57,0,18,0,152,0,174,0,105,0,241,0,209,0,183,0,76,0,143,0,216,0,209,0,218,0,182,0,0,0,56,0,34,0,237,0,0,0,21,0,0,0,78,0);
signal scenario_full  : scenario_type := (36,31,149,31,149,30,134,31,191,31,182,31,249,31,90,31,183,31,92,31,131,31,148,31,99,31,138,31,47,31,209,31,198,31,45,31,58,31,58,30,206,31,71,31,3,31,156,31,162,31,179,31,212,31,84,31,174,31,9,31,9,30,67,31,102,31,52,31,52,30,220,31,206,31,120,31,106,31,106,30,47,31,217,31,180,31,180,30,45,31,241,31,241,30,228,31,156,31,207,31,146,31,17,31,17,30,59,31,140,31,140,30,217,31,129,31,237,31,62,31,68,31,141,31,17,31,94,31,120,31,154,31,154,30,108,31,166,31,127,31,246,31,246,30,191,31,30,31,88,31,232,31,158,31,235,31,245,31,26,31,51,31,36,31,75,31,154,31,205,31,189,31,189,30,229,31,8,31,51,31,217,31,15,31,98,31,145,31,35,31,64,31,77,31,78,31,78,31,30,31,209,31,209,30,209,29,19,31,193,31,6,31,108,31,214,31,242,31,234,31,51,31,17,31,96,31,221,31,7,31,252,31,252,30,102,31,137,31,239,31,2,31,167,31,144,31,144,30,94,31,94,30,145,31,233,31,121,31,232,31,178,31,178,30,243,31,113,31,13,31,189,31,27,31,239,31,187,31,163,31,163,30,163,29,163,28,244,31,171,31,83,31,83,30,61,31,143,31,154,31,154,30,23,31,23,30,23,29,233,31,87,31,228,31,240,31,11,31,70,31,70,30,235,31,217,31,140,31,222,31,111,31,111,30,215,31,165,31,165,30,83,31,130,31,57,31,18,31,152,31,174,31,105,31,241,31,209,31,183,31,76,31,143,31,216,31,209,31,218,31,182,31,182,30,56,31,34,31,237,31,237,30,21,31,21,30,78,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
