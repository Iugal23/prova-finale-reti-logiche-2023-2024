-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_876 is
end project_tb_876;

architecture project_tb_arch_876 of project_tb_876 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 568;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,160,0,171,0,0,0,123,0,136,0,205,0,128,0,166,0,244,0,3,0,0,0,218,0,206,0,247,0,0,0,109,0,175,0,99,0,220,0,155,0,103,0,193,0,23,0,133,0,115,0,182,0,28,0,129,0,45,0,77,0,145,0,118,0,60,0,224,0,210,0,172,0,0,0,41,0,0,0,222,0,190,0,137,0,45,0,58,0,251,0,43,0,54,0,215,0,0,0,233,0,175,0,127,0,0,0,50,0,251,0,227,0,50,0,165,0,252,0,229,0,231,0,46,0,189,0,79,0,0,0,193,0,189,0,22,0,167,0,21,0,191,0,165,0,122,0,0,0,33,0,99,0,254,0,71,0,83,0,74,0,189,0,64,0,66,0,80,0,39,0,80,0,38,0,113,0,64,0,40,0,66,0,188,0,137,0,195,0,101,0,190,0,145,0,251,0,112,0,252,0,37,0,1,0,0,0,201,0,153,0,163,0,5,0,77,0,66,0,97,0,72,0,0,0,3,0,99,0,43,0,28,0,101,0,166,0,251,0,226,0,84,0,127,0,113,0,0,0,172,0,66,0,163,0,233,0,27,0,96,0,232,0,210,0,86,0,0,0,211,0,232,0,0,0,171,0,192,0,24,0,101,0,84,0,1,0,16,0,0,0,0,0,0,0,232,0,0,0,106,0,141,0,152,0,0,0,211,0,0,0,25,0,0,0,14,0,0,0,0,0,20,0,0,0,98,0,79,0,0,0,0,0,177,0,40,0,55,0,96,0,20,0,99,0,83,0,47,0,127,0,163,0,228,0,0,0,0,0,23,0,83,0,39,0,242,0,190,0,72,0,0,0,121,0,106,0,199,0,153,0,161,0,0,0,0,0,228,0,47,0,105,0,72,0,38,0,216,0,174,0,0,0,0,0,0,0,127,0,134,0,58,0,159,0,18,0,255,0,187,0,219,0,184,0,0,0,0,0,71,0,0,0,0,0,211,0,0,0,173,0,105,0,105,0,0,0,0,0,36,0,198,0,171,0,0,0,0,0,0,0,134,0,0,0,240,0,251,0,0,0,222,0,0,0,248,0,216,0,204,0,93,0,0,0,0,0,0,0,166,0,41,0,0,0,49,0,0,0,228,0,0,0,211,0,0,0,0,0,223,0,0,0,101,0,0,0,222,0,0,0,92,0,105,0,120,0,108,0,239,0,51,0,0,0,196,0,249,0,243,0,253,0,144,0,101,0,175,0,0,0,31,0,0,0,10,0,163,0,52,0,0,0,157,0,127,0,0,0,172,0,247,0,212,0,101,0,22,0,163,0,16,0,225,0,101,0,26,0,251,0,0,0,138,0,84,0,250,0,183,0,248,0,0,0,114,0,0,0,66,0,51,0,0,0,203,0,0,0,115,0,4,0,154,0,2,0,160,0,132,0,215,0,173,0,209,0,0,0,82,0,0,0,231,0,204,0,42,0,89,0,187,0,31,0,95,0,0,0,11,0,148,0,159,0,165,0,0,0,216,0,116,0,100,0,116,0,184,0,0,0,239,0,18,0,0,0,63,0,250,0,85,0,61,0,167,0,100,0,244,0,0,0,0,0,62,0,0,0,40,0,222,0,0,0,41,0,141,0,211,0,106,0,40,0,119,0,182,0,116,0,252,0,99,0,0,0,219,0,98,0,87,0,200,0,0,0,55,0,161,0,197,0,0,0,101,0,195,0,78,0,133,0,164,0,197,0,0,0,139,0,224,0,0,0,143,0,67,0,80,0,143,0,44,0,91,0,191,0,18,0,0,0,0,0,75,0,38,0,0,0,137,0,0,0,244,0,0,0,38,0,240,0,0,0,77,0,20,0,0,0,51,0,113,0,189,0,149,0,127,0,97,0,218,0,48,0,0,0,0,0,215,0,109,0,0,0,176,0,253,0,0,0,193,0,0,0,21,0,164,0,73,0,50,0,74,0,0,0,151,0,109,0,124,0,0,0,0,0,0,0,0,0,104,0,133,0,115,0,233,0,89,0,222,0,0,0,185,0,138,0,213,0,197,0,185,0,82,0,22,0,0,0,110,0,0,0,17,0,0,0,0,0,0,0,72,0,0,0,108,0,21,0,139,0,0,0,110,0,80,0,19,0,0,0,153,0,219,0,61,0,0,0,224,0,128,0,119,0,69,0,0,0,39,0,0,0,195,0,58,0,225,0,51,0,87,0,0,0,174,0,0,0,139,0,95,0,0,0,23,0,68,0,0,0,0,0,70,0,156,0,190,0,74,0,197,0,0,0,228,0,186,0,215,0,135,0,50,0,0,0,0,0,50,0,0,0,68,0,0,0,41,0,66,0,148,0,32,0,185,0,131,0,44,0,31,0,0,0,0,0,164,0,1,0,239,0,52,0,216,0,28,0,143,0,36,0,6,0,102,0,75,0,12,0,66,0,78,0,24,0,153,0,95,0,47,0,241,0,42,0,45,0,56,0,19,0,113,0,105,0,198,0,65,0,20,0,168,0,134,0,194,0,166,0,81,0,137,0,214,0,210,0,250,0,0,0,0,0,174,0,85,0,54,0);
signal scenario_full  : scenario_type := (0,0,160,31,171,31,171,30,123,31,136,31,205,31,128,31,166,31,244,31,3,31,3,30,218,31,206,31,247,31,247,30,109,31,175,31,99,31,220,31,155,31,103,31,193,31,23,31,133,31,115,31,182,31,28,31,129,31,45,31,77,31,145,31,118,31,60,31,224,31,210,31,172,31,172,30,41,31,41,30,222,31,190,31,137,31,45,31,58,31,251,31,43,31,54,31,215,31,215,30,233,31,175,31,127,31,127,30,50,31,251,31,227,31,50,31,165,31,252,31,229,31,231,31,46,31,189,31,79,31,79,30,193,31,189,31,22,31,167,31,21,31,191,31,165,31,122,31,122,30,33,31,99,31,254,31,71,31,83,31,74,31,189,31,64,31,66,31,80,31,39,31,80,31,38,31,113,31,64,31,40,31,66,31,188,31,137,31,195,31,101,31,190,31,145,31,251,31,112,31,252,31,37,31,1,31,1,30,201,31,153,31,163,31,5,31,77,31,66,31,97,31,72,31,72,30,3,31,99,31,43,31,28,31,101,31,166,31,251,31,226,31,84,31,127,31,113,31,113,30,172,31,66,31,163,31,233,31,27,31,96,31,232,31,210,31,86,31,86,30,211,31,232,31,232,30,171,31,192,31,24,31,101,31,84,31,1,31,16,31,16,30,16,29,16,28,232,31,232,30,106,31,141,31,152,31,152,30,211,31,211,30,25,31,25,30,14,31,14,30,14,29,20,31,20,30,98,31,79,31,79,30,79,29,177,31,40,31,55,31,96,31,20,31,99,31,83,31,47,31,127,31,163,31,228,31,228,30,228,29,23,31,83,31,39,31,242,31,190,31,72,31,72,30,121,31,106,31,199,31,153,31,161,31,161,30,161,29,228,31,47,31,105,31,72,31,38,31,216,31,174,31,174,30,174,29,174,28,127,31,134,31,58,31,159,31,18,31,255,31,187,31,219,31,184,31,184,30,184,29,71,31,71,30,71,29,211,31,211,30,173,31,105,31,105,31,105,30,105,29,36,31,198,31,171,31,171,30,171,29,171,28,134,31,134,30,240,31,251,31,251,30,222,31,222,30,248,31,216,31,204,31,93,31,93,30,93,29,93,28,166,31,41,31,41,30,49,31,49,30,228,31,228,30,211,31,211,30,211,29,223,31,223,30,101,31,101,30,222,31,222,30,92,31,105,31,120,31,108,31,239,31,51,31,51,30,196,31,249,31,243,31,253,31,144,31,101,31,175,31,175,30,31,31,31,30,10,31,163,31,52,31,52,30,157,31,127,31,127,30,172,31,247,31,212,31,101,31,22,31,163,31,16,31,225,31,101,31,26,31,251,31,251,30,138,31,84,31,250,31,183,31,248,31,248,30,114,31,114,30,66,31,51,31,51,30,203,31,203,30,115,31,4,31,154,31,2,31,160,31,132,31,215,31,173,31,209,31,209,30,82,31,82,30,231,31,204,31,42,31,89,31,187,31,31,31,95,31,95,30,11,31,148,31,159,31,165,31,165,30,216,31,116,31,100,31,116,31,184,31,184,30,239,31,18,31,18,30,63,31,250,31,85,31,61,31,167,31,100,31,244,31,244,30,244,29,62,31,62,30,40,31,222,31,222,30,41,31,141,31,211,31,106,31,40,31,119,31,182,31,116,31,252,31,99,31,99,30,219,31,98,31,87,31,200,31,200,30,55,31,161,31,197,31,197,30,101,31,195,31,78,31,133,31,164,31,197,31,197,30,139,31,224,31,224,30,143,31,67,31,80,31,143,31,44,31,91,31,191,31,18,31,18,30,18,29,75,31,38,31,38,30,137,31,137,30,244,31,244,30,38,31,240,31,240,30,77,31,20,31,20,30,51,31,113,31,189,31,149,31,127,31,97,31,218,31,48,31,48,30,48,29,215,31,109,31,109,30,176,31,253,31,253,30,193,31,193,30,21,31,164,31,73,31,50,31,74,31,74,30,151,31,109,31,124,31,124,30,124,29,124,28,124,27,104,31,133,31,115,31,233,31,89,31,222,31,222,30,185,31,138,31,213,31,197,31,185,31,82,31,22,31,22,30,110,31,110,30,17,31,17,30,17,29,17,28,72,31,72,30,108,31,21,31,139,31,139,30,110,31,80,31,19,31,19,30,153,31,219,31,61,31,61,30,224,31,128,31,119,31,69,31,69,30,39,31,39,30,195,31,58,31,225,31,51,31,87,31,87,30,174,31,174,30,139,31,95,31,95,30,23,31,68,31,68,30,68,29,70,31,156,31,190,31,74,31,197,31,197,30,228,31,186,31,215,31,135,31,50,31,50,30,50,29,50,31,50,30,68,31,68,30,41,31,66,31,148,31,32,31,185,31,131,31,44,31,31,31,31,30,31,29,164,31,1,31,239,31,52,31,216,31,28,31,143,31,36,31,6,31,102,31,75,31,12,31,66,31,78,31,24,31,153,31,95,31,47,31,241,31,42,31,45,31,56,31,19,31,113,31,105,31,198,31,65,31,20,31,168,31,134,31,194,31,166,31,81,31,137,31,214,31,210,31,250,31,250,30,250,29,174,31,85,31,54,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
