-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_600 is
end project_tb_600;

architecture project_tb_arch_600 of project_tb_600 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1021;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (228,0,0,0,193,0,118,0,26,0,85,0,71,0,0,0,170,0,202,0,76,0,0,0,159,0,153,0,35,0,226,0,213,0,36,0,80,0,0,0,125,0,19,0,27,0,0,0,24,0,224,0,170,0,0,0,183,0,39,0,130,0,188,0,237,0,223,0,127,0,0,0,100,0,16,0,107,0,6,0,120,0,34,0,0,0,170,0,0,0,0,0,0,0,96,0,144,0,185,0,152,0,159,0,154,0,30,0,210,0,103,0,0,0,32,0,242,0,55,0,242,0,231,0,118,0,246,0,0,0,44,0,145,0,120,0,0,0,188,0,13,0,0,0,0,0,162,0,86,0,97,0,0,0,85,0,198,0,0,0,0,0,175,0,110,0,0,0,203,0,0,0,249,0,249,0,237,0,0,0,30,0,0,0,0,0,202,0,222,0,184,0,0,0,136,0,0,0,0,0,93,0,107,0,46,0,33,0,0,0,170,0,0,0,217,0,239,0,0,0,0,0,0,0,108,0,231,0,2,0,244,0,0,0,221,0,121,0,44,0,103,0,247,0,193,0,0,0,203,0,211,0,209,0,235,0,249,0,58,0,78,0,20,0,28,0,176,0,156,0,244,0,0,0,83,0,103,0,0,0,208,0,150,0,60,0,18,0,139,0,0,0,25,0,226,0,66,0,112,0,48,0,0,0,230,0,240,0,189,0,0,0,50,0,0,0,254,0,121,0,0,0,107,0,166,0,163,0,90,0,180,0,19,0,227,0,88,0,218,0,159,0,240,0,30,0,66,0,0,0,99,0,107,0,32,0,167,0,150,0,243,0,179,0,170,0,29,0,74,0,0,0,175,0,178,0,0,0,205,0,148,0,0,0,160,0,0,0,140,0,223,0,0,0,53,0,57,0,154,0,0,0,70,0,141,0,78,0,135,0,31,0,0,0,92,0,197,0,223,0,236,0,0,0,146,0,0,0,0,0,248,0,20,0,183,0,0,0,87,0,200,0,19,0,23,0,215,0,104,0,183,0,129,0,228,0,132,0,206,0,0,0,225,0,64,0,0,0,110,0,102,0,12,0,0,0,194,0,0,0,0,0,27,0,47,0,97,0,203,0,162,0,214,0,2,0,146,0,8,0,93,0,255,0,105,0,90,0,0,0,168,0,167,0,155,0,124,0,186,0,44,0,45,0,19,0,148,0,163,0,11,0,176,0,182,0,114,0,40,0,0,0,85,0,199,0,0,0,161,0,48,0,186,0,109,0,42,0,108,0,130,0,46,0,249,0,0,0,0,0,210,0,77,0,0,0,0,0,211,0,155,0,0,0,115,0,0,0,236,0,117,0,210,0,67,0,132,0,47,0,78,0,195,0,121,0,87,0,0,0,169,0,107,0,115,0,209,0,162,0,53,0,111,0,86,0,250,0,63,0,34,0,26,0,45,0,209,0,108,0,87,0,10,0,121,0,145,0,242,0,0,0,0,0,181,0,118,0,131,0,120,0,254,0,0,0,16,0,71,0,186,0,244,0,64,0,240,0,28,0,219,0,121,0,146,0,124,0,185,0,31,0,108,0,123,0,91,0,240,0,119,0,106,0,7,0,147,0,26,0,0,0,124,0,26,0,91,0,66,0,0,0,71,0,255,0,200,0,0,0,255,0,138,0,98,0,212,0,25,0,159,0,9,0,64,0,247,0,167,0,8,0,51,0,162,0,75,0,153,0,0,0,102,0,165,0,123,0,130,0,214,0,190,0,102,0,0,0,91,0,0,0,0,0,205,0,19,0,163,0,66,0,167,0,16,0,150,0,141,0,101,0,0,0,0,0,0,0,95,0,109,0,179,0,26,0,202,0,144,0,29,0,132,0,121,0,94,0,0,0,246,0,102,0,0,0,0,0,110,0,42,0,133,0,34,0,219,0,177,0,74,0,126,0,129,0,0,0,0,0,0,0,0,0,0,0,13,0,63,0,99,0,105,0,97,0,221,0,192,0,124,0,110,0,149,0,37,0,81,0,0,0,157,0,130,0,0,0,0,0,0,0,87,0,0,0,0,0,145,0,195,0,125,0,42,0,162,0,0,0,0,0,110,0,0,0,87,0,25,0,130,0,200,0,110,0,0,0,0,0,174,0,0,0,0,0,0,0,245,0,75,0,0,0,69,0,197,0,174,0,0,0,110,0,167,0,93,0,60,0,94,0,23,0,94,0,212,0,240,0,215,0,0,0,140,0,0,0,0,0,190,0,223,0,0,0,0,0,61,0,215,0,0,0,175,0,190,0,194,0,90,0,28,0,45,0,110,0,0,0,107,0,130,0,139,0,212,0,186,0,194,0,82,0,121,0,0,0,139,0,24,0,83,0,28,0,88,0,0,0,164,0,222,0,224,0,0,0,247,0,155,0,0,0,163,0,1,0,192,0,126,0,109,0,1,0,9,0,167,0,31,0,186,0,216,0,231,0,224,0,153,0,200,0,186,0,0,0,86,0,62,0,37,0,0,0,212,0,0,0,207,0,114,0,18,0,0,0,0,0,6,0,136,0,0,0,118,0,136,0,0,0,0,0,143,0,0,0,94,0,59,0,73,0,102,0,0,0,87,0,0,0,171,0,0,0,0,0,199,0,171,0,44,0,254,0,47,0,114,0,59,0,0,0,68,0,0,0,33,0,55,0,0,0,48,0,215,0,120,0,47,0,13,0,0,0,133,0,150,0,199,0,86,0,244,0,211,0,93,0,151,0,93,0,37,0,114,0,173,0,45,0,0,0,29,0,184,0,0,0,68,0,82,0,171,0,104,0,190,0,0,0,170,0,164,0,243,0,251,0,36,0,82,0,56,0,0,0,9,0,38,0,137,0,0,0,165,0,0,0,176,0,173,0,158,0,64,0,0,0,53,0,119,0,71,0,168,0,30,0,131,0,59,0,191,0,224,0,103,0,255,0,169,0,149,0,107,0,199,0,97,0,14,0,210,0,114,0,150,0,143,0,0,0,187,0,200,0,70,0,76,0,0,0,23,0,224,0,178,0,191,0,0,0,122,0,167,0,0,0,13,0,97,0,212,0,0,0,109,0,69,0,213,0,247,0,71,0,0,0,219,0,35,0,0,0,27,0,166,0,16,0,0,0,77,0,184,0,244,0,42,0,124,0,0,0,40,0,128,0,180,0,19,0,61,0,33,0,216,0,0,0,128,0,0,0,141,0,26,0,191,0,201,0,158,0,85,0,98,0,11,0,127,0,0,0,203,0,234,0,217,0,109,0,0,0,106,0,111,0,0,0,15,0,7,0,239,0,6,0,164,0,173,0,182,0,0,0,84,0,38,0,0,0,0,0,127,0,0,0,72,0,0,0,29,0,83,0,129,0,101,0,204,0,0,0,135,0,176,0,34,0,0,0,218,0,0,0,25,0,16,0,166,0,0,0,107,0,0,0,38,0,0,0,106,0,0,0,0,0,143,0,35,0,177,0,206,0,0,0,40,0,0,0,0,0,154,0,8,0,15,0,98,0,57,0,93,0,186,0,127,0,190,0,0,0,0,0,174,0,249,0,132,0,0,0,0,0,170,0,8,0,214,0,0,0,0,0,22,0,0,0,212,0,0,0,13,0,77,0,0,0,110,0,195,0,145,0,0,0,4,0,94,0,51,0,47,0,0,0,164,0,31,0,254,0,0,0,160,0,103,0,36,0,0,0,22,0,218,0,163,0,125,0,115,0,106,0,30,0,203,0,49,0,255,0,19,0,169,0,61,0,57,0,163,0,115,0,97,0,121,0,46,0,141,0,38,0,0,0,223,0,11,0,0,0,190,0,133,0,0,0,0,0,220,0,50,0,95,0,246,0,29,0,0,0,230,0,0,0,153,0,32,0,0,0,92,0,153,0,0,0,249,0,114,0,0,0,145,0,100,0,0,0,2,0,162,0,0,0,0,0,225,0,139,0,202,0,42,0,231,0,0,0,180,0,178,0,24,0,253,0,242,0,102,0,47,0,20,0,156,0,178,0,219,0,0,0,127,0,0,0,0,0,0,0,102,0,10,0,212,0,174,0,0,0,0,0,237,0,199,0,9,0,0,0,248,0,10,0,0,0,133,0,181,0,122,0,177,0,56,0,11,0,93,0,132,0,252,0,0,0,155,0,60,0,69,0,193,0,226,0,23,0,52,0,0,0,247,0,0,0,137,0,2,0,72,0,0,0,14,0,119,0,25,0,0,0,139,0,118,0,166,0,0,0,19,0,124,0,174,0,103,0,22,0,100,0,0,0,72,0,213,0,103,0,111,0,75,0,149,0,46,0,66,0,50,0,112,0,34,0,107,0,221,0,200,0,80,0,25,0,0,0,80,0,109,0,152,0,171,0,116,0,0,0,200,0,147,0,7,0,51,0,153,0,0,0,0,0,0,0,0,0,189,0,1,0,0,0,172,0,189,0,140,0,103,0,150,0,5,0,31,0,108,0,100,0,49,0,215,0,0,0,0,0,244,0,203,0,155,0,200,0,201,0,0,0,119,0,235,0,222,0,0,0,183,0,0,0,31,0,237,0,8,0,0,0,146,0,194,0,63,0,221,0,141,0,73,0,36,0,30,0,109,0,0,0,222,0,126,0);
signal scenario_full  : scenario_type := (228,31,228,30,193,31,118,31,26,31,85,31,71,31,71,30,170,31,202,31,76,31,76,30,159,31,153,31,35,31,226,31,213,31,36,31,80,31,80,30,125,31,19,31,27,31,27,30,24,31,224,31,170,31,170,30,183,31,39,31,130,31,188,31,237,31,223,31,127,31,127,30,100,31,16,31,107,31,6,31,120,31,34,31,34,30,170,31,170,30,170,29,170,28,96,31,144,31,185,31,152,31,159,31,154,31,30,31,210,31,103,31,103,30,32,31,242,31,55,31,242,31,231,31,118,31,246,31,246,30,44,31,145,31,120,31,120,30,188,31,13,31,13,30,13,29,162,31,86,31,97,31,97,30,85,31,198,31,198,30,198,29,175,31,110,31,110,30,203,31,203,30,249,31,249,31,237,31,237,30,30,31,30,30,30,29,202,31,222,31,184,31,184,30,136,31,136,30,136,29,93,31,107,31,46,31,33,31,33,30,170,31,170,30,217,31,239,31,239,30,239,29,239,28,108,31,231,31,2,31,244,31,244,30,221,31,121,31,44,31,103,31,247,31,193,31,193,30,203,31,211,31,209,31,235,31,249,31,58,31,78,31,20,31,28,31,176,31,156,31,244,31,244,30,83,31,103,31,103,30,208,31,150,31,60,31,18,31,139,31,139,30,25,31,226,31,66,31,112,31,48,31,48,30,230,31,240,31,189,31,189,30,50,31,50,30,254,31,121,31,121,30,107,31,166,31,163,31,90,31,180,31,19,31,227,31,88,31,218,31,159,31,240,31,30,31,66,31,66,30,99,31,107,31,32,31,167,31,150,31,243,31,179,31,170,31,29,31,74,31,74,30,175,31,178,31,178,30,205,31,148,31,148,30,160,31,160,30,140,31,223,31,223,30,53,31,57,31,154,31,154,30,70,31,141,31,78,31,135,31,31,31,31,30,92,31,197,31,223,31,236,31,236,30,146,31,146,30,146,29,248,31,20,31,183,31,183,30,87,31,200,31,19,31,23,31,215,31,104,31,183,31,129,31,228,31,132,31,206,31,206,30,225,31,64,31,64,30,110,31,102,31,12,31,12,30,194,31,194,30,194,29,27,31,47,31,97,31,203,31,162,31,214,31,2,31,146,31,8,31,93,31,255,31,105,31,90,31,90,30,168,31,167,31,155,31,124,31,186,31,44,31,45,31,19,31,148,31,163,31,11,31,176,31,182,31,114,31,40,31,40,30,85,31,199,31,199,30,161,31,48,31,186,31,109,31,42,31,108,31,130,31,46,31,249,31,249,30,249,29,210,31,77,31,77,30,77,29,211,31,155,31,155,30,115,31,115,30,236,31,117,31,210,31,67,31,132,31,47,31,78,31,195,31,121,31,87,31,87,30,169,31,107,31,115,31,209,31,162,31,53,31,111,31,86,31,250,31,63,31,34,31,26,31,45,31,209,31,108,31,87,31,10,31,121,31,145,31,242,31,242,30,242,29,181,31,118,31,131,31,120,31,254,31,254,30,16,31,71,31,186,31,244,31,64,31,240,31,28,31,219,31,121,31,146,31,124,31,185,31,31,31,108,31,123,31,91,31,240,31,119,31,106,31,7,31,147,31,26,31,26,30,124,31,26,31,91,31,66,31,66,30,71,31,255,31,200,31,200,30,255,31,138,31,98,31,212,31,25,31,159,31,9,31,64,31,247,31,167,31,8,31,51,31,162,31,75,31,153,31,153,30,102,31,165,31,123,31,130,31,214,31,190,31,102,31,102,30,91,31,91,30,91,29,205,31,19,31,163,31,66,31,167,31,16,31,150,31,141,31,101,31,101,30,101,29,101,28,95,31,109,31,179,31,26,31,202,31,144,31,29,31,132,31,121,31,94,31,94,30,246,31,102,31,102,30,102,29,110,31,42,31,133,31,34,31,219,31,177,31,74,31,126,31,129,31,129,30,129,29,129,28,129,27,129,26,13,31,63,31,99,31,105,31,97,31,221,31,192,31,124,31,110,31,149,31,37,31,81,31,81,30,157,31,130,31,130,30,130,29,130,28,87,31,87,30,87,29,145,31,195,31,125,31,42,31,162,31,162,30,162,29,110,31,110,30,87,31,25,31,130,31,200,31,110,31,110,30,110,29,174,31,174,30,174,29,174,28,245,31,75,31,75,30,69,31,197,31,174,31,174,30,110,31,167,31,93,31,60,31,94,31,23,31,94,31,212,31,240,31,215,31,215,30,140,31,140,30,140,29,190,31,223,31,223,30,223,29,61,31,215,31,215,30,175,31,190,31,194,31,90,31,28,31,45,31,110,31,110,30,107,31,130,31,139,31,212,31,186,31,194,31,82,31,121,31,121,30,139,31,24,31,83,31,28,31,88,31,88,30,164,31,222,31,224,31,224,30,247,31,155,31,155,30,163,31,1,31,192,31,126,31,109,31,1,31,9,31,167,31,31,31,186,31,216,31,231,31,224,31,153,31,200,31,186,31,186,30,86,31,62,31,37,31,37,30,212,31,212,30,207,31,114,31,18,31,18,30,18,29,6,31,136,31,136,30,118,31,136,31,136,30,136,29,143,31,143,30,94,31,59,31,73,31,102,31,102,30,87,31,87,30,171,31,171,30,171,29,199,31,171,31,44,31,254,31,47,31,114,31,59,31,59,30,68,31,68,30,33,31,55,31,55,30,48,31,215,31,120,31,47,31,13,31,13,30,133,31,150,31,199,31,86,31,244,31,211,31,93,31,151,31,93,31,37,31,114,31,173,31,45,31,45,30,29,31,184,31,184,30,68,31,82,31,171,31,104,31,190,31,190,30,170,31,164,31,243,31,251,31,36,31,82,31,56,31,56,30,9,31,38,31,137,31,137,30,165,31,165,30,176,31,173,31,158,31,64,31,64,30,53,31,119,31,71,31,168,31,30,31,131,31,59,31,191,31,224,31,103,31,255,31,169,31,149,31,107,31,199,31,97,31,14,31,210,31,114,31,150,31,143,31,143,30,187,31,200,31,70,31,76,31,76,30,23,31,224,31,178,31,191,31,191,30,122,31,167,31,167,30,13,31,97,31,212,31,212,30,109,31,69,31,213,31,247,31,71,31,71,30,219,31,35,31,35,30,27,31,166,31,16,31,16,30,77,31,184,31,244,31,42,31,124,31,124,30,40,31,128,31,180,31,19,31,61,31,33,31,216,31,216,30,128,31,128,30,141,31,26,31,191,31,201,31,158,31,85,31,98,31,11,31,127,31,127,30,203,31,234,31,217,31,109,31,109,30,106,31,111,31,111,30,15,31,7,31,239,31,6,31,164,31,173,31,182,31,182,30,84,31,38,31,38,30,38,29,127,31,127,30,72,31,72,30,29,31,83,31,129,31,101,31,204,31,204,30,135,31,176,31,34,31,34,30,218,31,218,30,25,31,16,31,166,31,166,30,107,31,107,30,38,31,38,30,106,31,106,30,106,29,143,31,35,31,177,31,206,31,206,30,40,31,40,30,40,29,154,31,8,31,15,31,98,31,57,31,93,31,186,31,127,31,190,31,190,30,190,29,174,31,249,31,132,31,132,30,132,29,170,31,8,31,214,31,214,30,214,29,22,31,22,30,212,31,212,30,13,31,77,31,77,30,110,31,195,31,145,31,145,30,4,31,94,31,51,31,47,31,47,30,164,31,31,31,254,31,254,30,160,31,103,31,36,31,36,30,22,31,218,31,163,31,125,31,115,31,106,31,30,31,203,31,49,31,255,31,19,31,169,31,61,31,57,31,163,31,115,31,97,31,121,31,46,31,141,31,38,31,38,30,223,31,11,31,11,30,190,31,133,31,133,30,133,29,220,31,50,31,95,31,246,31,29,31,29,30,230,31,230,30,153,31,32,31,32,30,92,31,153,31,153,30,249,31,114,31,114,30,145,31,100,31,100,30,2,31,162,31,162,30,162,29,225,31,139,31,202,31,42,31,231,31,231,30,180,31,178,31,24,31,253,31,242,31,102,31,47,31,20,31,156,31,178,31,219,31,219,30,127,31,127,30,127,29,127,28,102,31,10,31,212,31,174,31,174,30,174,29,237,31,199,31,9,31,9,30,248,31,10,31,10,30,133,31,181,31,122,31,177,31,56,31,11,31,93,31,132,31,252,31,252,30,155,31,60,31,69,31,193,31,226,31,23,31,52,31,52,30,247,31,247,30,137,31,2,31,72,31,72,30,14,31,119,31,25,31,25,30,139,31,118,31,166,31,166,30,19,31,124,31,174,31,103,31,22,31,100,31,100,30,72,31,213,31,103,31,111,31,75,31,149,31,46,31,66,31,50,31,112,31,34,31,107,31,221,31,200,31,80,31,25,31,25,30,80,31,109,31,152,31,171,31,116,31,116,30,200,31,147,31,7,31,51,31,153,31,153,30,153,29,153,28,153,27,189,31,1,31,1,30,172,31,189,31,140,31,103,31,150,31,5,31,31,31,108,31,100,31,49,31,215,31,215,30,215,29,244,31,203,31,155,31,200,31,201,31,201,30,119,31,235,31,222,31,222,30,183,31,183,30,31,31,237,31,8,31,8,30,146,31,194,31,63,31,221,31,141,31,73,31,36,31,30,31,109,31,109,30,222,31,126,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
