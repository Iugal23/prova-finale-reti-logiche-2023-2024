-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 371;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (52,0,48,0,147,0,206,0,167,0,59,0,122,0,125,0,130,0,79,0,213,0,28,0,189,0,68,0,107,0,122,0,111,0,18,0,0,0,51,0,130,0,227,0,81,0,156,0,245,0,135,0,0,0,47,0,0,0,18,0,31,0,151,0,47,0,0,0,166,0,92,0,30,0,147,0,0,0,37,0,208,0,0,0,0,0,163,0,0,0,0,0,216,0,248,0,0,0,146,0,0,0,7,0,223,0,194,0,156,0,138,0,143,0,162,0,19,0,118,0,251,0,217,0,47,0,0,0,194,0,171,0,157,0,202,0,41,0,28,0,0,0,0,0,153,0,176,0,14,0,181,0,241,0,58,0,92,0,72,0,114,0,64,0,254,0,178,0,183,0,116,0,45,0,254,0,113,0,220,0,239,0,28,0,0,0,91,0,223,0,147,0,0,0,190,0,131,0,133,0,193,0,251,0,225,0,238,0,180,0,134,0,94,0,182,0,226,0,0,0,0,0,15,0,0,0,175,0,117,0,199,0,43,0,110,0,0,0,75,0,202,0,236,0,126,0,52,0,52,0,139,0,0,0,33,0,97,0,28,0,70,0,91,0,219,0,0,0,203,0,0,0,50,0,0,0,28,0,78,0,138,0,35,0,71,0,116,0,182,0,142,0,99,0,87,0,26,0,162,0,192,0,0,0,254,0,23,0,77,0,0,0,0,0,87,0,0,0,133,0,32,0,50,0,22,0,0,0,204,0,95,0,0,0,223,0,0,0,28,0,253,0,222,0,151,0,4,0,27,0,119,0,28,0,207,0,76,0,0,0,166,0,9,0,194,0,234,0,0,0,0,0,0,0,71,0,0,0,87,0,0,0,135,0,78,0,0,0,245,0,206,0,217,0,229,0,0,0,238,0,9,0,0,0,248,0,0,0,230,0,245,0,223,0,158,0,154,0,184,0,0,0,0,0,161,0,5,0,0,0,43,0,58,0,77,0,45,0,7,0,129,0,200,0,196,0,162,0,98,0,101,0,196,0,144,0,235,0,242,0,144,0,55,0,93,0,136,0,0,0,161,0,201,0,246,0,10,0,144,0,99,0,124,0,0,0,199,0,79,0,65,0,101,0,0,0,191,0,0,0,213,0,226,0,0,0,97,0,40,0,101,0,87,0,206,0,107,0,152,0,7,0,0,0,205,0,0,0,17,0,142,0,8,0,0,0,220,0,40,0,198,0,145,0,148,0,155,0,202,0,0,0,74,0,82,0,0,0,218,0,244,0,12,0,58,0,147,0,86,0,95,0,253,0,93,0,155,0,68,0,238,0,141,0,78,0,142,0,243,0,59,0,186,0,113,0,139,0,160,0,0,0,183,0,49,0,155,0,95,0,0,0,200,0,186,0,36,0,21,0,18,0,241,0,67,0,155,0,74,0,0,0,64,0,0,0,86,0,110,0,119,0,234,0,26,0,105,0,88,0,157,0,206,0,127,0,222,0,215,0,0,0,40,0,0,0,125,0,0,0,30,0,0,0,53,0,254,0,223,0,47,0,60,0,0,0,0,0,0,0,103,0,155,0,135,0,5,0,0,0,247,0,86,0,203,0,160,0,80,0,134,0,140,0,171,0,192,0,209,0,0,0,220,0,69,0,94,0,176,0,0,0,210,0,29,0,123,0,213,0,78,0);
signal scenario_full  : scenario_type := (52,31,48,31,147,31,206,31,167,31,59,31,122,31,125,31,130,31,79,31,213,31,28,31,189,31,68,31,107,31,122,31,111,31,18,31,18,30,51,31,130,31,227,31,81,31,156,31,245,31,135,31,135,30,47,31,47,30,18,31,31,31,151,31,47,31,47,30,166,31,92,31,30,31,147,31,147,30,37,31,208,31,208,30,208,29,163,31,163,30,163,29,216,31,248,31,248,30,146,31,146,30,7,31,223,31,194,31,156,31,138,31,143,31,162,31,19,31,118,31,251,31,217,31,47,31,47,30,194,31,171,31,157,31,202,31,41,31,28,31,28,30,28,29,153,31,176,31,14,31,181,31,241,31,58,31,92,31,72,31,114,31,64,31,254,31,178,31,183,31,116,31,45,31,254,31,113,31,220,31,239,31,28,31,28,30,91,31,223,31,147,31,147,30,190,31,131,31,133,31,193,31,251,31,225,31,238,31,180,31,134,31,94,31,182,31,226,31,226,30,226,29,15,31,15,30,175,31,117,31,199,31,43,31,110,31,110,30,75,31,202,31,236,31,126,31,52,31,52,31,139,31,139,30,33,31,97,31,28,31,70,31,91,31,219,31,219,30,203,31,203,30,50,31,50,30,28,31,78,31,138,31,35,31,71,31,116,31,182,31,142,31,99,31,87,31,26,31,162,31,192,31,192,30,254,31,23,31,77,31,77,30,77,29,87,31,87,30,133,31,32,31,50,31,22,31,22,30,204,31,95,31,95,30,223,31,223,30,28,31,253,31,222,31,151,31,4,31,27,31,119,31,28,31,207,31,76,31,76,30,166,31,9,31,194,31,234,31,234,30,234,29,234,28,71,31,71,30,87,31,87,30,135,31,78,31,78,30,245,31,206,31,217,31,229,31,229,30,238,31,9,31,9,30,248,31,248,30,230,31,245,31,223,31,158,31,154,31,184,31,184,30,184,29,161,31,5,31,5,30,43,31,58,31,77,31,45,31,7,31,129,31,200,31,196,31,162,31,98,31,101,31,196,31,144,31,235,31,242,31,144,31,55,31,93,31,136,31,136,30,161,31,201,31,246,31,10,31,144,31,99,31,124,31,124,30,199,31,79,31,65,31,101,31,101,30,191,31,191,30,213,31,226,31,226,30,97,31,40,31,101,31,87,31,206,31,107,31,152,31,7,31,7,30,205,31,205,30,17,31,142,31,8,31,8,30,220,31,40,31,198,31,145,31,148,31,155,31,202,31,202,30,74,31,82,31,82,30,218,31,244,31,12,31,58,31,147,31,86,31,95,31,253,31,93,31,155,31,68,31,238,31,141,31,78,31,142,31,243,31,59,31,186,31,113,31,139,31,160,31,160,30,183,31,49,31,155,31,95,31,95,30,200,31,186,31,36,31,21,31,18,31,241,31,67,31,155,31,74,31,74,30,64,31,64,30,86,31,110,31,119,31,234,31,26,31,105,31,88,31,157,31,206,31,127,31,222,31,215,31,215,30,40,31,40,30,125,31,125,30,30,31,30,30,53,31,254,31,223,31,47,31,60,31,60,30,60,29,60,28,103,31,155,31,135,31,5,31,5,30,247,31,86,31,203,31,160,31,80,31,134,31,140,31,171,31,192,31,209,31,209,30,220,31,69,31,94,31,176,31,176,30,210,31,29,31,123,31,213,31,78,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
