-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_472 is
end project_tb_472;

architecture project_tb_arch_472 of project_tb_472 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 310;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,245,0,38,0,251,0,0,0,59,0,143,0,91,0,29,0,85,0,210,0,0,0,0,0,0,0,164,0,192,0,0,0,19,0,194,0,0,0,125,0,0,0,196,0,251,0,16,0,0,0,240,0,176,0,20,0,131,0,0,0,205,0,170,0,0,0,232,0,90,0,30,0,106,0,0,0,147,0,244,0,149,0,56,0,0,0,134,0,242,0,120,0,95,0,155,0,0,0,144,0,241,0,77,0,79,0,52,0,173,0,81,0,26,0,15,0,178,0,175,0,255,0,228,0,206,0,85,0,0,0,225,0,184,0,152,0,128,0,246,0,132,0,253,0,218,0,252,0,191,0,0,0,126,0,53,0,26,0,145,0,0,0,247,0,105,0,62,0,0,0,0,0,197,0,112,0,0,0,10,0,225,0,0,0,121,0,10,0,245,0,141,0,0,0,251,0,198,0,148,0,166,0,131,0,82,0,191,0,113,0,0,0,0,0,23,0,23,0,208,0,120,0,1,0,100,0,25,0,226,0,103,0,120,0,84,0,32,0,28,0,160,0,0,0,102,0,117,0,42,0,131,0,246,0,121,0,20,0,94,0,47,0,154,0,31,0,101,0,75,0,149,0,118,0,5,0,156,0,206,0,152,0,0,0,0,0,0,0,44,0,0,0,193,0,151,0,1,0,0,0,0,0,0,0,201,0,129,0,0,0,0,0,211,0,240,0,7,0,118,0,102,0,125,0,192,0,247,0,19,0,0,0,193,0,252,0,38,0,202,0,84,0,0,0,61,0,179,0,133,0,12,0,9,0,64,0,195,0,202,0,0,0,0,0,243,0,24,0,101,0,169,0,28,0,0,0,176,0,85,0,35,0,167,0,0,0,226,0,225,0,0,0,202,0,138,0,32,0,76,0,0,0,0,0,78,0,129,0,176,0,83,0,66,0,214,0,109,0,126,0,156,0,86,0,39,0,102,0,220,0,205,0,231,0,21,0,225,0,234,0,118,0,166,0,86,0,187,0,182,0,201,0,235,0,0,0,0,0,0,0,107,0,121,0,201,0,0,0,157,0,50,0,0,0,9,0,169,0,99,0,0,0,196,0,232,0,55,0,57,0,179,0,213,0,61,0,15,0,155,0,0,0,154,0,83,0,70,0,188,0,125,0,0,0,19,0,94,0,101,0,0,0,15,0,246,0,208,0,197,0,192,0,0,0,70,0,122,0,94,0,3,0,0,0,171,0,63,0,24,0,122,0,56,0,49,0,140,0,248,0,0,0,142,0,0,0,0,0,96,0,197,0,38,0,245,0,145,0,83,0,0,0,199,0,0,0,56,0,94,0,0,0,228,0,0,0,134,0,186,0,225,0,0,0,106,0,0,0,27,0,143,0,172,0,0,0,242,0);
signal scenario_full  : scenario_type := (0,0,245,31,38,31,251,31,251,30,59,31,143,31,91,31,29,31,85,31,210,31,210,30,210,29,210,28,164,31,192,31,192,30,19,31,194,31,194,30,125,31,125,30,196,31,251,31,16,31,16,30,240,31,176,31,20,31,131,31,131,30,205,31,170,31,170,30,232,31,90,31,30,31,106,31,106,30,147,31,244,31,149,31,56,31,56,30,134,31,242,31,120,31,95,31,155,31,155,30,144,31,241,31,77,31,79,31,52,31,173,31,81,31,26,31,15,31,178,31,175,31,255,31,228,31,206,31,85,31,85,30,225,31,184,31,152,31,128,31,246,31,132,31,253,31,218,31,252,31,191,31,191,30,126,31,53,31,26,31,145,31,145,30,247,31,105,31,62,31,62,30,62,29,197,31,112,31,112,30,10,31,225,31,225,30,121,31,10,31,245,31,141,31,141,30,251,31,198,31,148,31,166,31,131,31,82,31,191,31,113,31,113,30,113,29,23,31,23,31,208,31,120,31,1,31,100,31,25,31,226,31,103,31,120,31,84,31,32,31,28,31,160,31,160,30,102,31,117,31,42,31,131,31,246,31,121,31,20,31,94,31,47,31,154,31,31,31,101,31,75,31,149,31,118,31,5,31,156,31,206,31,152,31,152,30,152,29,152,28,44,31,44,30,193,31,151,31,1,31,1,30,1,29,1,28,201,31,129,31,129,30,129,29,211,31,240,31,7,31,118,31,102,31,125,31,192,31,247,31,19,31,19,30,193,31,252,31,38,31,202,31,84,31,84,30,61,31,179,31,133,31,12,31,9,31,64,31,195,31,202,31,202,30,202,29,243,31,24,31,101,31,169,31,28,31,28,30,176,31,85,31,35,31,167,31,167,30,226,31,225,31,225,30,202,31,138,31,32,31,76,31,76,30,76,29,78,31,129,31,176,31,83,31,66,31,214,31,109,31,126,31,156,31,86,31,39,31,102,31,220,31,205,31,231,31,21,31,225,31,234,31,118,31,166,31,86,31,187,31,182,31,201,31,235,31,235,30,235,29,235,28,107,31,121,31,201,31,201,30,157,31,50,31,50,30,9,31,169,31,99,31,99,30,196,31,232,31,55,31,57,31,179,31,213,31,61,31,15,31,155,31,155,30,154,31,83,31,70,31,188,31,125,31,125,30,19,31,94,31,101,31,101,30,15,31,246,31,208,31,197,31,192,31,192,30,70,31,122,31,94,31,3,31,3,30,171,31,63,31,24,31,122,31,56,31,49,31,140,31,248,31,248,30,142,31,142,30,142,29,96,31,197,31,38,31,245,31,145,31,83,31,83,30,199,31,199,30,56,31,94,31,94,30,228,31,228,30,134,31,186,31,225,31,225,30,106,31,106,30,27,31,143,31,172,31,172,30,242,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
