-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_281 is
end project_tb_281;

architecture project_tb_arch_281 of project_tb_281 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 987;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (232,0,185,0,0,0,125,0,65,0,0,0,81,0,0,0,73,0,172,0,44,0,182,0,105,0,0,0,53,0,88,0,230,0,189,0,0,0,82,0,18,0,78,0,68,0,118,0,159,0,50,0,124,0,154,0,118,0,96,0,187,0,119,0,0,0,0,0,0,0,0,0,127,0,63,0,188,0,4,0,247,0,242,0,117,0,7,0,228,0,33,0,216,0,33,0,177,0,201,0,152,0,53,0,0,0,59,0,129,0,174,0,0,0,198,0,226,0,0,0,0,0,141,0,0,0,240,0,91,0,203,0,0,0,13,0,149,0,0,0,0,0,0,0,195,0,145,0,176,0,0,0,12,0,231,0,175,0,140,0,0,0,20,0,112,0,51,0,239,0,208,0,166,0,154,0,0,0,118,0,0,0,193,0,247,0,14,0,227,0,66,0,222,0,236,0,48,0,0,0,178,0,68,0,10,0,127,0,107,0,84,0,211,0,169,0,63,0,90,0,11,0,0,0,132,0,0,0,147,0,34,0,0,0,141,0,195,0,250,0,73,0,24,0,171,0,198,0,51,0,91,0,0,0,200,0,102,0,0,0,29,0,0,0,12,0,189,0,139,0,0,0,166,0,47,0,219,0,0,0,96,0,197,0,64,0,58,0,159,0,0,0,100,0,105,0,97,0,157,0,0,0,253,0,26,0,160,0,184,0,0,0,56,0,178,0,0,0,125,0,226,0,43,0,66,0,238,0,0,0,47,0,167,0,73,0,223,0,0,0,6,0,87,0,218,0,176,0,30,0,145,0,68,0,215,0,203,0,100,0,18,0,0,0,42,0,33,0,25,0,149,0,90,0,191,0,0,0,171,0,81,0,23,0,196,0,201,0,139,0,169,0,49,0,161,0,0,0,57,0,93,0,69,0,11,0,56,0,189,0,0,0,84,0,161,0,69,0,0,0,101,0,185,0,90,0,193,0,2,0,79,0,29,0,0,0,0,0,0,0,238,0,44,0,71,0,112,0,180,0,226,0,48,0,101,0,142,0,177,0,86,0,0,0,14,0,241,0,213,0,133,0,29,0,50,0,0,0,51,0,123,0,245,0,20,0,80,0,121,0,117,0,31,0,203,0,108,0,175,0,115,0,115,0,52,0,232,0,13,0,95,0,0,0,13,0,59,0,66,0,25,0,36,0,0,0,186,0,47,0,116,0,0,0,189,0,232,0,246,0,228,0,238,0,202,0,108,0,197,0,241,0,20,0,0,0,151,0,0,0,8,0,144,0,124,0,114,0,206,0,179,0,77,0,15,0,0,0,243,0,203,0,158,0,168,0,215,0,234,0,126,0,71,0,0,0,201,0,156,0,9,0,70,0,51,0,0,0,239,0,229,0,166,0,0,0,143,0,196,0,0,0,0,0,199,0,98,0,181,0,199,0,238,0,160,0,73,0,9,0,65,0,88,0,0,0,75,0,177,0,0,0,0,0,18,0,27,0,0,0,59,0,0,0,145,0,0,0,173,0,153,0,195,0,209,0,72,0,245,0,0,0,80,0,136,0,0,0,73,0,174,0,0,0,1,0,160,0,68,0,60,0,0,0,71,0,127,0,93,0,0,0,118,0,237,0,184,0,16,0,108,0,68,0,150,0,3,0,176,0,0,0,223,0,209,0,0,0,51,0,205,0,95,0,112,0,175,0,63,0,19,0,127,0,0,0,0,0,143,0,254,0,183,0,8,0,9,0,0,0,128,0,0,0,112,0,181,0,82,0,40,0,157,0,203,0,196,0,121,0,211,0,35,0,108,0,150,0,149,0,0,0,0,0,0,0,60,0,28,0,136,0,187,0,153,0,227,0,234,0,108,0,0,0,222,0,8,0,0,0,233,0,193,0,0,0,226,0,235,0,0,0,0,0,0,0,160,0,28,0,0,0,103,0,227,0,34,0,174,0,228,0,183,0,144,0,246,0,3,0,155,0,252,0,0,0,152,0,0,0,0,0,49,0,2,0,91,0,34,0,81,0,189,0,31,0,134,0,0,0,1,0,201,0,59,0,199,0,0,0,183,0,38,0,0,0,147,0,192,0,50,0,64,0,242,0,186,0,15,0,167,0,99,0,40,0,170,0,0,0,172,0,126,0,189,0,0,0,159,0,166,0,0,0,180,0,0,0,55,0,149,0,0,0,90,0,0,0,105,0,254,0,175,0,5,0,216,0,107,0,149,0,178,0,175,0,0,0,46,0,171,0,16,0,193,0,119,0,0,0,57,0,82,0,165,0,65,0,0,0,218,0,19,0,84,0,122,0,119,0,62,0,0,0,0,0,0,0,217,0,235,0,223,0,89,0,148,0,0,0,144,0,0,0,222,0,159,0,174,0,101,0,157,0,63,0,243,0,0,0,81,0,211,0,137,0,0,0,0,0,152,0,0,0,12,0,176,0,34,0,122,0,0,0,8,0,216,0,0,0,0,0,1,0,0,0,252,0,177,0,146,0,10,0,0,0,194,0,180,0,247,0,0,0,30,0,195,0,14,0,231,0,221,0,31,0,228,0,77,0,0,0,87,0,168,0,27,0,227,0,42,0,60,0,223,0,0,0,240,0,19,0,0,0,0,0,86,0,0,0,108,0,209,0,0,0,252,0,0,0,20,0,202,0,48,0,94,0,22,0,219,0,37,0,0,0,81,0,0,0,114,0,0,0,142,0,47,0,19,0,241,0,133,0,24,0,185,0,237,0,0,0,86,0,254,0,5,0,0,0,3,0,14,0,46,0,0,0,218,0,127,0,102,0,200,0,14,0,37,0,221,0,80,0,173,0,182,0,0,0,177,0,227,0,87,0,156,0,168,0,75,0,91,0,23,0,153,0,123,0,17,0,77,0,0,0,21,0,0,0,64,0,128,0,146,0,7,0,155,0,0,0,26,0,158,0,14,0,119,0,18,0,145,0,50,0,0,0,17,0,0,0,61,0,0,0,55,0,0,0,99,0,72,0,177,0,118,0,0,0,0,0,47,0,0,0,0,0,2,0,21,0,227,0,79,0,0,0,70,0,51,0,0,0,58,0,29,0,81,0,84,0,35,0,139,0,140,0,143,0,119,0,161,0,111,0,252,0,172,0,136,0,0,0,0,0,150,0,147,0,123,0,62,0,131,0,85,0,31,0,36,0,0,0,97,0,187,0,0,0,106,0,216,0,254,0,69,0,233,0,6,0,158,0,137,0,179,0,253,0,147,0,0,0,143,0,0,0,220,0,60,0,62,0,237,0,147,0,33,0,0,0,211,0,197,0,40,0,29,0,122,0,134,0,36,0,121,0,147,0,45,0,99,0,196,0,0,0,104,0,186,0,86,0,203,0,0,0,8,0,154,0,56,0,5,0,63,0,166,0,31,0,235,0,152,0,8,0,221,0,150,0,58,0,212,0,0,0,186,0,69,0,212,0,0,0,234,0,0,0,0,0,94,0,0,0,19,0,197,0,127,0,111,0,215,0,89,0,34,0,0,0,148,0,1,0,4,0,0,0,152,0,232,0,206,0,0,0,0,0,90,0,205,0,254,0,0,0,154,0,99,0,178,0,214,0,0,0,94,0,85,0,197,0,0,0,0,0,113,0,0,0,143,0,251,0,140,0,116,0,144,0,249,0,0,0,0,0,138,0,100,0,219,0,128,0,162,0,165,0,80,0,164,0,133,0,177,0,219,0,78,0,15,0,0,0,24,0,0,0,0,0,38,0,41,0,35,0,240,0,217,0,235,0,133,0,57,0,250,0,71,0,218,0,0,0,222,0,0,0,0,0,70,0,162,0,150,0,225,0,109,0,0,0,173,0,205,0,134,0,203,0,117,0,0,0,0,0,0,0,42,0,114,0,21,0,128,0,81,0,14,0,0,0,119,0,0,0,0,0,115,0,69,0,104,0,0,0,29,0,91,0,0,0,0,0,0,0,231,0,109,0,68,0,197,0,0,0,0,0,247,0,40,0,109,0,247,0,212,0,0,0,41,0,232,0,124,0,172,0,0,0,41,0,135,0,66,0,140,0,120,0,0,0,149,0,0,0,105,0,0,0,0,0,27,0,11,0,171,0,167,0,160,0,86,0,58,0,203,0,130,0,0,0,46,0,97,0,0,0,42,0,191,0,8,0,0,0,46,0,0,0,200,0,189,0,159,0,0,0,178,0,34,0,0,0,137,0,0,0,38,0,0,0,240,0,181,0,150,0,80,0,252,0,71,0,160,0,61,0,204,0,16,0,246,0,0,0,228,0,203,0,53,0,20,0,83,0,24,0,0,0,134,0,0,0,204,0,185,0,120,0,249,0,85,0,133,0,25,0,199,0,205,0,0,0,144,0,0,0,0,0,254,0,254,0,50,0,0,0,55,0,19,0,92,0,73,0,156,0,212,0,90,0,164,0,210,0,0,0,0,0,93,0,143,0,244,0,2,0,0,0,128,0);
signal scenario_full  : scenario_type := (232,31,185,31,185,30,125,31,65,31,65,30,81,31,81,30,73,31,172,31,44,31,182,31,105,31,105,30,53,31,88,31,230,31,189,31,189,30,82,31,18,31,78,31,68,31,118,31,159,31,50,31,124,31,154,31,118,31,96,31,187,31,119,31,119,30,119,29,119,28,119,27,127,31,63,31,188,31,4,31,247,31,242,31,117,31,7,31,228,31,33,31,216,31,33,31,177,31,201,31,152,31,53,31,53,30,59,31,129,31,174,31,174,30,198,31,226,31,226,30,226,29,141,31,141,30,240,31,91,31,203,31,203,30,13,31,149,31,149,30,149,29,149,28,195,31,145,31,176,31,176,30,12,31,231,31,175,31,140,31,140,30,20,31,112,31,51,31,239,31,208,31,166,31,154,31,154,30,118,31,118,30,193,31,247,31,14,31,227,31,66,31,222,31,236,31,48,31,48,30,178,31,68,31,10,31,127,31,107,31,84,31,211,31,169,31,63,31,90,31,11,31,11,30,132,31,132,30,147,31,34,31,34,30,141,31,195,31,250,31,73,31,24,31,171,31,198,31,51,31,91,31,91,30,200,31,102,31,102,30,29,31,29,30,12,31,189,31,139,31,139,30,166,31,47,31,219,31,219,30,96,31,197,31,64,31,58,31,159,31,159,30,100,31,105,31,97,31,157,31,157,30,253,31,26,31,160,31,184,31,184,30,56,31,178,31,178,30,125,31,226,31,43,31,66,31,238,31,238,30,47,31,167,31,73,31,223,31,223,30,6,31,87,31,218,31,176,31,30,31,145,31,68,31,215,31,203,31,100,31,18,31,18,30,42,31,33,31,25,31,149,31,90,31,191,31,191,30,171,31,81,31,23,31,196,31,201,31,139,31,169,31,49,31,161,31,161,30,57,31,93,31,69,31,11,31,56,31,189,31,189,30,84,31,161,31,69,31,69,30,101,31,185,31,90,31,193,31,2,31,79,31,29,31,29,30,29,29,29,28,238,31,44,31,71,31,112,31,180,31,226,31,48,31,101,31,142,31,177,31,86,31,86,30,14,31,241,31,213,31,133,31,29,31,50,31,50,30,51,31,123,31,245,31,20,31,80,31,121,31,117,31,31,31,203,31,108,31,175,31,115,31,115,31,52,31,232,31,13,31,95,31,95,30,13,31,59,31,66,31,25,31,36,31,36,30,186,31,47,31,116,31,116,30,189,31,232,31,246,31,228,31,238,31,202,31,108,31,197,31,241,31,20,31,20,30,151,31,151,30,8,31,144,31,124,31,114,31,206,31,179,31,77,31,15,31,15,30,243,31,203,31,158,31,168,31,215,31,234,31,126,31,71,31,71,30,201,31,156,31,9,31,70,31,51,31,51,30,239,31,229,31,166,31,166,30,143,31,196,31,196,30,196,29,199,31,98,31,181,31,199,31,238,31,160,31,73,31,9,31,65,31,88,31,88,30,75,31,177,31,177,30,177,29,18,31,27,31,27,30,59,31,59,30,145,31,145,30,173,31,153,31,195,31,209,31,72,31,245,31,245,30,80,31,136,31,136,30,73,31,174,31,174,30,1,31,160,31,68,31,60,31,60,30,71,31,127,31,93,31,93,30,118,31,237,31,184,31,16,31,108,31,68,31,150,31,3,31,176,31,176,30,223,31,209,31,209,30,51,31,205,31,95,31,112,31,175,31,63,31,19,31,127,31,127,30,127,29,143,31,254,31,183,31,8,31,9,31,9,30,128,31,128,30,112,31,181,31,82,31,40,31,157,31,203,31,196,31,121,31,211,31,35,31,108,31,150,31,149,31,149,30,149,29,149,28,60,31,28,31,136,31,187,31,153,31,227,31,234,31,108,31,108,30,222,31,8,31,8,30,233,31,193,31,193,30,226,31,235,31,235,30,235,29,235,28,160,31,28,31,28,30,103,31,227,31,34,31,174,31,228,31,183,31,144,31,246,31,3,31,155,31,252,31,252,30,152,31,152,30,152,29,49,31,2,31,91,31,34,31,81,31,189,31,31,31,134,31,134,30,1,31,201,31,59,31,199,31,199,30,183,31,38,31,38,30,147,31,192,31,50,31,64,31,242,31,186,31,15,31,167,31,99,31,40,31,170,31,170,30,172,31,126,31,189,31,189,30,159,31,166,31,166,30,180,31,180,30,55,31,149,31,149,30,90,31,90,30,105,31,254,31,175,31,5,31,216,31,107,31,149,31,178,31,175,31,175,30,46,31,171,31,16,31,193,31,119,31,119,30,57,31,82,31,165,31,65,31,65,30,218,31,19,31,84,31,122,31,119,31,62,31,62,30,62,29,62,28,217,31,235,31,223,31,89,31,148,31,148,30,144,31,144,30,222,31,159,31,174,31,101,31,157,31,63,31,243,31,243,30,81,31,211,31,137,31,137,30,137,29,152,31,152,30,12,31,176,31,34,31,122,31,122,30,8,31,216,31,216,30,216,29,1,31,1,30,252,31,177,31,146,31,10,31,10,30,194,31,180,31,247,31,247,30,30,31,195,31,14,31,231,31,221,31,31,31,228,31,77,31,77,30,87,31,168,31,27,31,227,31,42,31,60,31,223,31,223,30,240,31,19,31,19,30,19,29,86,31,86,30,108,31,209,31,209,30,252,31,252,30,20,31,202,31,48,31,94,31,22,31,219,31,37,31,37,30,81,31,81,30,114,31,114,30,142,31,47,31,19,31,241,31,133,31,24,31,185,31,237,31,237,30,86,31,254,31,5,31,5,30,3,31,14,31,46,31,46,30,218,31,127,31,102,31,200,31,14,31,37,31,221,31,80,31,173,31,182,31,182,30,177,31,227,31,87,31,156,31,168,31,75,31,91,31,23,31,153,31,123,31,17,31,77,31,77,30,21,31,21,30,64,31,128,31,146,31,7,31,155,31,155,30,26,31,158,31,14,31,119,31,18,31,145,31,50,31,50,30,17,31,17,30,61,31,61,30,55,31,55,30,99,31,72,31,177,31,118,31,118,30,118,29,47,31,47,30,47,29,2,31,21,31,227,31,79,31,79,30,70,31,51,31,51,30,58,31,29,31,81,31,84,31,35,31,139,31,140,31,143,31,119,31,161,31,111,31,252,31,172,31,136,31,136,30,136,29,150,31,147,31,123,31,62,31,131,31,85,31,31,31,36,31,36,30,97,31,187,31,187,30,106,31,216,31,254,31,69,31,233,31,6,31,158,31,137,31,179,31,253,31,147,31,147,30,143,31,143,30,220,31,60,31,62,31,237,31,147,31,33,31,33,30,211,31,197,31,40,31,29,31,122,31,134,31,36,31,121,31,147,31,45,31,99,31,196,31,196,30,104,31,186,31,86,31,203,31,203,30,8,31,154,31,56,31,5,31,63,31,166,31,31,31,235,31,152,31,8,31,221,31,150,31,58,31,212,31,212,30,186,31,69,31,212,31,212,30,234,31,234,30,234,29,94,31,94,30,19,31,197,31,127,31,111,31,215,31,89,31,34,31,34,30,148,31,1,31,4,31,4,30,152,31,232,31,206,31,206,30,206,29,90,31,205,31,254,31,254,30,154,31,99,31,178,31,214,31,214,30,94,31,85,31,197,31,197,30,197,29,113,31,113,30,143,31,251,31,140,31,116,31,144,31,249,31,249,30,249,29,138,31,100,31,219,31,128,31,162,31,165,31,80,31,164,31,133,31,177,31,219,31,78,31,15,31,15,30,24,31,24,30,24,29,38,31,41,31,35,31,240,31,217,31,235,31,133,31,57,31,250,31,71,31,218,31,218,30,222,31,222,30,222,29,70,31,162,31,150,31,225,31,109,31,109,30,173,31,205,31,134,31,203,31,117,31,117,30,117,29,117,28,42,31,114,31,21,31,128,31,81,31,14,31,14,30,119,31,119,30,119,29,115,31,69,31,104,31,104,30,29,31,91,31,91,30,91,29,91,28,231,31,109,31,68,31,197,31,197,30,197,29,247,31,40,31,109,31,247,31,212,31,212,30,41,31,232,31,124,31,172,31,172,30,41,31,135,31,66,31,140,31,120,31,120,30,149,31,149,30,105,31,105,30,105,29,27,31,11,31,171,31,167,31,160,31,86,31,58,31,203,31,130,31,130,30,46,31,97,31,97,30,42,31,191,31,8,31,8,30,46,31,46,30,200,31,189,31,159,31,159,30,178,31,34,31,34,30,137,31,137,30,38,31,38,30,240,31,181,31,150,31,80,31,252,31,71,31,160,31,61,31,204,31,16,31,246,31,246,30,228,31,203,31,53,31,20,31,83,31,24,31,24,30,134,31,134,30,204,31,185,31,120,31,249,31,85,31,133,31,25,31,199,31,205,31,205,30,144,31,144,30,144,29,254,31,254,31,50,31,50,30,55,31,19,31,92,31,73,31,156,31,212,31,90,31,164,31,210,31,210,30,210,29,93,31,143,31,244,31,2,31,2,30,128,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
