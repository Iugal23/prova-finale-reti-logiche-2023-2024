-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_298 is
end project_tb_298;

architecture project_tb_arch_298 of project_tb_298 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 232;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (250,0,98,0,100,0,0,0,98,0,64,0,0,0,0,0,164,0,19,0,96,0,194,0,6,0,0,0,57,0,68,0,70,0,18,0,227,0,62,0,121,0,214,0,0,0,0,0,135,0,0,0,0,0,149,0,153,0,98,0,181,0,21,0,0,0,54,0,36,0,170,0,202,0,191,0,46,0,183,0,74,0,217,0,0,0,246,0,70,0,46,0,51,0,11,0,120,0,30,0,0,0,215,0,0,0,149,0,107,0,0,0,39,0,149,0,0,0,16,0,253,0,201,0,206,0,198,0,255,0,20,0,64,0,190,0,153,0,220,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,165,0,0,0,106,0,217,0,37,0,241,0,4,0,0,0,0,0,0,0,173,0,0,0,47,0,0,0,73,0,10,0,71,0,8,0,233,0,148,0,150,0,223,0,47,0,106,0,53,0,141,0,214,0,134,0,185,0,96,0,214,0,232,0,237,0,40,0,233,0,0,0,102,0,239,0,37,0,0,0,190,0,66,0,188,0,0,0,101,0,0,0,18,0,62,0,0,0,46,0,110,0,86,0,177,0,39,0,250,0,211,0,17,0,4,0,68,0,104,0,93,0,0,0,218,0,37,0,224,0,251,0,155,0,118,0,72,0,0,0,29,0,138,0,173,0,231,0,185,0,186,0,105,0,98,0,39,0,244,0,118,0,129,0,20,0,0,0,191,0,69,0,82,0,244,0,0,0,181,0,157,0,226,0,66,0,212,0,111,0,108,0,116,0,190,0,225,0,185,0,174,0,154,0,219,0,190,0,167,0,165,0,202,0,16,0,160,0,7,0,4,0,237,0,136,0,150,0,48,0,7,0,23,0,118,0,0,0,49,0,43,0,111,0,128,0,207,0,218,0,77,0,196,0,0,0,85,0,203,0,144,0,131,0,66,0,0,0,0,0,221,0,55,0,246,0,113,0,0,0,0,0,27,0,64,0,212,0,248,0,0,0,121,0,192,0,0,0,39,0,164,0,17,0,197,0,123,0,42,0);
signal scenario_full  : scenario_type := (250,31,98,31,100,31,100,30,98,31,64,31,64,30,64,29,164,31,19,31,96,31,194,31,6,31,6,30,57,31,68,31,70,31,18,31,227,31,62,31,121,31,214,31,214,30,214,29,135,31,135,30,135,29,149,31,153,31,98,31,181,31,21,31,21,30,54,31,36,31,170,31,202,31,191,31,46,31,183,31,74,31,217,31,217,30,246,31,70,31,46,31,51,31,11,31,120,31,30,31,30,30,215,31,215,30,149,31,107,31,107,30,39,31,149,31,149,30,16,31,253,31,201,31,206,31,198,31,255,31,20,31,64,31,190,31,153,31,220,31,220,30,220,29,220,28,220,27,220,26,220,25,220,24,165,31,165,30,106,31,217,31,37,31,241,31,4,31,4,30,4,29,4,28,173,31,173,30,47,31,47,30,73,31,10,31,71,31,8,31,233,31,148,31,150,31,223,31,47,31,106,31,53,31,141,31,214,31,134,31,185,31,96,31,214,31,232,31,237,31,40,31,233,31,233,30,102,31,239,31,37,31,37,30,190,31,66,31,188,31,188,30,101,31,101,30,18,31,62,31,62,30,46,31,110,31,86,31,177,31,39,31,250,31,211,31,17,31,4,31,68,31,104,31,93,31,93,30,218,31,37,31,224,31,251,31,155,31,118,31,72,31,72,30,29,31,138,31,173,31,231,31,185,31,186,31,105,31,98,31,39,31,244,31,118,31,129,31,20,31,20,30,191,31,69,31,82,31,244,31,244,30,181,31,157,31,226,31,66,31,212,31,111,31,108,31,116,31,190,31,225,31,185,31,174,31,154,31,219,31,190,31,167,31,165,31,202,31,16,31,160,31,7,31,4,31,237,31,136,31,150,31,48,31,7,31,23,31,118,31,118,30,49,31,43,31,111,31,128,31,207,31,218,31,77,31,196,31,196,30,85,31,203,31,144,31,131,31,66,31,66,30,66,29,221,31,55,31,246,31,113,31,113,30,113,29,27,31,64,31,212,31,248,31,248,30,121,31,192,31,192,30,39,31,164,31,17,31,197,31,123,31,42,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
