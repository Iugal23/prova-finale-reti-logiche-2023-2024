-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_139 is
end project_tb_139;

architecture project_tb_arch_139 of project_tb_139 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 930;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (87,0,0,0,124,0,254,0,0,0,238,0,155,0,129,0,66,0,0,0,112,0,107,0,128,0,3,0,93,0,0,0,0,0,86,0,13,0,0,0,131,0,41,0,188,0,143,0,0,0,208,0,55,0,167,0,148,0,46,0,230,0,1,0,207,0,0,0,137,0,0,0,65,0,43,0,116,0,242,0,62,0,141,0,213,0,45,0,248,0,170,0,46,0,250,0,172,0,69,0,0,0,40,0,127,0,0,0,231,0,6,0,166,0,163,0,68,0,174,0,85,0,0,0,166,0,0,0,173,0,128,0,249,0,140,0,204,0,185,0,175,0,201,0,185,0,0,0,0,0,153,0,239,0,182,0,38,0,219,0,148,0,0,0,44,0,20,0,183,0,183,0,57,0,45,0,0,0,0,0,125,0,81,0,207,0,140,0,197,0,241,0,6,0,164,0,166,0,149,0,164,0,199,0,127,0,74,0,0,0,0,0,0,0,72,0,199,0,130,0,31,0,0,0,26,0,0,0,213,0,5,0,86,0,148,0,0,0,0,0,0,0,155,0,0,0,151,0,255,0,226,0,57,0,92,0,171,0,225,0,167,0,58,0,55,0,114,0,0,0,0,0,19,0,0,0,255,0,7,0,0,0,231,0,2,0,35,0,192,0,78,0,181,0,67,0,73,0,203,0,138,0,119,0,0,0,180,0,0,0,0,0,101,0,9,0,0,0,0,0,110,0,25,0,168,0,171,0,214,0,0,0,0,0,0,0,246,0,20,0,252,0,81,0,95,0,197,0,20,0,78,0,0,0,239,0,115,0,0,0,106,0,93,0,225,0,0,0,196,0,164,0,26,0,51,0,122,0,251,0,83,0,218,0,0,0,23,0,49,0,178,0,107,0,14,0,0,0,229,0,179,0,155,0,0,0,31,0,111,0,80,0,183,0,0,0,3,0,188,0,194,0,53,0,12,0,170,0,85,0,76,0,162,0,0,0,144,0,93,0,191,0,209,0,52,0,0,0,228,0,185,0,98,0,57,0,190,0,227,0,56,0,198,0,60,0,0,0,175,0,174,0,87,0,19,0,82,0,182,0,180,0,207,0,94,0,178,0,148,0,59,0,101,0,196,0,206,0,161,0,199,0,0,0,169,0,185,0,98,0,64,0,10,0,182,0,13,0,160,0,181,0,75,0,0,0,99,0,169,0,83,0,141,0,0,0,164,0,11,0,202,0,185,0,0,0,178,0,62,0,255,0,0,0,0,0,173,0,81,0,0,0,0,0,0,0,72,0,193,0,82,0,199,0,42,0,0,0,136,0,126,0,39,0,203,0,129,0,69,0,0,0,116,0,150,0,238,0,87,0,16,0,0,0,158,0,70,0,113,0,1,0,0,0,155,0,71,0,234,0,70,0,51,0,0,0,133,0,62,0,191,0,0,0,158,0,161,0,219,0,39,0,68,0,250,0,238,0,25,0,12,0,0,0,0,0,243,0,9,0,65,0,84,0,10,0,72,0,213,0,44,0,252,0,90,0,142,0,90,0,125,0,42,0,164,0,153,0,193,0,75,0,206,0,175,0,0,0,111,0,0,0,177,0,125,0,240,0,94,0,232,0,18,0,105,0,21,0,9,0,0,0,79,0,12,0,30,0,0,0,206,0,178,0,0,0,103,0,214,0,209,0,185,0,0,0,21,0,16,0,164,0,37,0,57,0,225,0,0,0,59,0,198,0,98,0,109,0,118,0,39,0,0,0,105,0,191,0,0,0,247,0,118,0,17,0,84,0,0,0,228,0,21,0,226,0,79,0,0,0,0,0,231,0,127,0,0,0,206,0,0,0,0,0,0,0,84,0,173,0,110,0,112,0,80,0,104,0,233,0,182,0,183,0,247,0,220,0,0,0,161,0,234,0,42,0,56,0,103,0,0,0,141,0,212,0,139,0,141,0,0,0,131,0,0,0,0,0,176,0,0,0,144,0,0,0,0,0,170,0,138,0,0,0,208,0,0,0,0,0,218,0,0,0,189,0,36,0,0,0,0,0,95,0,3,0,87,0,0,0,75,0,0,0,28,0,121,0,204,0,182,0,0,0,187,0,0,0,151,0,116,0,192,0,101,0,160,0,0,0,194,0,21,0,164,0,1,0,94,0,255,0,32,0,60,0,15,0,194,0,0,0,213,0,73,0,204,0,38,0,0,0,143,0,229,0,152,0,251,0,209,0,194,0,0,0,84,0,244,0,229,0,8,0,0,0,221,0,97,0,237,0,186,0,0,0,109,0,55,0,235,0,254,0,56,0,0,0,232,0,0,0,125,0,40,0,178,0,18,0,189,0,162,0,0,0,33,0,198,0,217,0,207,0,0,0,59,0,27,0,248,0,19,0,105,0,96,0,195,0,0,0,107,0,132,0,174,0,119,0,163,0,6,0,224,0,202,0,0,0,47,0,0,0,31,0,27,0,0,0,151,0,212,0,9,0,30,0,14,0,9,0,167,0,80,0,196,0,192,0,208,0,198,0,66,0,138,0,51,0,210,0,28,0,110,0,131,0,125,0,182,0,114,0,116,0,0,0,42,0,10,0,27,0,237,0,46,0,0,0,111,0,26,0,254,0,197,0,0,0,0,0,156,0,237,0,39,0,0,0,140,0,212,0,246,0,86,0,144,0,6,0,172,0,91,0,130,0,0,0,0,0,115,0,42,0,30,0,0,0,27,0,232,0,4,0,0,0,127,0,121,0,240,0,19,0,0,0,34,0,137,0,130,0,196,0,0,0,0,0,247,0,0,0,92,0,126,0,124,0,145,0,5,0,0,0,114,0,22,0,164,0,129,0,95,0,0,0,146,0,170,0,97,0,229,0,86,0,8,0,31,0,81,0,164,0,52,0,222,0,172,0,212,0,109,0,210,0,0,0,0,0,189,0,250,0,124,0,46,0,199,0,190,0,148,0,162,0,133,0,0,0,102,0,58,0,2,0,0,0,84,0,17,0,114,0,239,0,0,0,58,0,225,0,214,0,165,0,212,0,121,0,5,0,56,0,213,0,164,0,239,0,3,0,139,0,4,0,223,0,152,0,205,0,79,0,0,0,155,0,0,0,107,0,124,0,41,0,0,0,106,0,123,0,186,0,158,0,152,0,129,0,0,0,180,0,132,0,233,0,0,0,149,0,0,0,25,0,176,0,108,0,0,0,235,0,47,0,42,0,98,0,243,0,162,0,0,0,125,0,222,0,0,0,130,0,0,0,185,0,237,0,171,0,229,0,238,0,159,0,161,0,16,0,242,0,22,0,0,0,249,0,138,0,0,0,55,0,0,0,178,0,107,0,154,0,10,0,0,0,33,0,135,0,82,0,204,0,0,0,199,0,103,0,202,0,0,0,126,0,106,0,124,0,1,0,160,0,44,0,0,0,200,0,209,0,0,0,149,0,231,0,0,0,100,0,188,0,235,0,112,0,142,0,99,0,242,0,213,0,47,0,200,0,119,0,0,0,115,0,12,0,98,0,69,0,236,0,1,0,124,0,115,0,0,0,122,0,90,0,249,0,13,0,0,0,0,0,0,0,174,0,60,0,221,0,12,0,51,0,150,0,180,0,186,0,204,0,0,0,200,0,115,0,41,0,99,0,63,0,0,0,156,0,213,0,231,0,0,0,178,0,238,0,191,0,12,0,152,0,230,0,114,0,0,0,64,0,248,0,233,0,0,0,98,0,130,0,29,0,0,0,215,0,120,0,0,0,131,0,0,0,82,0,65,0,63,0,124,0,181,0,245,0,193,0,41,0,134,0,217,0,106,0,21,0,37,0,0,0,8,0,220,0,88,0,0,0,145,0,45,0,234,0,0,0,70,0,51,0,200,0,99,0,24,0,61,0,0,0,13,0,214,0,0,0,184,0,0,0,201,0,164,0,246,0,51,0,190,0,205,0,110,0,45,0,52,0,177,0,42,0,120,0,60,0,164,0,252,0,253,0,192,0,86,0,66,0,0,0,56,0,6,0,211,0,0,0,213,0,139,0,0,0,28,0,115,0,105,0,191,0,201,0,34,0,0,0,0,0,42,0,83,0,0,0,125,0,145,0,61,0,150,0,42,0,102,0,227,0,113,0,0,0,0,0,135,0,119,0,189,0,0,0,139,0,137,0,0,0,143,0,161,0,28,0,218,0,189,0,139,0,0,0,53,0,0,0,136,0);
signal scenario_full  : scenario_type := (87,31,87,30,124,31,254,31,254,30,238,31,155,31,129,31,66,31,66,30,112,31,107,31,128,31,3,31,93,31,93,30,93,29,86,31,13,31,13,30,131,31,41,31,188,31,143,31,143,30,208,31,55,31,167,31,148,31,46,31,230,31,1,31,207,31,207,30,137,31,137,30,65,31,43,31,116,31,242,31,62,31,141,31,213,31,45,31,248,31,170,31,46,31,250,31,172,31,69,31,69,30,40,31,127,31,127,30,231,31,6,31,166,31,163,31,68,31,174,31,85,31,85,30,166,31,166,30,173,31,128,31,249,31,140,31,204,31,185,31,175,31,201,31,185,31,185,30,185,29,153,31,239,31,182,31,38,31,219,31,148,31,148,30,44,31,20,31,183,31,183,31,57,31,45,31,45,30,45,29,125,31,81,31,207,31,140,31,197,31,241,31,6,31,164,31,166,31,149,31,164,31,199,31,127,31,74,31,74,30,74,29,74,28,72,31,199,31,130,31,31,31,31,30,26,31,26,30,213,31,5,31,86,31,148,31,148,30,148,29,148,28,155,31,155,30,151,31,255,31,226,31,57,31,92,31,171,31,225,31,167,31,58,31,55,31,114,31,114,30,114,29,19,31,19,30,255,31,7,31,7,30,231,31,2,31,35,31,192,31,78,31,181,31,67,31,73,31,203,31,138,31,119,31,119,30,180,31,180,30,180,29,101,31,9,31,9,30,9,29,110,31,25,31,168,31,171,31,214,31,214,30,214,29,214,28,246,31,20,31,252,31,81,31,95,31,197,31,20,31,78,31,78,30,239,31,115,31,115,30,106,31,93,31,225,31,225,30,196,31,164,31,26,31,51,31,122,31,251,31,83,31,218,31,218,30,23,31,49,31,178,31,107,31,14,31,14,30,229,31,179,31,155,31,155,30,31,31,111,31,80,31,183,31,183,30,3,31,188,31,194,31,53,31,12,31,170,31,85,31,76,31,162,31,162,30,144,31,93,31,191,31,209,31,52,31,52,30,228,31,185,31,98,31,57,31,190,31,227,31,56,31,198,31,60,31,60,30,175,31,174,31,87,31,19,31,82,31,182,31,180,31,207,31,94,31,178,31,148,31,59,31,101,31,196,31,206,31,161,31,199,31,199,30,169,31,185,31,98,31,64,31,10,31,182,31,13,31,160,31,181,31,75,31,75,30,99,31,169,31,83,31,141,31,141,30,164,31,11,31,202,31,185,31,185,30,178,31,62,31,255,31,255,30,255,29,173,31,81,31,81,30,81,29,81,28,72,31,193,31,82,31,199,31,42,31,42,30,136,31,126,31,39,31,203,31,129,31,69,31,69,30,116,31,150,31,238,31,87,31,16,31,16,30,158,31,70,31,113,31,1,31,1,30,155,31,71,31,234,31,70,31,51,31,51,30,133,31,62,31,191,31,191,30,158,31,161,31,219,31,39,31,68,31,250,31,238,31,25,31,12,31,12,30,12,29,243,31,9,31,65,31,84,31,10,31,72,31,213,31,44,31,252,31,90,31,142,31,90,31,125,31,42,31,164,31,153,31,193,31,75,31,206,31,175,31,175,30,111,31,111,30,177,31,125,31,240,31,94,31,232,31,18,31,105,31,21,31,9,31,9,30,79,31,12,31,30,31,30,30,206,31,178,31,178,30,103,31,214,31,209,31,185,31,185,30,21,31,16,31,164,31,37,31,57,31,225,31,225,30,59,31,198,31,98,31,109,31,118,31,39,31,39,30,105,31,191,31,191,30,247,31,118,31,17,31,84,31,84,30,228,31,21,31,226,31,79,31,79,30,79,29,231,31,127,31,127,30,206,31,206,30,206,29,206,28,84,31,173,31,110,31,112,31,80,31,104,31,233,31,182,31,183,31,247,31,220,31,220,30,161,31,234,31,42,31,56,31,103,31,103,30,141,31,212,31,139,31,141,31,141,30,131,31,131,30,131,29,176,31,176,30,144,31,144,30,144,29,170,31,138,31,138,30,208,31,208,30,208,29,218,31,218,30,189,31,36,31,36,30,36,29,95,31,3,31,87,31,87,30,75,31,75,30,28,31,121,31,204,31,182,31,182,30,187,31,187,30,151,31,116,31,192,31,101,31,160,31,160,30,194,31,21,31,164,31,1,31,94,31,255,31,32,31,60,31,15,31,194,31,194,30,213,31,73,31,204,31,38,31,38,30,143,31,229,31,152,31,251,31,209,31,194,31,194,30,84,31,244,31,229,31,8,31,8,30,221,31,97,31,237,31,186,31,186,30,109,31,55,31,235,31,254,31,56,31,56,30,232,31,232,30,125,31,40,31,178,31,18,31,189,31,162,31,162,30,33,31,198,31,217,31,207,31,207,30,59,31,27,31,248,31,19,31,105,31,96,31,195,31,195,30,107,31,132,31,174,31,119,31,163,31,6,31,224,31,202,31,202,30,47,31,47,30,31,31,27,31,27,30,151,31,212,31,9,31,30,31,14,31,9,31,167,31,80,31,196,31,192,31,208,31,198,31,66,31,138,31,51,31,210,31,28,31,110,31,131,31,125,31,182,31,114,31,116,31,116,30,42,31,10,31,27,31,237,31,46,31,46,30,111,31,26,31,254,31,197,31,197,30,197,29,156,31,237,31,39,31,39,30,140,31,212,31,246,31,86,31,144,31,6,31,172,31,91,31,130,31,130,30,130,29,115,31,42,31,30,31,30,30,27,31,232,31,4,31,4,30,127,31,121,31,240,31,19,31,19,30,34,31,137,31,130,31,196,31,196,30,196,29,247,31,247,30,92,31,126,31,124,31,145,31,5,31,5,30,114,31,22,31,164,31,129,31,95,31,95,30,146,31,170,31,97,31,229,31,86,31,8,31,31,31,81,31,164,31,52,31,222,31,172,31,212,31,109,31,210,31,210,30,210,29,189,31,250,31,124,31,46,31,199,31,190,31,148,31,162,31,133,31,133,30,102,31,58,31,2,31,2,30,84,31,17,31,114,31,239,31,239,30,58,31,225,31,214,31,165,31,212,31,121,31,5,31,56,31,213,31,164,31,239,31,3,31,139,31,4,31,223,31,152,31,205,31,79,31,79,30,155,31,155,30,107,31,124,31,41,31,41,30,106,31,123,31,186,31,158,31,152,31,129,31,129,30,180,31,132,31,233,31,233,30,149,31,149,30,25,31,176,31,108,31,108,30,235,31,47,31,42,31,98,31,243,31,162,31,162,30,125,31,222,31,222,30,130,31,130,30,185,31,237,31,171,31,229,31,238,31,159,31,161,31,16,31,242,31,22,31,22,30,249,31,138,31,138,30,55,31,55,30,178,31,107,31,154,31,10,31,10,30,33,31,135,31,82,31,204,31,204,30,199,31,103,31,202,31,202,30,126,31,106,31,124,31,1,31,160,31,44,31,44,30,200,31,209,31,209,30,149,31,231,31,231,30,100,31,188,31,235,31,112,31,142,31,99,31,242,31,213,31,47,31,200,31,119,31,119,30,115,31,12,31,98,31,69,31,236,31,1,31,124,31,115,31,115,30,122,31,90,31,249,31,13,31,13,30,13,29,13,28,174,31,60,31,221,31,12,31,51,31,150,31,180,31,186,31,204,31,204,30,200,31,115,31,41,31,99,31,63,31,63,30,156,31,213,31,231,31,231,30,178,31,238,31,191,31,12,31,152,31,230,31,114,31,114,30,64,31,248,31,233,31,233,30,98,31,130,31,29,31,29,30,215,31,120,31,120,30,131,31,131,30,82,31,65,31,63,31,124,31,181,31,245,31,193,31,41,31,134,31,217,31,106,31,21,31,37,31,37,30,8,31,220,31,88,31,88,30,145,31,45,31,234,31,234,30,70,31,51,31,200,31,99,31,24,31,61,31,61,30,13,31,214,31,214,30,184,31,184,30,201,31,164,31,246,31,51,31,190,31,205,31,110,31,45,31,52,31,177,31,42,31,120,31,60,31,164,31,252,31,253,31,192,31,86,31,66,31,66,30,56,31,6,31,211,31,211,30,213,31,139,31,139,30,28,31,115,31,105,31,191,31,201,31,34,31,34,30,34,29,42,31,83,31,83,30,125,31,145,31,61,31,150,31,42,31,102,31,227,31,113,31,113,30,113,29,135,31,119,31,189,31,189,30,139,31,137,31,137,30,143,31,161,31,28,31,218,31,189,31,139,31,139,30,53,31,53,30,136,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
