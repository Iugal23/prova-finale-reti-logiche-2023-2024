-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 684;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (200,0,0,0,229,0,30,0,123,0,124,0,0,0,155,0,0,0,48,0,173,0,108,0,95,0,27,0,181,0,135,0,167,0,69,0,0,0,0,0,98,0,112,0,169,0,204,0,34,0,19,0,155,0,173,0,230,0,90,0,205,0,37,0,0,0,0,0,26,0,254,0,47,0,0,0,0,0,74,0,0,0,23,0,17,0,37,0,245,0,38,0,110,0,233,0,0,0,233,0,45,0,117,0,183,0,108,0,125,0,230,0,0,0,157,0,123,0,145,0,16,0,138,0,182,0,170,0,186,0,176,0,216,0,0,0,132,0,156,0,191,0,20,0,223,0,9,0,94,0,224,0,222,0,0,0,0,0,0,0,67,0,4,0,0,0,104,0,140,0,136,0,0,0,197,0,244,0,195,0,80,0,0,0,29,0,60,0,0,0,53,0,243,0,230,0,0,0,178,0,128,0,237,0,221,0,170,0,0,0,86,0,201,0,30,0,202,0,188,0,60,0,148,0,167,0,159,0,221,0,253,0,56,0,96,0,105,0,27,0,90,0,78,0,88,0,222,0,180,0,214,0,112,0,0,0,0,0,141,0,253,0,169,0,0,0,171,0,163,0,197,0,94,0,109,0,0,0,0,0,21,0,147,0,66,0,0,0,106,0,78,0,127,0,0,0,79,0,90,0,49,0,64,0,0,0,73,0,230,0,203,0,215,0,63,0,250,0,193,0,126,0,124,0,98,0,183,0,194,0,17,0,63,0,129,0,198,0,226,0,185,0,74,0,255,0,0,0,56,0,107,0,16,0,132,0,177,0,76,0,193,0,15,0,164,0,0,0,17,0,238,0,210,0,186,0,213,0,0,0,63,0,188,0,177,0,117,0,232,0,96,0,232,0,167,0,212,0,231,0,179,0,134,0,50,0,180,0,180,0,0,0,0,0,4,0,130,0,20,0,212,0,153,0,0,0,78,0,0,0,173,0,89,0,0,0,228,0,74,0,114,0,20,0,19,0,0,0,169,0,71,0,25,0,155,0,0,0,97,0,146,0,249,0,119,0,54,0,37,0,228,0,54,0,226,0,37,0,213,0,0,0,46,0,167,0,166,0,93,0,149,0,0,0,0,0,9,0,2,0,0,0,44,0,164,0,248,0,170,0,38,0,43,0,107,0,105,0,212,0,0,0,73,0,0,0,0,0,13,0,94,0,133,0,95,0,246,0,92,0,46,0,123,0,252,0,0,0,18,0,223,0,78,0,188,0,236,0,0,0,0,0,0,0,0,0,72,0,128,0,0,0,117,0,168,0,23,0,67,0,84,0,189,0,46,0,11,0,0,0,19,0,0,0,84,0,217,0,29,0,55,0,197,0,181,0,223,0,182,0,105,0,253,0,0,0,0,0,208,0,215,0,62,0,244,0,192,0,105,0,212,0,221,0,33,0,121,0,221,0,109,0,137,0,116,0,214,0,80,0,85,0,175,0,63,0,234,0,143,0,9,0,173,0,0,0,0,0,87,0,0,0,0,0,0,0,0,0,153,0,34,0,254,0,38,0,35,0,0,0,125,0,23,0,70,0,66,0,148,0,0,0,213,0,140,0,0,0,216,0,40,0,0,0,93,0,236,0,0,0,113,0,244,0,193,0,185,0,209,0,0,0,163,0,112,0,3,0,192,0,53,0,49,0,0,0,179,0,63,0,74,0,231,0,0,0,0,0,0,0,255,0,58,0,70,0,97,0,37,0,222,0,67,0,0,0,141,0,0,0,91,0,156,0,46,0,133,0,200,0,252,0,6,0,130,0,28,0,21,0,161,0,234,0,177,0,192,0,60,0,129,0,0,0,237,0,158,0,230,0,52,0,215,0,136,0,117,0,160,0,87,0,214,0,0,0,6,0,0,0,223,0,51,0,107,0,164,0,237,0,196,0,102,0,0,0,148,0,187,0,254,0,208,0,104,0,0,0,56,0,0,0,177,0,0,0,18,0,14,0,86,0,35,0,198,0,218,0,241,0,214,0,42,0,65,0,0,0,155,0,237,0,0,0,97,0,0,0,0,0,235,0,183,0,87,0,63,0,77,0,160,0,162,0,128,0,18,0,179,0,249,0,150,0,215,0,83,0,137,0,45,0,231,0,111,0,71,0,45,0,225,0,3,0,201,0,222,0,236,0,192,0,0,0,111,0,232,0,49,0,242,0,0,0,114,0,0,0,18,0,0,0,194,0,247,0,252,0,52,0,0,0,144,0,227,0,154,0,228,0,0,0,207,0,8,0,97,0,159,0,73,0,103,0,183,0,107,0,0,0,204,0,201,0,0,0,52,0,42,0,50,0,0,0,29,0,0,0,124,0,0,0,178,0,223,0,225,0,143,0,254,0,166,0,168,0,115,0,40,0,49,0,251,0,0,0,213,0,195,0,252,0,169,0,149,0,88,0,129,0,251,0,19,0,142,0,187,0,55,0,140,0,149,0,48,0,8,0,0,0,124,0,106,0,218,0,0,0,0,0,164,0,0,0,219,0,0,0,213,0,33,0,121,0,0,0,48,0,0,0,139,0,37,0,247,0,71,0,221,0,51,0,0,0,0,0,212,0,95,0,199,0,0,0,151,0,47,0,214,0,150,0,0,0,115,0,87,0,222,0,64,0,92,0,98,0,73,0,56,0,62,0,242,0,141,0,215,0,124,0,160,0,0,0,55,0,0,0,39,0,237,0,49,0,139,0,118,0,0,0,132,0,115,0,8,0,0,0,107,0,226,0,175,0,239,0,248,0,134,0,13,0,196,0,26,0,0,0,173,0,254,0,140,0,119,0,0,0,0,0,0,0,236,0,85,0,243,0,0,0,100,0,237,0,164,0,6,0,139,0,0,0,148,0,26,0,204,0,119,0,239,0,226,0,69,0,25,0,150,0,195,0,139,0,1,0,0,0,0,0,62,0,137,0,23,0,250,0,0,0,53,0,39,0,161,0,0,0,212,0,187,0,116,0,30,0,0,0,38,0,103,0,119,0,0,0,0,0,244,0,251,0,52,0,162,0,215,0,58,0,0,0,216,0,64,0,20,0,59,0,0,0,120,0,33,0,0,0);
signal scenario_full  : scenario_type := (200,31,200,30,229,31,30,31,123,31,124,31,124,30,155,31,155,30,48,31,173,31,108,31,95,31,27,31,181,31,135,31,167,31,69,31,69,30,69,29,98,31,112,31,169,31,204,31,34,31,19,31,155,31,173,31,230,31,90,31,205,31,37,31,37,30,37,29,26,31,254,31,47,31,47,30,47,29,74,31,74,30,23,31,17,31,37,31,245,31,38,31,110,31,233,31,233,30,233,31,45,31,117,31,183,31,108,31,125,31,230,31,230,30,157,31,123,31,145,31,16,31,138,31,182,31,170,31,186,31,176,31,216,31,216,30,132,31,156,31,191,31,20,31,223,31,9,31,94,31,224,31,222,31,222,30,222,29,222,28,67,31,4,31,4,30,104,31,140,31,136,31,136,30,197,31,244,31,195,31,80,31,80,30,29,31,60,31,60,30,53,31,243,31,230,31,230,30,178,31,128,31,237,31,221,31,170,31,170,30,86,31,201,31,30,31,202,31,188,31,60,31,148,31,167,31,159,31,221,31,253,31,56,31,96,31,105,31,27,31,90,31,78,31,88,31,222,31,180,31,214,31,112,31,112,30,112,29,141,31,253,31,169,31,169,30,171,31,163,31,197,31,94,31,109,31,109,30,109,29,21,31,147,31,66,31,66,30,106,31,78,31,127,31,127,30,79,31,90,31,49,31,64,31,64,30,73,31,230,31,203,31,215,31,63,31,250,31,193,31,126,31,124,31,98,31,183,31,194,31,17,31,63,31,129,31,198,31,226,31,185,31,74,31,255,31,255,30,56,31,107,31,16,31,132,31,177,31,76,31,193,31,15,31,164,31,164,30,17,31,238,31,210,31,186,31,213,31,213,30,63,31,188,31,177,31,117,31,232,31,96,31,232,31,167,31,212,31,231,31,179,31,134,31,50,31,180,31,180,31,180,30,180,29,4,31,130,31,20,31,212,31,153,31,153,30,78,31,78,30,173,31,89,31,89,30,228,31,74,31,114,31,20,31,19,31,19,30,169,31,71,31,25,31,155,31,155,30,97,31,146,31,249,31,119,31,54,31,37,31,228,31,54,31,226,31,37,31,213,31,213,30,46,31,167,31,166,31,93,31,149,31,149,30,149,29,9,31,2,31,2,30,44,31,164,31,248,31,170,31,38,31,43,31,107,31,105,31,212,31,212,30,73,31,73,30,73,29,13,31,94,31,133,31,95,31,246,31,92,31,46,31,123,31,252,31,252,30,18,31,223,31,78,31,188,31,236,31,236,30,236,29,236,28,236,27,72,31,128,31,128,30,117,31,168,31,23,31,67,31,84,31,189,31,46,31,11,31,11,30,19,31,19,30,84,31,217,31,29,31,55,31,197,31,181,31,223,31,182,31,105,31,253,31,253,30,253,29,208,31,215,31,62,31,244,31,192,31,105,31,212,31,221,31,33,31,121,31,221,31,109,31,137,31,116,31,214,31,80,31,85,31,175,31,63,31,234,31,143,31,9,31,173,31,173,30,173,29,87,31,87,30,87,29,87,28,87,27,153,31,34,31,254,31,38,31,35,31,35,30,125,31,23,31,70,31,66,31,148,31,148,30,213,31,140,31,140,30,216,31,40,31,40,30,93,31,236,31,236,30,113,31,244,31,193,31,185,31,209,31,209,30,163,31,112,31,3,31,192,31,53,31,49,31,49,30,179,31,63,31,74,31,231,31,231,30,231,29,231,28,255,31,58,31,70,31,97,31,37,31,222,31,67,31,67,30,141,31,141,30,91,31,156,31,46,31,133,31,200,31,252,31,6,31,130,31,28,31,21,31,161,31,234,31,177,31,192,31,60,31,129,31,129,30,237,31,158,31,230,31,52,31,215,31,136,31,117,31,160,31,87,31,214,31,214,30,6,31,6,30,223,31,51,31,107,31,164,31,237,31,196,31,102,31,102,30,148,31,187,31,254,31,208,31,104,31,104,30,56,31,56,30,177,31,177,30,18,31,14,31,86,31,35,31,198,31,218,31,241,31,214,31,42,31,65,31,65,30,155,31,237,31,237,30,97,31,97,30,97,29,235,31,183,31,87,31,63,31,77,31,160,31,162,31,128,31,18,31,179,31,249,31,150,31,215,31,83,31,137,31,45,31,231,31,111,31,71,31,45,31,225,31,3,31,201,31,222,31,236,31,192,31,192,30,111,31,232,31,49,31,242,31,242,30,114,31,114,30,18,31,18,30,194,31,247,31,252,31,52,31,52,30,144,31,227,31,154,31,228,31,228,30,207,31,8,31,97,31,159,31,73,31,103,31,183,31,107,31,107,30,204,31,201,31,201,30,52,31,42,31,50,31,50,30,29,31,29,30,124,31,124,30,178,31,223,31,225,31,143,31,254,31,166,31,168,31,115,31,40,31,49,31,251,31,251,30,213,31,195,31,252,31,169,31,149,31,88,31,129,31,251,31,19,31,142,31,187,31,55,31,140,31,149,31,48,31,8,31,8,30,124,31,106,31,218,31,218,30,218,29,164,31,164,30,219,31,219,30,213,31,33,31,121,31,121,30,48,31,48,30,139,31,37,31,247,31,71,31,221,31,51,31,51,30,51,29,212,31,95,31,199,31,199,30,151,31,47,31,214,31,150,31,150,30,115,31,87,31,222,31,64,31,92,31,98,31,73,31,56,31,62,31,242,31,141,31,215,31,124,31,160,31,160,30,55,31,55,30,39,31,237,31,49,31,139,31,118,31,118,30,132,31,115,31,8,31,8,30,107,31,226,31,175,31,239,31,248,31,134,31,13,31,196,31,26,31,26,30,173,31,254,31,140,31,119,31,119,30,119,29,119,28,236,31,85,31,243,31,243,30,100,31,237,31,164,31,6,31,139,31,139,30,148,31,26,31,204,31,119,31,239,31,226,31,69,31,25,31,150,31,195,31,139,31,1,31,1,30,1,29,62,31,137,31,23,31,250,31,250,30,53,31,39,31,161,31,161,30,212,31,187,31,116,31,30,31,30,30,38,31,103,31,119,31,119,30,119,29,244,31,251,31,52,31,162,31,215,31,58,31,58,30,216,31,64,31,20,31,59,31,59,30,120,31,33,31,33,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
