-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 272;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (180,0,172,0,0,0,124,0,123,0,163,0,186,0,204,0,239,0,74,0,253,0,79,0,1,0,35,0,125,0,248,0,84,0,208,0,7,0,215,0,171,0,0,0,24,0,0,0,119,0,38,0,200,0,0,0,233,0,213,0,44,0,199,0,22,0,234,0,0,0,189,0,22,0,0,0,0,0,255,0,196,0,141,0,182,0,250,0,145,0,250,0,69,0,238,0,166,0,0,0,0,0,0,0,21,0,142,0,198,0,174,0,132,0,21,0,57,0,53,0,0,0,23,0,8,0,254,0,245,0,93,0,0,0,90,0,0,0,111,0,0,0,32,0,159,0,57,0,82,0,225,0,212,0,153,0,63,0,15,0,236,0,82,0,33,0,225,0,32,0,116,0,14,0,186,0,0,0,162,0,237,0,163,0,225,0,214,0,246,0,141,0,83,0,106,0,238,0,82,0,254,0,238,0,48,0,0,0,199,0,201,0,0,0,0,0,179,0,181,0,174,0,234,0,171,0,0,0,31,0,54,0,158,0,86,0,0,0,0,0,28,0,194,0,212,0,37,0,0,0,0,0,193,0,0,0,243,0,0,0,55,0,224,0,218,0,245,0,128,0,202,0,139,0,213,0,23,0,241,0,241,0,224,0,82,0,250,0,170,0,180,0,173,0,0,0,191,0,0,0,13,0,7,0,93,0,134,0,27,0,0,0,0,0,145,0,220,0,211,0,64,0,0,0,135,0,77,0,115,0,75,0,101,0,184,0,232,0,90,0,189,0,236,0,0,0,229,0,243,0,93,0,0,0,0,0,227,0,70,0,19,0,183,0,0,0,188,0,207,0,153,0,224,0,26,0,89,0,32,0,70,0,0,0,0,0,153,0,0,0,71,0,234,0,66,0,166,0,0,0,223,0,103,0,223,0,215,0,17,0,113,0,126,0,171,0,156,0,68,0,60,0,0,0,85,0,215,0,0,0,52,0,72,0,240,0,87,0,0,0,210,0,94,0,182,0,251,0,99,0,138,0,140,0,0,0,41,0,49,0,0,0,52,0,0,0,159,0,19,0,58,0,180,0,0,0,153,0,139,0,0,0,184,0,125,0,169,0,182,0,57,0,146,0,187,0,7,0,204,0,19,0,117,0,152,0,108,0,5,0,23,0,0,0,106,0,147,0,160,0,78,0,0,0,172,0,0,0,253,0,17,0,254,0,0,0,213,0,81,0,168,0,107,0);
signal scenario_full  : scenario_type := (180,31,172,31,172,30,124,31,123,31,163,31,186,31,204,31,239,31,74,31,253,31,79,31,1,31,35,31,125,31,248,31,84,31,208,31,7,31,215,31,171,31,171,30,24,31,24,30,119,31,38,31,200,31,200,30,233,31,213,31,44,31,199,31,22,31,234,31,234,30,189,31,22,31,22,30,22,29,255,31,196,31,141,31,182,31,250,31,145,31,250,31,69,31,238,31,166,31,166,30,166,29,166,28,21,31,142,31,198,31,174,31,132,31,21,31,57,31,53,31,53,30,23,31,8,31,254,31,245,31,93,31,93,30,90,31,90,30,111,31,111,30,32,31,159,31,57,31,82,31,225,31,212,31,153,31,63,31,15,31,236,31,82,31,33,31,225,31,32,31,116,31,14,31,186,31,186,30,162,31,237,31,163,31,225,31,214,31,246,31,141,31,83,31,106,31,238,31,82,31,254,31,238,31,48,31,48,30,199,31,201,31,201,30,201,29,179,31,181,31,174,31,234,31,171,31,171,30,31,31,54,31,158,31,86,31,86,30,86,29,28,31,194,31,212,31,37,31,37,30,37,29,193,31,193,30,243,31,243,30,55,31,224,31,218,31,245,31,128,31,202,31,139,31,213,31,23,31,241,31,241,31,224,31,82,31,250,31,170,31,180,31,173,31,173,30,191,31,191,30,13,31,7,31,93,31,134,31,27,31,27,30,27,29,145,31,220,31,211,31,64,31,64,30,135,31,77,31,115,31,75,31,101,31,184,31,232,31,90,31,189,31,236,31,236,30,229,31,243,31,93,31,93,30,93,29,227,31,70,31,19,31,183,31,183,30,188,31,207,31,153,31,224,31,26,31,89,31,32,31,70,31,70,30,70,29,153,31,153,30,71,31,234,31,66,31,166,31,166,30,223,31,103,31,223,31,215,31,17,31,113,31,126,31,171,31,156,31,68,31,60,31,60,30,85,31,215,31,215,30,52,31,72,31,240,31,87,31,87,30,210,31,94,31,182,31,251,31,99,31,138,31,140,31,140,30,41,31,49,31,49,30,52,31,52,30,159,31,19,31,58,31,180,31,180,30,153,31,139,31,139,30,184,31,125,31,169,31,182,31,57,31,146,31,187,31,7,31,204,31,19,31,117,31,152,31,108,31,5,31,23,31,23,30,106,31,147,31,160,31,78,31,78,30,172,31,172,30,253,31,17,31,254,31,254,30,213,31,81,31,168,31,107,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
