-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 356;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (24,0,60,0,104,0,254,0,122,0,78,0,149,0,140,0,0,0,0,0,255,0,0,0,46,0,52,0,245,0,0,0,5,0,49,0,29,0,32,0,74,0,181,0,0,0,56,0,151,0,92,0,254,0,218,0,234,0,101,0,0,0,224,0,253,0,86,0,0,0,242,0,0,0,0,0,0,0,220,0,57,0,46,0,2,0,0,0,13,0,235,0,208,0,145,0,66,0,18,0,248,0,127,0,79,0,30,0,47,0,188,0,254,0,58,0,0,0,99,0,21,0,217,0,96,0,81,0,0,0,184,0,0,0,0,0,0,0,214,0,79,0,188,0,140,0,103,0,253,0,0,0,76,0,5,0,0,0,176,0,24,0,8,0,231,0,0,0,248,0,0,0,233,0,87,0,152,0,197,0,152,0,229,0,0,0,65,0,192,0,0,0,65,0,108,0,86,0,0,0,40,0,39,0,213,0,154,0,0,0,132,0,44,0,118,0,168,0,92,0,53,0,96,0,153,0,188,0,0,0,0,0,100,0,161,0,170,0,219,0,68,0,0,0,227,0,196,0,0,0,61,0,66,0,234,0,207,0,60,0,164,0,202,0,106,0,0,0,114,0,247,0,183,0,38,0,238,0,255,0,143,0,249,0,11,0,123,0,0,0,207,0,184,0,165,0,163,0,152,0,67,0,189,0,150,0,171,0,227,0,0,0,0,0,201,0,215,0,66,0,19,0,237,0,95,0,155,0,55,0,93,0,44,0,123,0,0,0,0,0,0,0,133,0,183,0,91,0,23,0,116,0,73,0,194,0,194,0,68,0,87,0,180,0,0,0,11,0,93,0,0,0,50,0,2,0,0,0,209,0,67,0,225,0,43,0,90,0,255,0,200,0,234,0,118,0,0,0,152,0,127,0,134,0,107,0,0,0,0,0,0,0,169,0,0,0,87,0,215,0,18,0,0,0,191,0,80,0,165,0,0,0,206,0,1,0,184,0,0,0,244,0,62,0,0,0,0,0,232,0,0,0,178,0,236,0,42,0,199,0,0,0,0,0,143,0,0,0,233,0,231,0,0,0,199,0,0,0,0,0,67,0,165,0,208,0,54,0,170,0,199,0,157,0,144,0,211,0,100,0,0,0,93,0,198,0,0,0,9,0,108,0,197,0,55,0,232,0,15,0,225,0,0,0,141,0,0,0,203,0,80,0,132,0,0,0,170,0,53,0,186,0,6,0,181,0,89,0,0,0,0,0,217,0,27,0,85,0,76,0,0,0,0,0,141,0,122,0,157,0,34,0,124,0,0,0,235,0,64,0,130,0,35,0,34,0,141,0,0,0,130,0,113,0,91,0,58,0,0,0,193,0,13,0,0,0,191,0,252,0,120,0,0,0,0,0,60,0,136,0,146,0,213,0,0,0,197,0,204,0,116,0,188,0,56,0,187,0,115,0,250,0,140,0,233,0,133,0,96,0,0,0,56,0,0,0,105,0,252,0,85,0,233,0,0,0,156,0,0,0,247,0,142,0,188,0,141,0,0,0,163,0,170,0,139,0,131,0,0,0,44,0,47,0,234,0,0,0,37,0,0,0,0,0,66,0,101,0,5,0,178,0);
signal scenario_full  : scenario_type := (24,31,60,31,104,31,254,31,122,31,78,31,149,31,140,31,140,30,140,29,255,31,255,30,46,31,52,31,245,31,245,30,5,31,49,31,29,31,32,31,74,31,181,31,181,30,56,31,151,31,92,31,254,31,218,31,234,31,101,31,101,30,224,31,253,31,86,31,86,30,242,31,242,30,242,29,242,28,220,31,57,31,46,31,2,31,2,30,13,31,235,31,208,31,145,31,66,31,18,31,248,31,127,31,79,31,30,31,47,31,188,31,254,31,58,31,58,30,99,31,21,31,217,31,96,31,81,31,81,30,184,31,184,30,184,29,184,28,214,31,79,31,188,31,140,31,103,31,253,31,253,30,76,31,5,31,5,30,176,31,24,31,8,31,231,31,231,30,248,31,248,30,233,31,87,31,152,31,197,31,152,31,229,31,229,30,65,31,192,31,192,30,65,31,108,31,86,31,86,30,40,31,39,31,213,31,154,31,154,30,132,31,44,31,118,31,168,31,92,31,53,31,96,31,153,31,188,31,188,30,188,29,100,31,161,31,170,31,219,31,68,31,68,30,227,31,196,31,196,30,61,31,66,31,234,31,207,31,60,31,164,31,202,31,106,31,106,30,114,31,247,31,183,31,38,31,238,31,255,31,143,31,249,31,11,31,123,31,123,30,207,31,184,31,165,31,163,31,152,31,67,31,189,31,150,31,171,31,227,31,227,30,227,29,201,31,215,31,66,31,19,31,237,31,95,31,155,31,55,31,93,31,44,31,123,31,123,30,123,29,123,28,133,31,183,31,91,31,23,31,116,31,73,31,194,31,194,31,68,31,87,31,180,31,180,30,11,31,93,31,93,30,50,31,2,31,2,30,209,31,67,31,225,31,43,31,90,31,255,31,200,31,234,31,118,31,118,30,152,31,127,31,134,31,107,31,107,30,107,29,107,28,169,31,169,30,87,31,215,31,18,31,18,30,191,31,80,31,165,31,165,30,206,31,1,31,184,31,184,30,244,31,62,31,62,30,62,29,232,31,232,30,178,31,236,31,42,31,199,31,199,30,199,29,143,31,143,30,233,31,231,31,231,30,199,31,199,30,199,29,67,31,165,31,208,31,54,31,170,31,199,31,157,31,144,31,211,31,100,31,100,30,93,31,198,31,198,30,9,31,108,31,197,31,55,31,232,31,15,31,225,31,225,30,141,31,141,30,203,31,80,31,132,31,132,30,170,31,53,31,186,31,6,31,181,31,89,31,89,30,89,29,217,31,27,31,85,31,76,31,76,30,76,29,141,31,122,31,157,31,34,31,124,31,124,30,235,31,64,31,130,31,35,31,34,31,141,31,141,30,130,31,113,31,91,31,58,31,58,30,193,31,13,31,13,30,191,31,252,31,120,31,120,30,120,29,60,31,136,31,146,31,213,31,213,30,197,31,204,31,116,31,188,31,56,31,187,31,115,31,250,31,140,31,233,31,133,31,96,31,96,30,56,31,56,30,105,31,252,31,85,31,233,31,233,30,156,31,156,30,247,31,142,31,188,31,141,31,141,30,163,31,170,31,139,31,131,31,131,30,44,31,47,31,234,31,234,30,37,31,37,30,37,29,66,31,101,31,5,31,178,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
