-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 951;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (110,0,241,0,0,0,193,0,61,0,76,0,0,0,97,0,187,0,61,0,98,0,0,0,181,0,206,0,38,0,68,0,61,0,211,0,59,0,0,0,195,0,40,0,0,0,115,0,243,0,0,0,48,0,188,0,233,0,0,0,7,0,111,0,24,0,25,0,84,0,175,0,56,0,210,0,0,0,0,0,150,0,160,0,156,0,34,0,0,0,79,0,246,0,44,0,177,0,0,0,164,0,0,0,255,0,30,0,167,0,0,0,133,0,236,0,150,0,2,0,162,0,129,0,131,0,0,0,117,0,146,0,85,0,100,0,149,0,255,0,8,0,197,0,99,0,6,0,0,0,100,0,12,0,232,0,206,0,46,0,118,0,0,0,0,0,9,0,0,0,66,0,253,0,115,0,87,0,0,0,147,0,105,0,249,0,209,0,0,0,228,0,22,0,14,0,16,0,0,0,179,0,212,0,51,0,15,0,191,0,160,0,194,0,12,0,102,0,240,0,18,0,169,0,0,0,146,0,0,0,179,0,15,0,0,0,0,0,176,0,0,0,190,0,81,0,168,0,184,0,0,0,114,0,5,0,202,0,194,0,141,0,38,0,181,0,220,0,228,0,216,0,108,0,0,0,0,0,166,0,67,0,182,0,76,0,0,0,135,0,0,0,107,0,204,0,128,0,0,0,108,0,0,0,77,0,84,0,0,0,0,0,54,0,10,0,183,0,0,0,76,0,233,0,145,0,146,0,0,0,0,0,211,0,176,0,0,0,0,0,161,0,24,0,0,0,59,0,128,0,181,0,186,0,132,0,76,0,199,0,0,0,200,0,138,0,0,0,29,0,101,0,133,0,0,0,178,0,0,0,209,0,101,0,2,0,158,0,0,0,102,0,55,0,159,0,243,0,18,0,197,0,198,0,245,0,39,0,246,0,141,0,0,0,175,0,133,0,127,0,91,0,163,0,48,0,110,0,60,0,0,0,110,0,0,0,64,0,17,0,50,0,206,0,48,0,141,0,58,0,32,0,0,0,183,0,0,0,106,0,136,0,221,0,191,0,0,0,54,0,248,0,231,0,28,0,52,0,77,0,202,0,0,0,231,0,32,0,0,0,0,0,92,0,189,0,43,0,137,0,79,0,183,0,255,0,36,0,210,0,88,0,111,0,91,0,0,0,0,0,51,0,185,0,223,0,63,0,175,0,71,0,2,0,0,0,198,0,167,0,0,0,208,0,180,0,127,0,0,0,78,0,207,0,27,0,0,0,99,0,232,0,6,0,65,0,161,0,30,0,198,0,185,0,177,0,247,0,0,0,127,0,193,0,234,0,201,0,133,0,38,0,113,0,0,0,0,0,0,0,153,0,185,0,130,0,10,0,50,0,65,0,255,0,0,0,195,0,197,0,0,0,0,0,252,0,25,0,186,0,0,0,0,0,130,0,189,0,250,0,153,0,240,0,39,0,143,0,213,0,135,0,151,0,215,0,223,0,75,0,255,0,45,0,0,0,245,0,222,0,184,0,171,0,8,0,236,0,240,0,54,0,155,0,107,0,34,0,210,0,244,0,122,0,0,0,52,0,0,0,34,0,176,0,140,0,0,0,116,0,44,0,251,0,114,0,237,0,164,0,251,0,109,0,0,0,34,0,186,0,0,0,215,0,20,0,142,0,25,0,2,0,2,0,0,0,79,0,196,0,141,0,0,0,9,0,81,0,58,0,0,0,65,0,115,0,129,0,199,0,251,0,248,0,0,0,94,0,198,0,73,0,118,0,123,0,0,0,176,0,94,0,56,0,0,0,204,0,142,0,196,0,49,0,61,0,61,0,102,0,54,0,209,0,77,0,193,0,202,0,219,0,0,0,0,0,149,0,98,0,8,0,143,0,109,0,79,0,0,0,138,0,164,0,102,0,53,0,167,0,141,0,54,0,172,0,250,0,91,0,234,0,208,0,0,0,233,0,188,0,217,0,180,0,226,0,113,0,55,0,238,0,108,0,20,0,255,0,180,0,0,0,23,0,0,0,61,0,0,0,202,0,19,0,227,0,102,0,222,0,46,0,181,0,112,0,121,0,0,0,5,0,69,0,126,0,145,0,79,0,207,0,172,0,0,0,156,0,188,0,8,0,0,0,0,0,165,0,200,0,0,0,1,0,118,0,49,0,178,0,204,0,192,0,168,0,136,0,29,0,76,0,10,0,0,0,39,0,0,0,81,0,0,0,228,0,111,0,232,0,243,0,208,0,31,0,0,0,0,0,252,0,0,0,0,0,0,0,226,0,0,0,0,0,104,0,0,0,34,0,0,0,173,0,145,0,0,0,69,0,166,0,25,0,118,0,18,0,218,0,115,0,192,0,254,0,127,0,0,0,0,0,0,0,104,0,38,0,0,0,45,0,32,0,39,0,228,0,238,0,178,0,170,0,150,0,11,0,63,0,149,0,33,0,0,0,3,0,106,0,220,0,63,0,0,0,214,0,0,0,0,0,99,0,151,0,84,0,235,0,53,0,89,0,75,0,120,0,250,0,42,0,155,0,54,0,192,0,37,0,102,0,35,0,138,0,0,0,253,0,0,0,186,0,59,0,117,0,0,0,96,0,0,0,191,0,133,0,0,0,142,0,115,0,45,0,91,0,85,0,0,0,229,0,147,0,121,0,34,0,57,0,13,0,159,0,181,0,161,0,244,0,112,0,62,0,96,0,0,0,81,0,0,0,37,0,46,0,0,0,130,0,129,0,67,0,239,0,0,0,114,0,43,0,0,0,148,0,0,0,62,0,130,0,0,0,78,0,253,0,87,0,91,0,81,0,128,0,0,0,187,0,185,0,43,0,80,0,27,0,0,0,37,0,6,0,170,0,153,0,27,0,173,0,31,0,0,0,88,0,130,0,0,0,251,0,4,0,17,0,230,0,0,0,243,0,185,0,166,0,0,0,227,0,17,0,165,0,0,0,8,0,109,0,62,0,5,0,4,0,31,0,151,0,0,0,0,0,83,0,196,0,0,0,141,0,0,0,0,0,0,0,91,0,195,0,110,0,245,0,0,0,0,0,176,0,55,0,128,0,218,0,145,0,0,0,192,0,0,0,0,0,66,0,0,0,0,0,144,0,0,0,9,0,0,0,215,0,43,0,188,0,143,0,180,0,175,0,127,0,77,0,56,0,0,0,0,0,210,0,19,0,197,0,0,0,0,0,141,0,9,0,101,0,92,0,0,0,167,0,12,0,233,0,0,0,137,0,21,0,45,0,0,0,53,0,220,0,84,0,0,0,225,0,70,0,68,0,74,0,111,0,0,0,14,0,99,0,185,0,45,0,0,0,0,0,233,0,227,0,0,0,121,0,171,0,0,0,186,0,156,0,136,0,0,0,202,0,0,0,0,0,151,0,65,0,48,0,0,0,72,0,169,0,12,0,50,0,179,0,119,0,40,0,95,0,0,0,30,0,24,0,185,0,0,0,2,0,15,0,148,0,134,0,169,0,0,0,0,0,149,0,0,0,59,0,219,0,246,0,54,0,96,0,240,0,21,0,247,0,0,0,93,0,0,0,167,0,173,0,152,0,0,0,253,0,158,0,187,0,175,0,0,0,75,0,0,0,25,0,254,0,129,0,73,0,246,0,138,0,174,0,18,0,0,0,232,0,159,0,0,0,39,0,179,0,198,0,75,0,253,0,5,0,0,0,72,0,153,0,85,0,36,0,51,0,78,0,172,0,122,0,0,0,97,0,116,0,63,0,77,0,0,0,35,0,0,0,203,0,180,0,205,0,132,0,29,0,0,0,0,0,209,0,255,0,164,0,58,0,46,0,130,0,22,0,226,0,74,0,78,0,0,0,54,0,0,0,210,0,0,0,20,0,145,0,0,0,225,0,209,0,0,0,12,0,238,0,0,0,251,0,11,0,95,0,68,0,17,0,0,0,104,0,125,0,119,0,0,0,43,0,131,0,161,0,68,0,245,0,181,0,177,0,48,0,0,0,48,0,209,0,0,0,0,0,39,0,0,0,0,0,168,0,220,0,87,0,71,0,109,0,210,0,214,0,181,0,33,0,60,0,173,0,75,0,0,0,8,0,165,0,229,0,15,0,199,0,221,0,156,0,188,0,27,0,0,0,0,0,0,0,249,0,17,0,89,0,200,0,130,0,244,0,0,0,125,0,119,0,165,0,212,0,122,0,19,0,147,0,70,0,107,0,213,0,35,0,0,0,215,0,232,0,0,0,100,0,255,0,185,0,188,0,60,0,180,0,27,0,179,0,220,0,106,0,87,0,69,0,0,0);
signal scenario_full  : scenario_type := (110,31,241,31,241,30,193,31,61,31,76,31,76,30,97,31,187,31,61,31,98,31,98,30,181,31,206,31,38,31,68,31,61,31,211,31,59,31,59,30,195,31,40,31,40,30,115,31,243,31,243,30,48,31,188,31,233,31,233,30,7,31,111,31,24,31,25,31,84,31,175,31,56,31,210,31,210,30,210,29,150,31,160,31,156,31,34,31,34,30,79,31,246,31,44,31,177,31,177,30,164,31,164,30,255,31,30,31,167,31,167,30,133,31,236,31,150,31,2,31,162,31,129,31,131,31,131,30,117,31,146,31,85,31,100,31,149,31,255,31,8,31,197,31,99,31,6,31,6,30,100,31,12,31,232,31,206,31,46,31,118,31,118,30,118,29,9,31,9,30,66,31,253,31,115,31,87,31,87,30,147,31,105,31,249,31,209,31,209,30,228,31,22,31,14,31,16,31,16,30,179,31,212,31,51,31,15,31,191,31,160,31,194,31,12,31,102,31,240,31,18,31,169,31,169,30,146,31,146,30,179,31,15,31,15,30,15,29,176,31,176,30,190,31,81,31,168,31,184,31,184,30,114,31,5,31,202,31,194,31,141,31,38,31,181,31,220,31,228,31,216,31,108,31,108,30,108,29,166,31,67,31,182,31,76,31,76,30,135,31,135,30,107,31,204,31,128,31,128,30,108,31,108,30,77,31,84,31,84,30,84,29,54,31,10,31,183,31,183,30,76,31,233,31,145,31,146,31,146,30,146,29,211,31,176,31,176,30,176,29,161,31,24,31,24,30,59,31,128,31,181,31,186,31,132,31,76,31,199,31,199,30,200,31,138,31,138,30,29,31,101,31,133,31,133,30,178,31,178,30,209,31,101,31,2,31,158,31,158,30,102,31,55,31,159,31,243,31,18,31,197,31,198,31,245,31,39,31,246,31,141,31,141,30,175,31,133,31,127,31,91,31,163,31,48,31,110,31,60,31,60,30,110,31,110,30,64,31,17,31,50,31,206,31,48,31,141,31,58,31,32,31,32,30,183,31,183,30,106,31,136,31,221,31,191,31,191,30,54,31,248,31,231,31,28,31,52,31,77,31,202,31,202,30,231,31,32,31,32,30,32,29,92,31,189,31,43,31,137,31,79,31,183,31,255,31,36,31,210,31,88,31,111,31,91,31,91,30,91,29,51,31,185,31,223,31,63,31,175,31,71,31,2,31,2,30,198,31,167,31,167,30,208,31,180,31,127,31,127,30,78,31,207,31,27,31,27,30,99,31,232,31,6,31,65,31,161,31,30,31,198,31,185,31,177,31,247,31,247,30,127,31,193,31,234,31,201,31,133,31,38,31,113,31,113,30,113,29,113,28,153,31,185,31,130,31,10,31,50,31,65,31,255,31,255,30,195,31,197,31,197,30,197,29,252,31,25,31,186,31,186,30,186,29,130,31,189,31,250,31,153,31,240,31,39,31,143,31,213,31,135,31,151,31,215,31,223,31,75,31,255,31,45,31,45,30,245,31,222,31,184,31,171,31,8,31,236,31,240,31,54,31,155,31,107,31,34,31,210,31,244,31,122,31,122,30,52,31,52,30,34,31,176,31,140,31,140,30,116,31,44,31,251,31,114,31,237,31,164,31,251,31,109,31,109,30,34,31,186,31,186,30,215,31,20,31,142,31,25,31,2,31,2,31,2,30,79,31,196,31,141,31,141,30,9,31,81,31,58,31,58,30,65,31,115,31,129,31,199,31,251,31,248,31,248,30,94,31,198,31,73,31,118,31,123,31,123,30,176,31,94,31,56,31,56,30,204,31,142,31,196,31,49,31,61,31,61,31,102,31,54,31,209,31,77,31,193,31,202,31,219,31,219,30,219,29,149,31,98,31,8,31,143,31,109,31,79,31,79,30,138,31,164,31,102,31,53,31,167,31,141,31,54,31,172,31,250,31,91,31,234,31,208,31,208,30,233,31,188,31,217,31,180,31,226,31,113,31,55,31,238,31,108,31,20,31,255,31,180,31,180,30,23,31,23,30,61,31,61,30,202,31,19,31,227,31,102,31,222,31,46,31,181,31,112,31,121,31,121,30,5,31,69,31,126,31,145,31,79,31,207,31,172,31,172,30,156,31,188,31,8,31,8,30,8,29,165,31,200,31,200,30,1,31,118,31,49,31,178,31,204,31,192,31,168,31,136,31,29,31,76,31,10,31,10,30,39,31,39,30,81,31,81,30,228,31,111,31,232,31,243,31,208,31,31,31,31,30,31,29,252,31,252,30,252,29,252,28,226,31,226,30,226,29,104,31,104,30,34,31,34,30,173,31,145,31,145,30,69,31,166,31,25,31,118,31,18,31,218,31,115,31,192,31,254,31,127,31,127,30,127,29,127,28,104,31,38,31,38,30,45,31,32,31,39,31,228,31,238,31,178,31,170,31,150,31,11,31,63,31,149,31,33,31,33,30,3,31,106,31,220,31,63,31,63,30,214,31,214,30,214,29,99,31,151,31,84,31,235,31,53,31,89,31,75,31,120,31,250,31,42,31,155,31,54,31,192,31,37,31,102,31,35,31,138,31,138,30,253,31,253,30,186,31,59,31,117,31,117,30,96,31,96,30,191,31,133,31,133,30,142,31,115,31,45,31,91,31,85,31,85,30,229,31,147,31,121,31,34,31,57,31,13,31,159,31,181,31,161,31,244,31,112,31,62,31,96,31,96,30,81,31,81,30,37,31,46,31,46,30,130,31,129,31,67,31,239,31,239,30,114,31,43,31,43,30,148,31,148,30,62,31,130,31,130,30,78,31,253,31,87,31,91,31,81,31,128,31,128,30,187,31,185,31,43,31,80,31,27,31,27,30,37,31,6,31,170,31,153,31,27,31,173,31,31,31,31,30,88,31,130,31,130,30,251,31,4,31,17,31,230,31,230,30,243,31,185,31,166,31,166,30,227,31,17,31,165,31,165,30,8,31,109,31,62,31,5,31,4,31,31,31,151,31,151,30,151,29,83,31,196,31,196,30,141,31,141,30,141,29,141,28,91,31,195,31,110,31,245,31,245,30,245,29,176,31,55,31,128,31,218,31,145,31,145,30,192,31,192,30,192,29,66,31,66,30,66,29,144,31,144,30,9,31,9,30,215,31,43,31,188,31,143,31,180,31,175,31,127,31,77,31,56,31,56,30,56,29,210,31,19,31,197,31,197,30,197,29,141,31,9,31,101,31,92,31,92,30,167,31,12,31,233,31,233,30,137,31,21,31,45,31,45,30,53,31,220,31,84,31,84,30,225,31,70,31,68,31,74,31,111,31,111,30,14,31,99,31,185,31,45,31,45,30,45,29,233,31,227,31,227,30,121,31,171,31,171,30,186,31,156,31,136,31,136,30,202,31,202,30,202,29,151,31,65,31,48,31,48,30,72,31,169,31,12,31,50,31,179,31,119,31,40,31,95,31,95,30,30,31,24,31,185,31,185,30,2,31,15,31,148,31,134,31,169,31,169,30,169,29,149,31,149,30,59,31,219,31,246,31,54,31,96,31,240,31,21,31,247,31,247,30,93,31,93,30,167,31,173,31,152,31,152,30,253,31,158,31,187,31,175,31,175,30,75,31,75,30,25,31,254,31,129,31,73,31,246,31,138,31,174,31,18,31,18,30,232,31,159,31,159,30,39,31,179,31,198,31,75,31,253,31,5,31,5,30,72,31,153,31,85,31,36,31,51,31,78,31,172,31,122,31,122,30,97,31,116,31,63,31,77,31,77,30,35,31,35,30,203,31,180,31,205,31,132,31,29,31,29,30,29,29,209,31,255,31,164,31,58,31,46,31,130,31,22,31,226,31,74,31,78,31,78,30,54,31,54,30,210,31,210,30,20,31,145,31,145,30,225,31,209,31,209,30,12,31,238,31,238,30,251,31,11,31,95,31,68,31,17,31,17,30,104,31,125,31,119,31,119,30,43,31,131,31,161,31,68,31,245,31,181,31,177,31,48,31,48,30,48,31,209,31,209,30,209,29,39,31,39,30,39,29,168,31,220,31,87,31,71,31,109,31,210,31,214,31,181,31,33,31,60,31,173,31,75,31,75,30,8,31,165,31,229,31,15,31,199,31,221,31,156,31,188,31,27,31,27,30,27,29,27,28,249,31,17,31,89,31,200,31,130,31,244,31,244,30,125,31,119,31,165,31,212,31,122,31,19,31,147,31,70,31,107,31,213,31,35,31,35,30,215,31,232,31,232,30,100,31,255,31,185,31,188,31,60,31,180,31,27,31,179,31,220,31,106,31,87,31,69,31,69,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
