-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_640 is
end project_tb_640;

architecture project_tb_arch_640 of project_tb_640 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 208;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (120,0,0,0,52,0,78,0,216,0,198,0,0,0,112,0,1,0,243,0,98,0,205,0,77,0,182,0,143,0,170,0,236,0,99,0,227,0,139,0,103,0,226,0,222,0,142,0,0,0,0,0,208,0,112,0,0,0,0,0,203,0,213,0,54,0,0,0,135,0,0,0,174,0,197,0,49,0,169,0,0,0,62,0,34,0,31,0,141,0,228,0,0,0,212,0,128,0,0,0,40,0,110,0,79,0,0,0,0,0,88,0,244,0,0,0,233,0,221,0,221,0,217,0,214,0,46,0,0,0,0,0,85,0,0,0,111,0,24,0,253,0,68,0,238,0,140,0,197,0,12,0,197,0,0,0,71,0,97,0,240,0,24,0,217,0,7,0,215,0,0,0,124,0,39,0,132,0,165,0,0,0,207,0,96,0,82,0,0,0,0,0,198,0,14,0,168,0,58,0,5,0,174,0,237,0,168,0,96,0,211,0,38,0,17,0,165,0,0,0,0,0,0,0,0,0,0,0,71,0,173,0,89,0,85,0,157,0,54,0,177,0,80,0,37,0,119,0,213,0,0,0,44,0,233,0,8,0,90,0,0,0,182,0,109,0,162,0,14,0,15,0,0,0,120,0,0,0,147,0,73,0,17,0,142,0,0,0,0,0,0,0,0,0,0,0,113,0,51,0,55,0,160,0,224,0,243,0,0,0,152,0,162,0,192,0,0,0,48,0,239,0,60,0,206,0,33,0,145,0,156,0,116,0,79,0,0,0,0,0,133,0,20,0,244,0,111,0,0,0,132,0,76,0,63,0,32,0,88,0,55,0,159,0,20,0,71,0,231,0,0,0,199,0,32,0,0,0,39,0,90,0,45,0,0,0,0,0,233,0,6,0,161,0,0,0,237,0,196,0,0,0,206,0,12,0,103,0,113,0,122,0,254,0,0,0);
signal scenario_full  : scenario_type := (120,31,120,30,52,31,78,31,216,31,198,31,198,30,112,31,1,31,243,31,98,31,205,31,77,31,182,31,143,31,170,31,236,31,99,31,227,31,139,31,103,31,226,31,222,31,142,31,142,30,142,29,208,31,112,31,112,30,112,29,203,31,213,31,54,31,54,30,135,31,135,30,174,31,197,31,49,31,169,31,169,30,62,31,34,31,31,31,141,31,228,31,228,30,212,31,128,31,128,30,40,31,110,31,79,31,79,30,79,29,88,31,244,31,244,30,233,31,221,31,221,31,217,31,214,31,46,31,46,30,46,29,85,31,85,30,111,31,24,31,253,31,68,31,238,31,140,31,197,31,12,31,197,31,197,30,71,31,97,31,240,31,24,31,217,31,7,31,215,31,215,30,124,31,39,31,132,31,165,31,165,30,207,31,96,31,82,31,82,30,82,29,198,31,14,31,168,31,58,31,5,31,174,31,237,31,168,31,96,31,211,31,38,31,17,31,165,31,165,30,165,29,165,28,165,27,165,26,71,31,173,31,89,31,85,31,157,31,54,31,177,31,80,31,37,31,119,31,213,31,213,30,44,31,233,31,8,31,90,31,90,30,182,31,109,31,162,31,14,31,15,31,15,30,120,31,120,30,147,31,73,31,17,31,142,31,142,30,142,29,142,28,142,27,142,26,113,31,51,31,55,31,160,31,224,31,243,31,243,30,152,31,162,31,192,31,192,30,48,31,239,31,60,31,206,31,33,31,145,31,156,31,116,31,79,31,79,30,79,29,133,31,20,31,244,31,111,31,111,30,132,31,76,31,63,31,32,31,88,31,55,31,159,31,20,31,71,31,231,31,231,30,199,31,32,31,32,30,39,31,90,31,45,31,45,30,45,29,233,31,6,31,161,31,161,30,237,31,196,31,196,30,206,31,12,31,103,31,113,31,122,31,254,31,254,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
