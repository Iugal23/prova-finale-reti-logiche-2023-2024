-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_842 is
end project_tb_842;

architecture project_tb_arch_842 of project_tb_842 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 964;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (242,0,65,0,209,0,6,0,199,0,112,0,104,0,100,0,209,0,116,0,158,0,233,0,25,0,57,0,96,0,59,0,149,0,65,0,157,0,0,0,217,0,219,0,128,0,0,0,0,0,160,0,225,0,68,0,0,0,0,0,95,0,0,0,0,0,59,0,0,0,0,0,6,0,57,0,169,0,128,0,114,0,32,0,79,0,28,0,223,0,0,0,190,0,19,0,77,0,120,0,0,0,56,0,221,0,147,0,2,0,77,0,80,0,237,0,127,0,18,0,70,0,213,0,220,0,0,0,0,0,188,0,0,0,176,0,122,0,180,0,186,0,165,0,190,0,150,0,100,0,255,0,143,0,35,0,70,0,0,0,46,0,0,0,130,0,88,0,251,0,0,0,112,0,0,0,46,0,39,0,0,0,130,0,252,0,199,0,16,0,0,0,0,0,11,0,46,0,181,0,218,0,131,0,76,0,0,0,114,0,0,0,246,0,164,0,87,0,2,0,62,0,218,0,0,0,0,0,0,0,223,0,46,0,44,0,150,0,183,0,143,0,4,0,130,0,147,0,60,0,60,0,83,0,17,0,204,0,235,0,25,0,249,0,59,0,109,0,176,0,148,0,77,0,91,0,160,0,0,0,233,0,97,0,238,0,179,0,10,0,142,0,0,0,187,0,0,0,0,0,0,0,239,0,72,0,215,0,146,0,84,0,88,0,123,0,0,0,204,0,214,0,85,0,185,0,120,0,39,0,168,0,73,0,65,0,61,0,126,0,61,0,196,0,19,0,193,0,223,0,52,0,57,0,221,0,68,0,59,0,36,0,112,0,155,0,186,0,76,0,25,0,56,0,88,0,82,0,217,0,137,0,203,0,231,0,226,0,0,0,70,0,29,0,0,0,159,0,198,0,219,0,240,0,236,0,207,0,0,0,26,0,0,0,199,0,0,0,43,0,200,0,56,0,25,0,0,0,103,0,0,0,66,0,57,0,130,0,34,0,227,0,99,0,192,0,185,0,49,0,0,0,0,0,180,0,16,0,185,0,0,0,0,0,122,0,193,0,242,0,0,0,86,0,108,0,6,0,13,0,0,0,120,0,246,0,65,0,134,0,0,0,165,0,30,0,246,0,94,0,45,0,0,0,120,0,3,0,167,0,33,0,61,0,163,0,25,0,92,0,88,0,166,0,239,0,232,0,167,0,112,0,181,0,210,0,118,0,0,0,5,0,30,0,0,0,0,0,209,0,71,0,5,0,53,0,209,0,0,0,188,0,56,0,0,0,112,0,12,0,138,0,0,0,48,0,94,0,127,0,121,0,44,0,200,0,0,0,184,0,148,0,74,0,0,0,0,0,126,0,113,0,149,0,84,0,143,0,165,0,172,0,157,0,154,0,50,0,3,0,239,0,194,0,227,0,0,0,130,0,122,0,248,0,242,0,147,0,37,0,111,0,196,0,0,0,138,0,245,0,60,0,0,0,113,0,205,0,80,0,150,0,211,0,254,0,254,0,78,0,53,0,37,0,53,0,0,0,241,0,177,0,80,0,54,0,0,0,95,0,66,0,58,0,106,0,0,0,105,0,209,0,187,0,0,0,13,0,41,0,0,0,166,0,35,0,59,0,84,0,112,0,85,0,194,0,7,0,73,0,58,0,0,0,0,0,127,0,0,0,191,0,0,0,224,0,34,0,55,0,0,0,220,0,246,0,243,0,0,0,60,0,29,0,159,0,0,0,181,0,111,0,1,0,195,0,29,0,164,0,175,0,129,0,11,0,0,0,172,0,200,0,94,0,37,0,112,0,180,0,175,0,200,0,214,0,0,0,0,0,0,0,0,0,0,0,0,0,30,0,0,0,153,0,253,0,42,0,79,0,127,0,124,0,0,0,58,0,13,0,120,0,60,0,187,0,0,0,0,0,60,0,156,0,185,0,8,0,123,0,238,0,246,0,159,0,123,0,48,0,154,0,0,0,0,0,231,0,235,0,123,0,6,0,0,0,74,0,57,0,93,0,0,0,134,0,19,0,0,0,58,0,0,0,128,0,251,0,0,0,214,0,130,0,169,0,233,0,162,0,64,0,66,0,133,0,18,0,0,0,217,0,61,0,41,0,227,0,152,0,93,0,93,0,0,0,172,0,68,0,0,0,69,0,142,0,0,0,248,0,130,0,181,0,244,0,0,0,224,0,181,0,72,0,0,0,156,0,114,0,0,0,57,0,151,0,234,0,149,0,0,0,129,0,29,0,185,0,153,0,46,0,82,0,179,0,100,0,161,0,231,0,221,0,211,0,1,0,153,0,0,0,156,0,22,0,123,0,168,0,166,0,0,0,0,0,206,0,116,0,51,0,0,0,139,0,167,0,0,0,239,0,117,0,0,0,189,0,90,0,163,0,167,0,94,0,236,0,236,0,223,0,150,0,25,0,238,0,177,0,70,0,0,0,196,0,176,0,187,0,216,0,184,0,8,0,0,0,48,0,104,0,10,0,0,0,229,0,239,0,115,0,0,0,140,0,229,0,116,0,0,0,56,0,243,0,59,0,234,0,130,0,0,0,217,0,207,0,94,0,0,0,0,0,82,0,115,0,245,0,245,0,0,0,0,0,91,0,7,0,28,0,0,0,0,0,99,0,189,0,0,0,159,0,67,0,144,0,107,0,46,0,66,0,165,0,241,0,0,0,48,0,197,0,160,0,155,0,168,0,0,0,160,0,234,0,100,0,99,0,50,0,172,0,223,0,221,0,211,0,196,0,45,0,118,0,25,0,128,0,176,0,203,0,74,0,255,0,106,0,0,0,64,0,187,0,68,0,163,0,186,0,32,0,24,0,84,0,115,0,241,0,71,0,136,0,171,0,79,0,0,0,142,0,100,0,0,0,132,0,0,0,187,0,105,0,175,0,255,0,0,0,0,0,179,0,122,0,247,0,0,0,0,0,14,0,0,0,0,0,136,0,48,0,25,0,177,0,0,0,0,0,171,0,62,0,50,0,0,0,0,0,0,0,129,0,36,0,0,0,0,0,165,0,253,0,145,0,0,0,153,0,95,0,11,0,33,0,123,0,204,0,231,0,207,0,206,0,38,0,112,0,45,0,128,0,160,0,0,0,24,0,123,0,38,0,141,0,182,0,162,0,5,0,203,0,220,0,76,0,170,0,28,0,129,0,67,0,151,0,61,0,110,0,79,0,39,0,154,0,104,0,0,0,104,0,30,0,144,0,99,0,0,0,166,0,0,0,0,0,123,0,163,0,60,0,16,0,136,0,180,0,152,0,0,0,117,0,111,0,232,0,152,0,21,0,208,0,109,0,0,0,134,0,40,0,255,0,242,0,209,0,211,0,1,0,201,0,130,0,67,0,0,0,70,0,51,0,140,0,62,0,5,0,211,0,34,0,192,0,217,0,68,0,185,0,13,0,0,0,100,0,0,0,16,0,103,0,135,0,0,0,10,0,234,0,120,0,150,0,69,0,123,0,124,0,217,0,40,0,65,0,94,0,127,0,198,0,176,0,250,0,0,0,165,0,137,0,1,0,14,0,251,0,188,0,214,0,123,0,55,0,194,0,147,0,217,0,241,0,144,0,0,0,238,0,216,0,112,0,48,0,132,0,224,0,78,0,198,0,138,0,87,0,224,0,133,0,56,0,5,0,45,0,225,0,253,0,126,0,111,0,105,0,31,0,0,0,0,0,108,0,0,0,116,0,0,0,49,0,235,0,142,0,69,0,146,0,0,0,166,0,169,0,205,0,0,0,221,0,0,0,203,0,220,0,182,0,176,0,68,0,82,0,91,0,194,0,53,0,17,0,12,0,171,0,89,0,202,0,0,0,41,0,178,0,0,0,3,0,51,0,253,0,0,0,97,0,106,0,240,0,207,0,66,0,222,0,9,0,7,0,199,0,0,0,71,0,218,0,161,0,193,0,171,0,147,0,0,0,25,0,89,0,186,0,45,0,78,0,188,0,239,0,140,0,0,0,207,0,202,0,244,0,31,0,76,0,206,0,166,0,248,0,0,0,204,0,160,0,250,0,209,0,96,0,105,0,180,0,185,0,234,0,95,0,216,0,0,0,194,0,118,0,99,0,143,0,133,0,0,0,172,0,218,0,141,0,239,0,198,0,0,0,166,0,7,0,111,0,0,0,240,0,26,0,32,0,203,0,106,0,0,0,119,0,0,0,178,0,105,0,0,0,248,0,205,0,27,0,194,0,10,0,126,0,50,0,133,0,249,0,0,0,63,0,0,0,175,0,11,0,134,0,30,0,93,0,195,0,0,0,159,0,220,0,95,0,83,0,73,0,7,0,131,0,1,0,106,0,226,0,253,0,0,0,118,0);
signal scenario_full  : scenario_type := (242,31,65,31,209,31,6,31,199,31,112,31,104,31,100,31,209,31,116,31,158,31,233,31,25,31,57,31,96,31,59,31,149,31,65,31,157,31,157,30,217,31,219,31,128,31,128,30,128,29,160,31,225,31,68,31,68,30,68,29,95,31,95,30,95,29,59,31,59,30,59,29,6,31,57,31,169,31,128,31,114,31,32,31,79,31,28,31,223,31,223,30,190,31,19,31,77,31,120,31,120,30,56,31,221,31,147,31,2,31,77,31,80,31,237,31,127,31,18,31,70,31,213,31,220,31,220,30,220,29,188,31,188,30,176,31,122,31,180,31,186,31,165,31,190,31,150,31,100,31,255,31,143,31,35,31,70,31,70,30,46,31,46,30,130,31,88,31,251,31,251,30,112,31,112,30,46,31,39,31,39,30,130,31,252,31,199,31,16,31,16,30,16,29,11,31,46,31,181,31,218,31,131,31,76,31,76,30,114,31,114,30,246,31,164,31,87,31,2,31,62,31,218,31,218,30,218,29,218,28,223,31,46,31,44,31,150,31,183,31,143,31,4,31,130,31,147,31,60,31,60,31,83,31,17,31,204,31,235,31,25,31,249,31,59,31,109,31,176,31,148,31,77,31,91,31,160,31,160,30,233,31,97,31,238,31,179,31,10,31,142,31,142,30,187,31,187,30,187,29,187,28,239,31,72,31,215,31,146,31,84,31,88,31,123,31,123,30,204,31,214,31,85,31,185,31,120,31,39,31,168,31,73,31,65,31,61,31,126,31,61,31,196,31,19,31,193,31,223,31,52,31,57,31,221,31,68,31,59,31,36,31,112,31,155,31,186,31,76,31,25,31,56,31,88,31,82,31,217,31,137,31,203,31,231,31,226,31,226,30,70,31,29,31,29,30,159,31,198,31,219,31,240,31,236,31,207,31,207,30,26,31,26,30,199,31,199,30,43,31,200,31,56,31,25,31,25,30,103,31,103,30,66,31,57,31,130,31,34,31,227,31,99,31,192,31,185,31,49,31,49,30,49,29,180,31,16,31,185,31,185,30,185,29,122,31,193,31,242,31,242,30,86,31,108,31,6,31,13,31,13,30,120,31,246,31,65,31,134,31,134,30,165,31,30,31,246,31,94,31,45,31,45,30,120,31,3,31,167,31,33,31,61,31,163,31,25,31,92,31,88,31,166,31,239,31,232,31,167,31,112,31,181,31,210,31,118,31,118,30,5,31,30,31,30,30,30,29,209,31,71,31,5,31,53,31,209,31,209,30,188,31,56,31,56,30,112,31,12,31,138,31,138,30,48,31,94,31,127,31,121,31,44,31,200,31,200,30,184,31,148,31,74,31,74,30,74,29,126,31,113,31,149,31,84,31,143,31,165,31,172,31,157,31,154,31,50,31,3,31,239,31,194,31,227,31,227,30,130,31,122,31,248,31,242,31,147,31,37,31,111,31,196,31,196,30,138,31,245,31,60,31,60,30,113,31,205,31,80,31,150,31,211,31,254,31,254,31,78,31,53,31,37,31,53,31,53,30,241,31,177,31,80,31,54,31,54,30,95,31,66,31,58,31,106,31,106,30,105,31,209,31,187,31,187,30,13,31,41,31,41,30,166,31,35,31,59,31,84,31,112,31,85,31,194,31,7,31,73,31,58,31,58,30,58,29,127,31,127,30,191,31,191,30,224,31,34,31,55,31,55,30,220,31,246,31,243,31,243,30,60,31,29,31,159,31,159,30,181,31,111,31,1,31,195,31,29,31,164,31,175,31,129,31,11,31,11,30,172,31,200,31,94,31,37,31,112,31,180,31,175,31,200,31,214,31,214,30,214,29,214,28,214,27,214,26,214,25,30,31,30,30,153,31,253,31,42,31,79,31,127,31,124,31,124,30,58,31,13,31,120,31,60,31,187,31,187,30,187,29,60,31,156,31,185,31,8,31,123,31,238,31,246,31,159,31,123,31,48,31,154,31,154,30,154,29,231,31,235,31,123,31,6,31,6,30,74,31,57,31,93,31,93,30,134,31,19,31,19,30,58,31,58,30,128,31,251,31,251,30,214,31,130,31,169,31,233,31,162,31,64,31,66,31,133,31,18,31,18,30,217,31,61,31,41,31,227,31,152,31,93,31,93,31,93,30,172,31,68,31,68,30,69,31,142,31,142,30,248,31,130,31,181,31,244,31,244,30,224,31,181,31,72,31,72,30,156,31,114,31,114,30,57,31,151,31,234,31,149,31,149,30,129,31,29,31,185,31,153,31,46,31,82,31,179,31,100,31,161,31,231,31,221,31,211,31,1,31,153,31,153,30,156,31,22,31,123,31,168,31,166,31,166,30,166,29,206,31,116,31,51,31,51,30,139,31,167,31,167,30,239,31,117,31,117,30,189,31,90,31,163,31,167,31,94,31,236,31,236,31,223,31,150,31,25,31,238,31,177,31,70,31,70,30,196,31,176,31,187,31,216,31,184,31,8,31,8,30,48,31,104,31,10,31,10,30,229,31,239,31,115,31,115,30,140,31,229,31,116,31,116,30,56,31,243,31,59,31,234,31,130,31,130,30,217,31,207,31,94,31,94,30,94,29,82,31,115,31,245,31,245,31,245,30,245,29,91,31,7,31,28,31,28,30,28,29,99,31,189,31,189,30,159,31,67,31,144,31,107,31,46,31,66,31,165,31,241,31,241,30,48,31,197,31,160,31,155,31,168,31,168,30,160,31,234,31,100,31,99,31,50,31,172,31,223,31,221,31,211,31,196,31,45,31,118,31,25,31,128,31,176,31,203,31,74,31,255,31,106,31,106,30,64,31,187,31,68,31,163,31,186,31,32,31,24,31,84,31,115,31,241,31,71,31,136,31,171,31,79,31,79,30,142,31,100,31,100,30,132,31,132,30,187,31,105,31,175,31,255,31,255,30,255,29,179,31,122,31,247,31,247,30,247,29,14,31,14,30,14,29,136,31,48,31,25,31,177,31,177,30,177,29,171,31,62,31,50,31,50,30,50,29,50,28,129,31,36,31,36,30,36,29,165,31,253,31,145,31,145,30,153,31,95,31,11,31,33,31,123,31,204,31,231,31,207,31,206,31,38,31,112,31,45,31,128,31,160,31,160,30,24,31,123,31,38,31,141,31,182,31,162,31,5,31,203,31,220,31,76,31,170,31,28,31,129,31,67,31,151,31,61,31,110,31,79,31,39,31,154,31,104,31,104,30,104,31,30,31,144,31,99,31,99,30,166,31,166,30,166,29,123,31,163,31,60,31,16,31,136,31,180,31,152,31,152,30,117,31,111,31,232,31,152,31,21,31,208,31,109,31,109,30,134,31,40,31,255,31,242,31,209,31,211,31,1,31,201,31,130,31,67,31,67,30,70,31,51,31,140,31,62,31,5,31,211,31,34,31,192,31,217,31,68,31,185,31,13,31,13,30,100,31,100,30,16,31,103,31,135,31,135,30,10,31,234,31,120,31,150,31,69,31,123,31,124,31,217,31,40,31,65,31,94,31,127,31,198,31,176,31,250,31,250,30,165,31,137,31,1,31,14,31,251,31,188,31,214,31,123,31,55,31,194,31,147,31,217,31,241,31,144,31,144,30,238,31,216,31,112,31,48,31,132,31,224,31,78,31,198,31,138,31,87,31,224,31,133,31,56,31,5,31,45,31,225,31,253,31,126,31,111,31,105,31,31,31,31,30,31,29,108,31,108,30,116,31,116,30,49,31,235,31,142,31,69,31,146,31,146,30,166,31,169,31,205,31,205,30,221,31,221,30,203,31,220,31,182,31,176,31,68,31,82,31,91,31,194,31,53,31,17,31,12,31,171,31,89,31,202,31,202,30,41,31,178,31,178,30,3,31,51,31,253,31,253,30,97,31,106,31,240,31,207,31,66,31,222,31,9,31,7,31,199,31,199,30,71,31,218,31,161,31,193,31,171,31,147,31,147,30,25,31,89,31,186,31,45,31,78,31,188,31,239,31,140,31,140,30,207,31,202,31,244,31,31,31,76,31,206,31,166,31,248,31,248,30,204,31,160,31,250,31,209,31,96,31,105,31,180,31,185,31,234,31,95,31,216,31,216,30,194,31,118,31,99,31,143,31,133,31,133,30,172,31,218,31,141,31,239,31,198,31,198,30,166,31,7,31,111,31,111,30,240,31,26,31,32,31,203,31,106,31,106,30,119,31,119,30,178,31,105,31,105,30,248,31,205,31,27,31,194,31,10,31,126,31,50,31,133,31,249,31,249,30,63,31,63,30,175,31,11,31,134,31,30,31,93,31,195,31,195,30,159,31,220,31,95,31,83,31,73,31,7,31,131,31,1,31,106,31,226,31,253,31,253,30,118,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
