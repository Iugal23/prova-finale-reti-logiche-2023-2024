-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 851;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (124,0,227,0,125,0,202,0,0,0,0,0,86,0,21,0,0,0,164,0,194,0,184,0,10,0,125,0,212,0,96,0,62,0,209,0,223,0,254,0,0,0,56,0,19,0,144,0,209,0,58,0,0,0,76,0,253,0,134,0,220,0,183,0,63,0,54,0,0,0,108,0,66,0,21,0,148,0,3,0,162,0,233,0,86,0,0,0,209,0,0,0,52,0,240,0,227,0,184,0,103,0,68,0,45,0,0,0,0,0,21,0,194,0,95,0,141,0,30,0,151,0,228,0,92,0,168,0,53,0,130,0,54,0,236,0,12,0,27,0,161,0,1,0,120,0,39,0,240,0,0,0,0,0,0,0,42,0,145,0,68,0,104,0,187,0,0,0,214,0,242,0,152,0,0,0,0,0,0,0,45,0,0,0,0,0,92,0,0,0,226,0,97,0,120,0,235,0,223,0,52,0,0,0,131,0,0,0,0,0,51,0,201,0,65,0,216,0,140,0,60,0,0,0,0,0,149,0,142,0,53,0,55,0,194,0,0,0,131,0,0,0,182,0,0,0,174,0,69,0,201,0,141,0,16,0,0,0,229,0,240,0,198,0,249,0,46,0,0,0,179,0,121,0,4,0,0,0,156,0,223,0,189,0,3,0,133,0,207,0,163,0,221,0,157,0,216,0,152,0,162,0,0,0,0,0,209,0,212,0,245,0,230,0,187,0,190,0,125,0,224,0,167,0,0,0,108,0,9,0,50,0,0,0,188,0,0,0,37,0,202,0,0,0,0,0,0,0,0,0,0,0,175,0,0,0,3,0,238,0,63,0,140,0,0,0,120,0,29,0,0,0,156,0,177,0,238,0,99,0,70,0,0,0,14,0,191,0,0,0,248,0,234,0,227,0,174,0,72,0,0,0,242,0,51,0,59,0,143,0,203,0,62,0,0,0,0,0,177,0,80,0,0,0,137,0,73,0,170,0,118,0,12,0,30,0,0,0,246,0,0,0,50,0,34,0,26,0,106,0,73,0,21,0,104,0,0,0,0,0,117,0,238,0,0,0,122,0,0,0,0,0,0,0,85,0,189,0,116,0,160,0,0,0,102,0,14,0,78,0,4,0,0,0,0,0,169,0,218,0,137,0,34,0,249,0,156,0,170,0,252,0,98,0,68,0,67,0,134,0,0,0,106,0,213,0,0,0,151,0,0,0,0,0,101,0,0,0,0,0,170,0,130,0,20,0,0,0,0,0,150,0,211,0,216,0,115,0,74,0,219,0,0,0,0,0,135,0,161,0,209,0,138,0,44,0,176,0,138,0,0,0,66,0,26,0,19,0,0,0,41,0,69,0,141,0,58,0,208,0,0,0,81,0,33,0,0,0,240,0,9,0,52,0,226,0,64,0,253,0,73,0,93,0,194,0,0,0,65,0,167,0,0,0,90,0,184,0,30,0,164,0,210,0,0,0,229,0,59,0,51,0,0,0,0,0,208,0,0,0,208,0,18,0,34,0,151,0,251,0,0,0,232,0,0,0,0,0,76,0,247,0,219,0,198,0,234,0,0,0,0,0,0,0,0,0,28,0,218,0,119,0,125,0,90,0,182,0,0,0,59,0,63,0,14,0,107,0,186,0,221,0,238,0,175,0,0,0,0,0,11,0,194,0,150,0,158,0,87,0,42,0,11,0,139,0,204,0,227,0,97,0,221,0,69,0,0,0,148,0,52,0,169,0,40,0,255,0,0,0,115,0,48,0,0,0,177,0,65,0,251,0,70,0,0,0,180,0,201,0,0,0,239,0,164,0,220,0,54,0,213,0,243,0,141,0,0,0,0,0,220,0,0,0,17,0,0,0,0,0,0,0,214,0,166,0,229,0,237,0,150,0,156,0,171,0,33,0,162,0,158,0,201,0,0,0,68,0,0,0,211,0,16,0,134,0,0,0,19,0,174,0,167,0,110,0,0,0,30,0,189,0,202,0,114,0,221,0,119,0,0,0,57,0,125,0,113,0,241,0,219,0,13,0,43,0,0,0,0,0,110,0,170,0,125,0,10,0,103,0,53,0,192,0,222,0,188,0,0,0,93,0,0,0,221,0,109,0,35,0,73,0,184,0,110,0,255,0,152,0,0,0,83,0,198,0,164,0,59,0,21,0,2,0,0,0,195,0,0,0,35,0,163,0,103,0,223,0,71,0,102,0,104,0,219,0,182,0,67,0,180,0,38,0,38,0,5,0,7,0,209,0,135,0,147,0,16,0,35,0,0,0,182,0,55,0,0,0,107,0,4,0,159,0,141,0,243,0,0,0,0,0,161,0,122,0,153,0,182,0,0,0,113,0,11,0,158,0,228,0,162,0,17,0,247,0,58,0,199,0,213,0,75,0,125,0,221,0,119,0,164,0,22,0,220,0,162,0,203,0,29,0,17,0,46,0,5,0,104,0,236,0,137,0,24,0,155,0,247,0,172,0,249,0,116,0,214,0,23,0,148,0,196,0,94,0,228,0,212,0,124,0,149,0,0,0,62,0,0,0,0,0,0,0,42,0,66,0,132,0,180,0,226,0,0,0,8,0,152,0,31,0,191,0,223,0,14,0,222,0,0,0,79,0,1,0,105,0,0,0,38,0,249,0,235,0,10,0,98,0,68,0,224,0,111,0,19,0,0,0,67,0,0,0,35,0,210,0,0,0,123,0,74,0,0,0,157,0,86,0,141,0,108,0,107,0,171,0,89,0,43,0,85,0,113,0,168,0,244,0,175,0,240,0,237,0,188,0,0,0,19,0,55,0,21,0,147,0,207,0,22,0,4,0,0,0,0,0,53,0,24,0,88,0,110,0,0,0,117,0,0,0,56,0,0,0,9,0,80,0,0,0,136,0,179,0,0,0,0,0,126,0,0,0,0,0,246,0,67,0,167,0,153,0,0,0,187,0,34,0,84,0,4,0,231,0,40,0,77,0,127,0,57,0,156,0,71,0,240,0,158,0,7,0,164,0,49,0,45,0,78,0,50,0,225,0,0,0,51,0,186,0,54,0,220,0,0,0,20,0,156,0,0,0,94,0,231,0,65,0,195,0,42,0,36,0,93,0,134,0,74,0,37,0,0,0,227,0,10,0,180,0,142,0,207,0,0,0,59,0,245,0,15,0,99,0,78,0,32,0,187,0,0,0,224,0,0,0,0,0,0,0,0,0,203,0,0,0,64,0,77,0,130,0,85,0,39,0,103,0,36,0,132,0,123,0,179,0,0,0,104,0,143,0,52,0,18,0,152,0,127,0,238,0,0,0,201,0,0,0,247,0,139,0,226,0,138,0,43,0,119,0,234,0,96,0,0,0,0,0,242,0,215,0,92,0,63,0,240,0,93,0,135,0,0,0,115,0,102,0,73,0,197,0,131,0,136,0,205,0,250,0,244,0,167,0,152,0,198,0,160,0,0,0,52,0,248,0,133,0,141,0,0,0,203,0,228,0,19,0,0,0,90,0,144,0,224,0,46,0,0,0,134,0,104,0,54,0,56,0,212,0,0,0,181,0,84,0,143,0,112,0,95,0,75,0,176,0,209,0,171,0,0,0,4,0,40,0,102,0,188,0,78,0,0,0,99,0,22,0,40,0,0,0,251,0,22,0,229,0,21,0,13,0,57,0,39,0,0,0,166,0,149,0,0,0,154,0,202,0,0,0,0,0,43,0,103,0,0,0,148,0,219,0,169,0,27,0,31,0,0,0,16,0,0,0,181,0,0,0,100,0,29,0,233,0,247,0,65,0,134,0,141,0,159,0,200,0,0,0,0,0,190,0,0,0,45,0,190,0,201,0,233,0,241,0,194,0,159,0,94,0);
signal scenario_full  : scenario_type := (124,31,227,31,125,31,202,31,202,30,202,29,86,31,21,31,21,30,164,31,194,31,184,31,10,31,125,31,212,31,96,31,62,31,209,31,223,31,254,31,254,30,56,31,19,31,144,31,209,31,58,31,58,30,76,31,253,31,134,31,220,31,183,31,63,31,54,31,54,30,108,31,66,31,21,31,148,31,3,31,162,31,233,31,86,31,86,30,209,31,209,30,52,31,240,31,227,31,184,31,103,31,68,31,45,31,45,30,45,29,21,31,194,31,95,31,141,31,30,31,151,31,228,31,92,31,168,31,53,31,130,31,54,31,236,31,12,31,27,31,161,31,1,31,120,31,39,31,240,31,240,30,240,29,240,28,42,31,145,31,68,31,104,31,187,31,187,30,214,31,242,31,152,31,152,30,152,29,152,28,45,31,45,30,45,29,92,31,92,30,226,31,97,31,120,31,235,31,223,31,52,31,52,30,131,31,131,30,131,29,51,31,201,31,65,31,216,31,140,31,60,31,60,30,60,29,149,31,142,31,53,31,55,31,194,31,194,30,131,31,131,30,182,31,182,30,174,31,69,31,201,31,141,31,16,31,16,30,229,31,240,31,198,31,249,31,46,31,46,30,179,31,121,31,4,31,4,30,156,31,223,31,189,31,3,31,133,31,207,31,163,31,221,31,157,31,216,31,152,31,162,31,162,30,162,29,209,31,212,31,245,31,230,31,187,31,190,31,125,31,224,31,167,31,167,30,108,31,9,31,50,31,50,30,188,31,188,30,37,31,202,31,202,30,202,29,202,28,202,27,202,26,175,31,175,30,3,31,238,31,63,31,140,31,140,30,120,31,29,31,29,30,156,31,177,31,238,31,99,31,70,31,70,30,14,31,191,31,191,30,248,31,234,31,227,31,174,31,72,31,72,30,242,31,51,31,59,31,143,31,203,31,62,31,62,30,62,29,177,31,80,31,80,30,137,31,73,31,170,31,118,31,12,31,30,31,30,30,246,31,246,30,50,31,34,31,26,31,106,31,73,31,21,31,104,31,104,30,104,29,117,31,238,31,238,30,122,31,122,30,122,29,122,28,85,31,189,31,116,31,160,31,160,30,102,31,14,31,78,31,4,31,4,30,4,29,169,31,218,31,137,31,34,31,249,31,156,31,170,31,252,31,98,31,68,31,67,31,134,31,134,30,106,31,213,31,213,30,151,31,151,30,151,29,101,31,101,30,101,29,170,31,130,31,20,31,20,30,20,29,150,31,211,31,216,31,115,31,74,31,219,31,219,30,219,29,135,31,161,31,209,31,138,31,44,31,176,31,138,31,138,30,66,31,26,31,19,31,19,30,41,31,69,31,141,31,58,31,208,31,208,30,81,31,33,31,33,30,240,31,9,31,52,31,226,31,64,31,253,31,73,31,93,31,194,31,194,30,65,31,167,31,167,30,90,31,184,31,30,31,164,31,210,31,210,30,229,31,59,31,51,31,51,30,51,29,208,31,208,30,208,31,18,31,34,31,151,31,251,31,251,30,232,31,232,30,232,29,76,31,247,31,219,31,198,31,234,31,234,30,234,29,234,28,234,27,28,31,218,31,119,31,125,31,90,31,182,31,182,30,59,31,63,31,14,31,107,31,186,31,221,31,238,31,175,31,175,30,175,29,11,31,194,31,150,31,158,31,87,31,42,31,11,31,139,31,204,31,227,31,97,31,221,31,69,31,69,30,148,31,52,31,169,31,40,31,255,31,255,30,115,31,48,31,48,30,177,31,65,31,251,31,70,31,70,30,180,31,201,31,201,30,239,31,164,31,220,31,54,31,213,31,243,31,141,31,141,30,141,29,220,31,220,30,17,31,17,30,17,29,17,28,214,31,166,31,229,31,237,31,150,31,156,31,171,31,33,31,162,31,158,31,201,31,201,30,68,31,68,30,211,31,16,31,134,31,134,30,19,31,174,31,167,31,110,31,110,30,30,31,189,31,202,31,114,31,221,31,119,31,119,30,57,31,125,31,113,31,241,31,219,31,13,31,43,31,43,30,43,29,110,31,170,31,125,31,10,31,103,31,53,31,192,31,222,31,188,31,188,30,93,31,93,30,221,31,109,31,35,31,73,31,184,31,110,31,255,31,152,31,152,30,83,31,198,31,164,31,59,31,21,31,2,31,2,30,195,31,195,30,35,31,163,31,103,31,223,31,71,31,102,31,104,31,219,31,182,31,67,31,180,31,38,31,38,31,5,31,7,31,209,31,135,31,147,31,16,31,35,31,35,30,182,31,55,31,55,30,107,31,4,31,159,31,141,31,243,31,243,30,243,29,161,31,122,31,153,31,182,31,182,30,113,31,11,31,158,31,228,31,162,31,17,31,247,31,58,31,199,31,213,31,75,31,125,31,221,31,119,31,164,31,22,31,220,31,162,31,203,31,29,31,17,31,46,31,5,31,104,31,236,31,137,31,24,31,155,31,247,31,172,31,249,31,116,31,214,31,23,31,148,31,196,31,94,31,228,31,212,31,124,31,149,31,149,30,62,31,62,30,62,29,62,28,42,31,66,31,132,31,180,31,226,31,226,30,8,31,152,31,31,31,191,31,223,31,14,31,222,31,222,30,79,31,1,31,105,31,105,30,38,31,249,31,235,31,10,31,98,31,68,31,224,31,111,31,19,31,19,30,67,31,67,30,35,31,210,31,210,30,123,31,74,31,74,30,157,31,86,31,141,31,108,31,107,31,171,31,89,31,43,31,85,31,113,31,168,31,244,31,175,31,240,31,237,31,188,31,188,30,19,31,55,31,21,31,147,31,207,31,22,31,4,31,4,30,4,29,53,31,24,31,88,31,110,31,110,30,117,31,117,30,56,31,56,30,9,31,80,31,80,30,136,31,179,31,179,30,179,29,126,31,126,30,126,29,246,31,67,31,167,31,153,31,153,30,187,31,34,31,84,31,4,31,231,31,40,31,77,31,127,31,57,31,156,31,71,31,240,31,158,31,7,31,164,31,49,31,45,31,78,31,50,31,225,31,225,30,51,31,186,31,54,31,220,31,220,30,20,31,156,31,156,30,94,31,231,31,65,31,195,31,42,31,36,31,93,31,134,31,74,31,37,31,37,30,227,31,10,31,180,31,142,31,207,31,207,30,59,31,245,31,15,31,99,31,78,31,32,31,187,31,187,30,224,31,224,30,224,29,224,28,224,27,203,31,203,30,64,31,77,31,130,31,85,31,39,31,103,31,36,31,132,31,123,31,179,31,179,30,104,31,143,31,52,31,18,31,152,31,127,31,238,31,238,30,201,31,201,30,247,31,139,31,226,31,138,31,43,31,119,31,234,31,96,31,96,30,96,29,242,31,215,31,92,31,63,31,240,31,93,31,135,31,135,30,115,31,102,31,73,31,197,31,131,31,136,31,205,31,250,31,244,31,167,31,152,31,198,31,160,31,160,30,52,31,248,31,133,31,141,31,141,30,203,31,228,31,19,31,19,30,90,31,144,31,224,31,46,31,46,30,134,31,104,31,54,31,56,31,212,31,212,30,181,31,84,31,143,31,112,31,95,31,75,31,176,31,209,31,171,31,171,30,4,31,40,31,102,31,188,31,78,31,78,30,99,31,22,31,40,31,40,30,251,31,22,31,229,31,21,31,13,31,57,31,39,31,39,30,166,31,149,31,149,30,154,31,202,31,202,30,202,29,43,31,103,31,103,30,148,31,219,31,169,31,27,31,31,31,31,30,16,31,16,30,181,31,181,30,100,31,29,31,233,31,247,31,65,31,134,31,141,31,159,31,200,31,200,30,200,29,190,31,190,30,45,31,190,31,201,31,233,31,241,31,194,31,159,31,94,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
