-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1003;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (218,0,81,0,83,0,0,0,223,0,250,0,21,0,116,0,106,0,53,0,136,0,2,0,143,0,15,0,31,0,0,0,0,0,158,0,0,0,164,0,0,0,143,0,31,0,0,0,226,0,84,0,0,0,6,0,141,0,0,0,36,0,198,0,0,0,104,0,198,0,170,0,42,0,0,0,218,0,167,0,207,0,132,0,141,0,152,0,152,0,0,0,37,0,7,0,230,0,122,0,89,0,188,0,125,0,156,0,0,0,0,0,2,0,219,0,234,0,191,0,217,0,225,0,104,0,140,0,0,0,67,0,195,0,140,0,177,0,0,0,45,0,0,0,224,0,0,0,0,0,155,0,132,0,144,0,0,0,159,0,96,0,148,0,208,0,180,0,152,0,0,0,227,0,142,0,151,0,22,0,15,0,220,0,126,0,0,0,0,0,170,0,189,0,176,0,202,0,100,0,20,0,237,0,97,0,41,0,167,0,41,0,164,0,145,0,222,0,255,0,64,0,84,0,0,0,150,0,70,0,142,0,31,0,154,0,254,0,149,0,54,0,42,0,0,0,149,0,0,0,167,0,158,0,112,0,0,0,0,0,175,0,223,0,102,0,0,0,255,0,13,0,171,0,170,0,131,0,172,0,250,0,192,0,228,0,218,0,0,0,69,0,17,0,61,0,75,0,212,0,243,0,47,0,189,0,3,0,212,0,186,0,111,0,51,0,62,0,214,0,62,0,204,0,143,0,27,0,0,0,22,0,0,0,210,0,214,0,149,0,8,0,5,0,34,0,23,0,0,0,35,0,0,0,0,0,243,0,0,0,88,0,242,0,242,0,124,0,167,0,100,0,0,0,130,0,253,0,0,0,56,0,0,0,180,0,0,0,181,0,0,0,50,0,140,0,0,0,239,0,0,0,0,0,240,0,82,0,160,0,222,0,93,0,17,0,108,0,0,0,194,0,223,0,123,0,206,0,51,0,0,0,76,0,145,0,113,0,165,0,242,0,110,0,0,0,241,0,178,0,28,0,247,0,176,0,154,0,39,0,42,0,5,0,7,0,191,0,14,0,0,0,0,0,0,0,66,0,62,0,31,0,168,0,40,0,77,0,45,0,179,0,179,0,0,0,180,0,226,0,113,0,0,0,201,0,157,0,0,0,144,0,166,0,180,0,0,0,69,0,64,0,105,0,0,0,194,0,150,0,164,0,60,0,0,0,172,0,109,0,189,0,121,0,202,0,0,0,146,0,22,0,16,0,119,0,92,0,0,0,187,0,185,0,131,0,254,0,112,0,182,0,209,0,176,0,223,0,254,0,23,0,193,0,125,0,5,0,84,0,123,0,48,0,0,0,22,0,34,0,85,0,0,0,95,0,163,0,166,0,247,0,183,0,99,0,213,0,12,0,44,0,123,0,231,0,63,0,35,0,28,0,232,0,99,0,29,0,5,0,0,0,0,0,46,0,21,0,228,0,170,0,74,0,0,0,255,0,232,0,78,0,152,0,130,0,121,0,129,0,0,0,87,0,181,0,0,0,88,0,162,0,0,0,239,0,57,0,53,0,34,0,59,0,109,0,22,0,97,0,85,0,228,0,113,0,0,0,84,0,0,0,0,0,188,0,70,0,107,0,201,0,83,0,41,0,0,0,23,0,56,0,218,0,187,0,206,0,0,0,187,0,0,0,201,0,0,0,254,0,156,0,1,0,0,0,198,0,100,0,117,0,59,0,164,0,37,0,114,0,255,0,194,0,6,0,0,0,185,0,0,0,114,0,204,0,0,0,90,0,78,0,217,0,100,0,0,0,0,0,121,0,47,0,175,0,193,0,0,0,127,0,0,0,192,0,65,0,87,0,116,0,0,0,33,0,0,0,43,0,15,0,45,0,238,0,205,0,73,0,245,0,0,0,9,0,28,0,244,0,36,0,208,0,0,0,56,0,0,0,0,0,90,0,60,0,53,0,88,0,149,0,45,0,165,0,94,0,0,0,238,0,13,0,1,0,121,0,66,0,149,0,55,0,26,0,0,0,102,0,131,0,96,0,26,0,80,0,130,0,228,0,52,0,238,0,191,0,108,0,0,0,0,0,193,0,88,0,0,0,99,0,148,0,0,0,192,0,76,0,145,0,186,0,161,0,0,0,52,0,197,0,183,0,68,0,33,0,15,0,25,0,55,0,0,0,184,0,213,0,0,0,139,0,151,0,160,0,233,0,229,0,200,0,8,0,172,0,63,0,0,0,224,0,0,0,29,0,0,0,47,0,0,0,129,0,53,0,122,0,210,0,169,0,146,0,83,0,113,0,0,0,5,0,187,0,47,0,0,0,169,0,33,0,183,0,228,0,218,0,248,0,168,0,194,0,92,0,0,0,212,0,0,0,6,0,0,0,153,0,246,0,0,0,79,0,187,0,0,0,30,0,131,0,50,0,46,0,161,0,0,0,179,0,252,0,50,0,117,0,121,0,0,0,0,0,39,0,48,0,36,0,0,0,0,0,60,0,0,0,181,0,83,0,108,0,221,0,50,0,42,0,74,0,57,0,0,0,0,0,0,0,185,0,154,0,84,0,155,0,95,0,66,0,0,0,69,0,219,0,249,0,19,0,0,0,140,0,29,0,58,0,197,0,40,0,121,0,185,0,141,0,0,0,0,0,56,0,0,0,45,0,12,0,84,0,253,0,54,0,91,0,160,0,160,0,35,0,254,0,118,0,56,0,211,0,0,0,43,0,117,0,16,0,34,0,164,0,123,0,0,0,0,0,210,0,9,0,193,0,0,0,0,0,0,0,101,0,13,0,23,0,32,0,119,0,90,0,149,0,22,0,43,0,0,0,136,0,86,0,0,0,3,0,210,0,4,0,60,0,0,0,192,0,0,0,56,0,6,0,113,0,0,0,121,0,0,0,0,0,57,0,0,0,197,0,64,0,81,0,103,0,160,0,140,0,0,0,107,0,4,0,212,0,237,0,103,0,200,0,80,0,203,0,118,0,161,0,49,0,0,0,246,0,52,0,31,0,101,0,81,0,118,0,0,0,28,0,99,0,0,0,189,0,31,0,0,0,229,0,55,0,47,0,188,0,12,0,231,0,97,0,153,0,110,0,0,0,167,0,206,0,120,0,191,0,81,0,0,0,32,0,0,0,2,0,63,0,0,0,5,0,153,0,118,0,0,0,126,0,0,0,217,0,0,0,137,0,6,0,231,0,52,0,0,0,0,0,68,0,181,0,32,0,216,0,0,0,0,0,161,0,77,0,238,0,118,0,60,0,118,0,79,0,0,0,76,0,151,0,6,0,68,0,63,0,229,0,182,0,232,0,151,0,50,0,164,0,243,0,52,0,0,0,0,0,246,0,183,0,206,0,252,0,39,0,111,0,0,0,99,0,210,0,57,0,22,0,143,0,78,0,103,0,128,0,212,0,239,0,214,0,40,0,16,0,217,0,121,0,220,0,0,0,0,0,96,0,138,0,0,0,55,0,158,0,121,0,0,0,209,0,106,0,215,0,176,0,32,0,134,0,115,0,71,0,203,0,38,0,58,0,177,0,70,0,12,0,231,0,151,0,0,0,152,0,154,0,161,0,220,0,0,0,196,0,18,0,150,0,188,0,188,0,204,0,95,0,74,0,0,0,166,0,115,0,127,0,69,0,229,0,210,0,0,0,221,0,8,0,143,0,0,0,227,0,220,0,0,0,253,0,255,0,197,0,65,0,88,0,0,0,14,0,0,0,0,0,253,0,173,0,0,0,251,0,0,0,182,0,7,0,33,0,77,0,97,0,177,0,0,0,245,0,45,0,0,0,178,0,140,0,87,0,147,0,85,0,0,0,186,0,0,0,206,0,0,0,0,0,222,0,34,0,192,0,65,0,0,0,24,0,114,0,73,0,33,0,226,0,207,0,34,0,0,0,52,0,14,0,216,0,214,0,212,0,193,0,157,0,202,0,154,0,73,0,117,0,147,0,105,0,193,0,233,0,232,0,208,0,141,0,0,0,95,0,182,0,215,0,0,0,232,0,49,0,22,0,185,0,164,0,0,0,173,0,143,0,65,0,58,0,138,0,0,0,5,0,251,0,67,0,179,0,81,0,20,0,78,0,0,0,0,0,131,0,0,0,206,0,116,0,186,0,47,0,77,0,0,0,40,0,26,0,214,0,94,0,82,0,89,0,148,0,83,0,59,0,138,0,67,0,1,0,0,0,0,0,0,0,129,0,166,0,0,0,100,0,133,0,0,0,181,0,88,0,131,0,56,0,39,0,244,0,223,0,1,0,19,0,79,0,157,0,204,0,0,0,206,0,166,0,0,0,236,0,19,0,0,0,0,0,98,0,201,0,98,0,63,0,239,0,0,0,0,0,88,0,199,0,53,0,103,0,150,0,34,0,86,0,105,0,198,0,228,0,0,0,25,0,65,0,0,0,223,0,255,0,0,0,51,0,0,0,205,0,0,0,91,0,160,0,44,0,0,0,7,0,2,0,54,0,30,0,255,0,0,0,4,0,74,0,69,0,250,0);
signal scenario_full  : scenario_type := (218,31,81,31,83,31,83,30,223,31,250,31,21,31,116,31,106,31,53,31,136,31,2,31,143,31,15,31,31,31,31,30,31,29,158,31,158,30,164,31,164,30,143,31,31,31,31,30,226,31,84,31,84,30,6,31,141,31,141,30,36,31,198,31,198,30,104,31,198,31,170,31,42,31,42,30,218,31,167,31,207,31,132,31,141,31,152,31,152,31,152,30,37,31,7,31,230,31,122,31,89,31,188,31,125,31,156,31,156,30,156,29,2,31,219,31,234,31,191,31,217,31,225,31,104,31,140,31,140,30,67,31,195,31,140,31,177,31,177,30,45,31,45,30,224,31,224,30,224,29,155,31,132,31,144,31,144,30,159,31,96,31,148,31,208,31,180,31,152,31,152,30,227,31,142,31,151,31,22,31,15,31,220,31,126,31,126,30,126,29,170,31,189,31,176,31,202,31,100,31,20,31,237,31,97,31,41,31,167,31,41,31,164,31,145,31,222,31,255,31,64,31,84,31,84,30,150,31,70,31,142,31,31,31,154,31,254,31,149,31,54,31,42,31,42,30,149,31,149,30,167,31,158,31,112,31,112,30,112,29,175,31,223,31,102,31,102,30,255,31,13,31,171,31,170,31,131,31,172,31,250,31,192,31,228,31,218,31,218,30,69,31,17,31,61,31,75,31,212,31,243,31,47,31,189,31,3,31,212,31,186,31,111,31,51,31,62,31,214,31,62,31,204,31,143,31,27,31,27,30,22,31,22,30,210,31,214,31,149,31,8,31,5,31,34,31,23,31,23,30,35,31,35,30,35,29,243,31,243,30,88,31,242,31,242,31,124,31,167,31,100,31,100,30,130,31,253,31,253,30,56,31,56,30,180,31,180,30,181,31,181,30,50,31,140,31,140,30,239,31,239,30,239,29,240,31,82,31,160,31,222,31,93,31,17,31,108,31,108,30,194,31,223,31,123,31,206,31,51,31,51,30,76,31,145,31,113,31,165,31,242,31,110,31,110,30,241,31,178,31,28,31,247,31,176,31,154,31,39,31,42,31,5,31,7,31,191,31,14,31,14,30,14,29,14,28,66,31,62,31,31,31,168,31,40,31,77,31,45,31,179,31,179,31,179,30,180,31,226,31,113,31,113,30,201,31,157,31,157,30,144,31,166,31,180,31,180,30,69,31,64,31,105,31,105,30,194,31,150,31,164,31,60,31,60,30,172,31,109,31,189,31,121,31,202,31,202,30,146,31,22,31,16,31,119,31,92,31,92,30,187,31,185,31,131,31,254,31,112,31,182,31,209,31,176,31,223,31,254,31,23,31,193,31,125,31,5,31,84,31,123,31,48,31,48,30,22,31,34,31,85,31,85,30,95,31,163,31,166,31,247,31,183,31,99,31,213,31,12,31,44,31,123,31,231,31,63,31,35,31,28,31,232,31,99,31,29,31,5,31,5,30,5,29,46,31,21,31,228,31,170,31,74,31,74,30,255,31,232,31,78,31,152,31,130,31,121,31,129,31,129,30,87,31,181,31,181,30,88,31,162,31,162,30,239,31,57,31,53,31,34,31,59,31,109,31,22,31,97,31,85,31,228,31,113,31,113,30,84,31,84,30,84,29,188,31,70,31,107,31,201,31,83,31,41,31,41,30,23,31,56,31,218,31,187,31,206,31,206,30,187,31,187,30,201,31,201,30,254,31,156,31,1,31,1,30,198,31,100,31,117,31,59,31,164,31,37,31,114,31,255,31,194,31,6,31,6,30,185,31,185,30,114,31,204,31,204,30,90,31,78,31,217,31,100,31,100,30,100,29,121,31,47,31,175,31,193,31,193,30,127,31,127,30,192,31,65,31,87,31,116,31,116,30,33,31,33,30,43,31,15,31,45,31,238,31,205,31,73,31,245,31,245,30,9,31,28,31,244,31,36,31,208,31,208,30,56,31,56,30,56,29,90,31,60,31,53,31,88,31,149,31,45,31,165,31,94,31,94,30,238,31,13,31,1,31,121,31,66,31,149,31,55,31,26,31,26,30,102,31,131,31,96,31,26,31,80,31,130,31,228,31,52,31,238,31,191,31,108,31,108,30,108,29,193,31,88,31,88,30,99,31,148,31,148,30,192,31,76,31,145,31,186,31,161,31,161,30,52,31,197,31,183,31,68,31,33,31,15,31,25,31,55,31,55,30,184,31,213,31,213,30,139,31,151,31,160,31,233,31,229,31,200,31,8,31,172,31,63,31,63,30,224,31,224,30,29,31,29,30,47,31,47,30,129,31,53,31,122,31,210,31,169,31,146,31,83,31,113,31,113,30,5,31,187,31,47,31,47,30,169,31,33,31,183,31,228,31,218,31,248,31,168,31,194,31,92,31,92,30,212,31,212,30,6,31,6,30,153,31,246,31,246,30,79,31,187,31,187,30,30,31,131,31,50,31,46,31,161,31,161,30,179,31,252,31,50,31,117,31,121,31,121,30,121,29,39,31,48,31,36,31,36,30,36,29,60,31,60,30,181,31,83,31,108,31,221,31,50,31,42,31,74,31,57,31,57,30,57,29,57,28,185,31,154,31,84,31,155,31,95,31,66,31,66,30,69,31,219,31,249,31,19,31,19,30,140,31,29,31,58,31,197,31,40,31,121,31,185,31,141,31,141,30,141,29,56,31,56,30,45,31,12,31,84,31,253,31,54,31,91,31,160,31,160,31,35,31,254,31,118,31,56,31,211,31,211,30,43,31,117,31,16,31,34,31,164,31,123,31,123,30,123,29,210,31,9,31,193,31,193,30,193,29,193,28,101,31,13,31,23,31,32,31,119,31,90,31,149,31,22,31,43,31,43,30,136,31,86,31,86,30,3,31,210,31,4,31,60,31,60,30,192,31,192,30,56,31,6,31,113,31,113,30,121,31,121,30,121,29,57,31,57,30,197,31,64,31,81,31,103,31,160,31,140,31,140,30,107,31,4,31,212,31,237,31,103,31,200,31,80,31,203,31,118,31,161,31,49,31,49,30,246,31,52,31,31,31,101,31,81,31,118,31,118,30,28,31,99,31,99,30,189,31,31,31,31,30,229,31,55,31,47,31,188,31,12,31,231,31,97,31,153,31,110,31,110,30,167,31,206,31,120,31,191,31,81,31,81,30,32,31,32,30,2,31,63,31,63,30,5,31,153,31,118,31,118,30,126,31,126,30,217,31,217,30,137,31,6,31,231,31,52,31,52,30,52,29,68,31,181,31,32,31,216,31,216,30,216,29,161,31,77,31,238,31,118,31,60,31,118,31,79,31,79,30,76,31,151,31,6,31,68,31,63,31,229,31,182,31,232,31,151,31,50,31,164,31,243,31,52,31,52,30,52,29,246,31,183,31,206,31,252,31,39,31,111,31,111,30,99,31,210,31,57,31,22,31,143,31,78,31,103,31,128,31,212,31,239,31,214,31,40,31,16,31,217,31,121,31,220,31,220,30,220,29,96,31,138,31,138,30,55,31,158,31,121,31,121,30,209,31,106,31,215,31,176,31,32,31,134,31,115,31,71,31,203,31,38,31,58,31,177,31,70,31,12,31,231,31,151,31,151,30,152,31,154,31,161,31,220,31,220,30,196,31,18,31,150,31,188,31,188,31,204,31,95,31,74,31,74,30,166,31,115,31,127,31,69,31,229,31,210,31,210,30,221,31,8,31,143,31,143,30,227,31,220,31,220,30,253,31,255,31,197,31,65,31,88,31,88,30,14,31,14,30,14,29,253,31,173,31,173,30,251,31,251,30,182,31,7,31,33,31,77,31,97,31,177,31,177,30,245,31,45,31,45,30,178,31,140,31,87,31,147,31,85,31,85,30,186,31,186,30,206,31,206,30,206,29,222,31,34,31,192,31,65,31,65,30,24,31,114,31,73,31,33,31,226,31,207,31,34,31,34,30,52,31,14,31,216,31,214,31,212,31,193,31,157,31,202,31,154,31,73,31,117,31,147,31,105,31,193,31,233,31,232,31,208,31,141,31,141,30,95,31,182,31,215,31,215,30,232,31,49,31,22,31,185,31,164,31,164,30,173,31,143,31,65,31,58,31,138,31,138,30,5,31,251,31,67,31,179,31,81,31,20,31,78,31,78,30,78,29,131,31,131,30,206,31,116,31,186,31,47,31,77,31,77,30,40,31,26,31,214,31,94,31,82,31,89,31,148,31,83,31,59,31,138,31,67,31,1,31,1,30,1,29,1,28,129,31,166,31,166,30,100,31,133,31,133,30,181,31,88,31,131,31,56,31,39,31,244,31,223,31,1,31,19,31,79,31,157,31,204,31,204,30,206,31,166,31,166,30,236,31,19,31,19,30,19,29,98,31,201,31,98,31,63,31,239,31,239,30,239,29,88,31,199,31,53,31,103,31,150,31,34,31,86,31,105,31,198,31,228,31,228,30,25,31,65,31,65,30,223,31,255,31,255,30,51,31,51,30,205,31,205,30,91,31,160,31,44,31,44,30,7,31,2,31,54,31,30,31,255,31,255,30,4,31,74,31,69,31,250,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
