-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 986;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (32,0,3,0,167,0,87,0,31,0,82,0,241,0,189,0,180,0,139,0,207,0,71,0,135,0,56,0,204,0,122,0,0,0,0,0,65,0,70,0,0,0,0,0,122,0,44,0,0,0,221,0,122,0,59,0,243,0,0,0,136,0,205,0,0,0,20,0,103,0,51,0,127,0,0,0,62,0,111,0,250,0,247,0,188,0,0,0,205,0,151,0,17,0,215,0,182,0,98,0,0,0,0,0,220,0,25,0,0,0,47,0,206,0,15,0,7,0,99,0,0,0,30,0,204,0,206,0,196,0,46,0,22,0,0,0,174,0,0,0,199,0,240,0,111,0,0,0,171,0,3,0,113,0,16,0,47,0,248,0,2,0,57,0,83,0,238,0,0,0,4,0,187,0,135,0,152,0,202,0,155,0,201,0,65,0,209,0,135,0,40,0,252,0,19,0,224,0,220,0,56,0,230,0,181,0,41,0,198,0,1,0,180,0,124,0,0,0,26,0,34,0,147,0,157,0,29,0,0,0,217,0,0,0,109,0,61,0,148,0,0,0,0,0,60,0,97,0,0,0,238,0,168,0,99,0,65,0,230,0,0,0,248,0,0,0,10,0,197,0,107,0,128,0,64,0,243,0,160,0,81,0,218,0,0,0,0,0,133,0,119,0,45,0,117,0,169,0,109,0,42,0,0,0,21,0,147,0,129,0,121,0,141,0,180,0,132,0,248,0,219,0,0,0,0,0,0,0,47,0,42,0,19,0,99,0,148,0,178,0,78,0,154,0,146,0,135,0,176,0,0,0,0,0,112,0,129,0,0,0,104,0,88,0,215,0,149,0,250,0,76,0,149,0,103,0,175,0,31,0,110,0,117,0,77,0,248,0,100,0,15,0,228,0,73,0,0,0,55,0,0,0,198,0,78,0,233,0,80,0,18,0,94,0,205,0,179,0,15,0,58,0,194,0,228,0,9,0,171,0,173,0,202,0,202,0,115,0,249,0,162,0,28,0,0,0,164,0,0,0,56,0,211,0,196,0,37,0,0,0,37,0,113,0,145,0,198,0,0,0,9,0,0,0,111,0,0,0,250,0,151,0,109,0,186,0,167,0,184,0,22,0,231,0,117,0,28,0,56,0,0,0,179,0,234,0,38,0,184,0,152,0,216,0,18,0,200,0,129,0,195,0,173,0,27,0,26,0,0,0,0,0,223,0,86,0,139,0,120,0,244,0,0,0,161,0,125,0,0,0,107,0,125,0,232,0,0,0,153,0,192,0,0,0,138,0,0,0,94,0,98,0,0,0,0,0,13,0,0,0,185,0,186,0,0,0,33,0,224,0,0,0,223,0,203,0,105,0,10,0,41,0,63,0,19,0,0,0,176,0,59,0,160,0,211,0,227,0,73,0,0,0,37,0,137,0,92,0,0,0,43,0,129,0,178,0,17,0,57,0,175,0,129,0,0,0,76,0,84,0,218,0,47,0,89,0,0,0,216,0,202,0,189,0,249,0,165,0,0,0,0,0,240,0,0,0,89,0,80,0,233,0,60,0,36,0,162,0,184,0,214,0,85,0,29,0,18,0,197,0,130,0,154,0,200,0,223,0,0,0,190,0,190,0,247,0,69,0,234,0,182,0,230,0,235,0,187,0,0,0,34,0,221,0,160,0,106,0,117,0,0,0,186,0,219,0,0,0,123,0,130,0,253,0,61,0,0,0,171,0,213,0,219,0,0,0,74,0,0,0,110,0,188,0,51,0,83,0,33,0,141,0,0,0,235,0,61,0,113,0,255,0,0,0,140,0,201,0,61,0,85,0,29,0,161,0,124,0,5,0,67,0,189,0,174,0,122,0,66,0,0,0,141,0,45,0,106,0,193,0,96,0,102,0,210,0,48,0,200,0,0,0,29,0,129,0,251,0,228,0,202,0,22,0,0,0,0,0,60,0,0,0,0,0,124,0,0,0,231,0,0,0,0,0,0,0,51,0,5,0,0,0,204,0,246,0,192,0,0,0,249,0,106,0,250,0,162,0,0,0,80,0,147,0,211,0,99,0,163,0,114,0,0,0,192,0,164,0,148,0,190,0,69,0,0,0,209,0,106,0,85,0,0,0,29,0,61,0,47,0,0,0,57,0,24,0,0,0,119,0,222,0,191,0,93,0,158,0,140,0,48,0,179,0,0,0,215,0,0,0,233,0,107,0,89,0,212,0,0,0,250,0,48,0,213,0,76,0,35,0,179,0,31,0,186,0,112,0,134,0,240,0,42,0,84,0,47,0,217,0,82,0,254,0,210,0,66,0,138,0,81,0,100,0,0,0,144,0,0,0,153,0,49,0,176,0,2,0,194,0,81,0,226,0,230,0,45,0,0,0,132,0,0,0,173,0,166,0,186,0,163,0,0,0,80,0,54,0,0,0,218,0,45,0,163,0,0,0,109,0,188,0,127,0,177,0,0,0,202,0,153,0,1,0,48,0,41,0,130,0,63,0,79,0,0,0,131,0,140,0,101,0,253,0,43,0,178,0,0,0,22,0,0,0,212,0,6,0,169,0,160,0,39,0,0,0,182,0,0,0,142,0,39,0,153,0,0,0,183,0,0,0,31,0,223,0,0,0,244,0,144,0,210,0,21,0,125,0,195,0,72,0,0,0,206,0,68,0,228,0,152,0,0,0,232,0,0,0,163,0,247,0,0,0,0,0,169,0,144,0,101,0,47,0,239,0,107,0,188,0,7,0,37,0,0,0,100,0,230,0,207,0,171,0,31,0,219,0,144,0,0,0,4,0,228,0,165,0,8,0,253,0,0,0,5,0,229,0,73,0,0,0,0,0,0,0,187,0,58,0,0,0,0,0,204,0,118,0,244,0,89,0,0,0,0,0,208,0,0,0,30,0,223,0,1,0,83,0,229,0,0,0,0,0,0,0,246,0,238,0,144,0,0,0,67,0,0,0,234,0,78,0,116,0,116,0,95,0,37,0,148,0,117,0,19,0,250,0,194,0,0,0,103,0,58,0,72,0,145,0,237,0,51,0,82,0,236,0,175,0,110,0,167,0,0,0,0,0,34,0,0,0,91,0,4,0,16,0,90,0,74,0,164,0,66,0,156,0,138,0,254,0,58,0,233,0,108,0,191,0,114,0,50,0,121,0,186,0,38,0,65,0,227,0,105,0,0,0,0,0,0,0,164,0,40,0,119,0,188,0,58,0,218,0,0,0,102,0,253,0,39,0,0,0,129,0,0,0,221,0,184,0,102,0,160,0,182,0,0,0,62,0,135,0,109,0,71,0,0,0,176,0,0,0,136,0,146,0,0,0,22,0,228,0,105,0,92,0,164,0,10,0,0,0,104,0,176,0,182,0,0,0,228,0,0,0,7,0,192,0,0,0,229,0,21,0,0,0,0,0,251,0,123,0,49,0,0,0,153,0,84,0,0,0,250,0,76,0,83,0,0,0,249,0,82,0,210,0,51,0,0,0,0,0,205,0,0,0,0,0,142,0,125,0,0,0,11,0,97,0,49,0,179,0,29,0,0,0,99,0,43,0,0,0,69,0,0,0,0,0,12,0,200,0,229,0,152,0,142,0,0,0,13,0,44,0,11,0,26,0,37,0,107,0,159,0,117,0,3,0,4,0,0,0,172,0,13,0,161,0,165,0,145,0,44,0,197,0,50,0,170,0,172,0,219,0,0,0,44,0,10,0,154,0,223,0,142,0,0,0,190,0,25,0,239,0,103,0,112,0,9,0,150,0,72,0,0,0,38,0,83,0,150,0,140,0,45,0,99,0,206,0,76,0,121,0,184,0,105,0,148,0,0,0,21,0,14,0,205,0,169,0,0,0,0,0,119,0,201,0,92,0,124,0,0,0,98,0,117,0,174,0,186,0,0,0,0,0,134,0,0,0,193,0,0,0,93,0,128,0,17,0,0,0,0,0,0,0,183,0,119,0,247,0,183,0,0,0,173,0,190,0,0,0,125,0,202,0,63,0,90,0,186,0,40,0,158,0,220,0,160,0,0,0,47,0,74,0,0,0,193,0,0,0,204,0,59,0,155,0,202,0,0,0,111,0,100,0,203,0,23,0,0,0,0,0,0,0,173,0,169,0,53,0,222,0,151,0,0,0,139,0,112,0,207,0,0,0,49,0,182,0,109,0,219,0,40,0,138,0,194,0,209,0,0,0,238,0,245,0,25,0,135,0,34,0,2,0,0,0,183,0,18,0,24,0,96,0,198,0,250,0,147,0,183,0,179,0,0,0,0,0,154,0,60,0,0,0,176,0,105,0,254,0,42,0,188,0,41,0,0,0,234,0,226,0,12,0,0,0,54,0,0,0,12,0,125,0,0,0,37,0,0,0,238,0,176,0,229,0,58,0,241,0,0,0,197,0,234,0,0,0,0,0,219,0,0,0,0,0,216,0,121,0,0,0,46,0,16,0,117,0);
signal scenario_full  : scenario_type := (32,31,3,31,167,31,87,31,31,31,82,31,241,31,189,31,180,31,139,31,207,31,71,31,135,31,56,31,204,31,122,31,122,30,122,29,65,31,70,31,70,30,70,29,122,31,44,31,44,30,221,31,122,31,59,31,243,31,243,30,136,31,205,31,205,30,20,31,103,31,51,31,127,31,127,30,62,31,111,31,250,31,247,31,188,31,188,30,205,31,151,31,17,31,215,31,182,31,98,31,98,30,98,29,220,31,25,31,25,30,47,31,206,31,15,31,7,31,99,31,99,30,30,31,204,31,206,31,196,31,46,31,22,31,22,30,174,31,174,30,199,31,240,31,111,31,111,30,171,31,3,31,113,31,16,31,47,31,248,31,2,31,57,31,83,31,238,31,238,30,4,31,187,31,135,31,152,31,202,31,155,31,201,31,65,31,209,31,135,31,40,31,252,31,19,31,224,31,220,31,56,31,230,31,181,31,41,31,198,31,1,31,180,31,124,31,124,30,26,31,34,31,147,31,157,31,29,31,29,30,217,31,217,30,109,31,61,31,148,31,148,30,148,29,60,31,97,31,97,30,238,31,168,31,99,31,65,31,230,31,230,30,248,31,248,30,10,31,197,31,107,31,128,31,64,31,243,31,160,31,81,31,218,31,218,30,218,29,133,31,119,31,45,31,117,31,169,31,109,31,42,31,42,30,21,31,147,31,129,31,121,31,141,31,180,31,132,31,248,31,219,31,219,30,219,29,219,28,47,31,42,31,19,31,99,31,148,31,178,31,78,31,154,31,146,31,135,31,176,31,176,30,176,29,112,31,129,31,129,30,104,31,88,31,215,31,149,31,250,31,76,31,149,31,103,31,175,31,31,31,110,31,117,31,77,31,248,31,100,31,15,31,228,31,73,31,73,30,55,31,55,30,198,31,78,31,233,31,80,31,18,31,94,31,205,31,179,31,15,31,58,31,194,31,228,31,9,31,171,31,173,31,202,31,202,31,115,31,249,31,162,31,28,31,28,30,164,31,164,30,56,31,211,31,196,31,37,31,37,30,37,31,113,31,145,31,198,31,198,30,9,31,9,30,111,31,111,30,250,31,151,31,109,31,186,31,167,31,184,31,22,31,231,31,117,31,28,31,56,31,56,30,179,31,234,31,38,31,184,31,152,31,216,31,18,31,200,31,129,31,195,31,173,31,27,31,26,31,26,30,26,29,223,31,86,31,139,31,120,31,244,31,244,30,161,31,125,31,125,30,107,31,125,31,232,31,232,30,153,31,192,31,192,30,138,31,138,30,94,31,98,31,98,30,98,29,13,31,13,30,185,31,186,31,186,30,33,31,224,31,224,30,223,31,203,31,105,31,10,31,41,31,63,31,19,31,19,30,176,31,59,31,160,31,211,31,227,31,73,31,73,30,37,31,137,31,92,31,92,30,43,31,129,31,178,31,17,31,57,31,175,31,129,31,129,30,76,31,84,31,218,31,47,31,89,31,89,30,216,31,202,31,189,31,249,31,165,31,165,30,165,29,240,31,240,30,89,31,80,31,233,31,60,31,36,31,162,31,184,31,214,31,85,31,29,31,18,31,197,31,130,31,154,31,200,31,223,31,223,30,190,31,190,31,247,31,69,31,234,31,182,31,230,31,235,31,187,31,187,30,34,31,221,31,160,31,106,31,117,31,117,30,186,31,219,31,219,30,123,31,130,31,253,31,61,31,61,30,171,31,213,31,219,31,219,30,74,31,74,30,110,31,188,31,51,31,83,31,33,31,141,31,141,30,235,31,61,31,113,31,255,31,255,30,140,31,201,31,61,31,85,31,29,31,161,31,124,31,5,31,67,31,189,31,174,31,122,31,66,31,66,30,141,31,45,31,106,31,193,31,96,31,102,31,210,31,48,31,200,31,200,30,29,31,129,31,251,31,228,31,202,31,22,31,22,30,22,29,60,31,60,30,60,29,124,31,124,30,231,31,231,30,231,29,231,28,51,31,5,31,5,30,204,31,246,31,192,31,192,30,249,31,106,31,250,31,162,31,162,30,80,31,147,31,211,31,99,31,163,31,114,31,114,30,192,31,164,31,148,31,190,31,69,31,69,30,209,31,106,31,85,31,85,30,29,31,61,31,47,31,47,30,57,31,24,31,24,30,119,31,222,31,191,31,93,31,158,31,140,31,48,31,179,31,179,30,215,31,215,30,233,31,107,31,89,31,212,31,212,30,250,31,48,31,213,31,76,31,35,31,179,31,31,31,186,31,112,31,134,31,240,31,42,31,84,31,47,31,217,31,82,31,254,31,210,31,66,31,138,31,81,31,100,31,100,30,144,31,144,30,153,31,49,31,176,31,2,31,194,31,81,31,226,31,230,31,45,31,45,30,132,31,132,30,173,31,166,31,186,31,163,31,163,30,80,31,54,31,54,30,218,31,45,31,163,31,163,30,109,31,188,31,127,31,177,31,177,30,202,31,153,31,1,31,48,31,41,31,130,31,63,31,79,31,79,30,131,31,140,31,101,31,253,31,43,31,178,31,178,30,22,31,22,30,212,31,6,31,169,31,160,31,39,31,39,30,182,31,182,30,142,31,39,31,153,31,153,30,183,31,183,30,31,31,223,31,223,30,244,31,144,31,210,31,21,31,125,31,195,31,72,31,72,30,206,31,68,31,228,31,152,31,152,30,232,31,232,30,163,31,247,31,247,30,247,29,169,31,144,31,101,31,47,31,239,31,107,31,188,31,7,31,37,31,37,30,100,31,230,31,207,31,171,31,31,31,219,31,144,31,144,30,4,31,228,31,165,31,8,31,253,31,253,30,5,31,229,31,73,31,73,30,73,29,73,28,187,31,58,31,58,30,58,29,204,31,118,31,244,31,89,31,89,30,89,29,208,31,208,30,30,31,223,31,1,31,83,31,229,31,229,30,229,29,229,28,246,31,238,31,144,31,144,30,67,31,67,30,234,31,78,31,116,31,116,31,95,31,37,31,148,31,117,31,19,31,250,31,194,31,194,30,103,31,58,31,72,31,145,31,237,31,51,31,82,31,236,31,175,31,110,31,167,31,167,30,167,29,34,31,34,30,91,31,4,31,16,31,90,31,74,31,164,31,66,31,156,31,138,31,254,31,58,31,233,31,108,31,191,31,114,31,50,31,121,31,186,31,38,31,65,31,227,31,105,31,105,30,105,29,105,28,164,31,40,31,119,31,188,31,58,31,218,31,218,30,102,31,253,31,39,31,39,30,129,31,129,30,221,31,184,31,102,31,160,31,182,31,182,30,62,31,135,31,109,31,71,31,71,30,176,31,176,30,136,31,146,31,146,30,22,31,228,31,105,31,92,31,164,31,10,31,10,30,104,31,176,31,182,31,182,30,228,31,228,30,7,31,192,31,192,30,229,31,21,31,21,30,21,29,251,31,123,31,49,31,49,30,153,31,84,31,84,30,250,31,76,31,83,31,83,30,249,31,82,31,210,31,51,31,51,30,51,29,205,31,205,30,205,29,142,31,125,31,125,30,11,31,97,31,49,31,179,31,29,31,29,30,99,31,43,31,43,30,69,31,69,30,69,29,12,31,200,31,229,31,152,31,142,31,142,30,13,31,44,31,11,31,26,31,37,31,107,31,159,31,117,31,3,31,4,31,4,30,172,31,13,31,161,31,165,31,145,31,44,31,197,31,50,31,170,31,172,31,219,31,219,30,44,31,10,31,154,31,223,31,142,31,142,30,190,31,25,31,239,31,103,31,112,31,9,31,150,31,72,31,72,30,38,31,83,31,150,31,140,31,45,31,99,31,206,31,76,31,121,31,184,31,105,31,148,31,148,30,21,31,14,31,205,31,169,31,169,30,169,29,119,31,201,31,92,31,124,31,124,30,98,31,117,31,174,31,186,31,186,30,186,29,134,31,134,30,193,31,193,30,93,31,128,31,17,31,17,30,17,29,17,28,183,31,119,31,247,31,183,31,183,30,173,31,190,31,190,30,125,31,202,31,63,31,90,31,186,31,40,31,158,31,220,31,160,31,160,30,47,31,74,31,74,30,193,31,193,30,204,31,59,31,155,31,202,31,202,30,111,31,100,31,203,31,23,31,23,30,23,29,23,28,173,31,169,31,53,31,222,31,151,31,151,30,139,31,112,31,207,31,207,30,49,31,182,31,109,31,219,31,40,31,138,31,194,31,209,31,209,30,238,31,245,31,25,31,135,31,34,31,2,31,2,30,183,31,18,31,24,31,96,31,198,31,250,31,147,31,183,31,179,31,179,30,179,29,154,31,60,31,60,30,176,31,105,31,254,31,42,31,188,31,41,31,41,30,234,31,226,31,12,31,12,30,54,31,54,30,12,31,125,31,125,30,37,31,37,30,238,31,176,31,229,31,58,31,241,31,241,30,197,31,234,31,234,30,234,29,219,31,219,30,219,29,216,31,121,31,121,30,46,31,16,31,117,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
