-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 830;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (111,0,186,0,233,0,77,0,197,0,0,0,174,0,240,0,57,0,0,0,148,0,137,0,4,0,182,0,7,0,0,0,15,0,135,0,145,0,71,0,67,0,62,0,62,0,4,0,0,0,64,0,241,0,0,0,134,0,34,0,83,0,0,0,192,0,97,0,178,0,57,0,163,0,159,0,71,0,0,0,46,0,138,0,126,0,174,0,255,0,135,0,2,0,0,0,148,0,0,0,0,0,0,0,8,0,0,0,228,0,22,0,0,0,165,0,122,0,76,0,116,0,88,0,111,0,101,0,63,0,0,0,185,0,0,0,0,0,0,0,0,0,0,0,106,0,84,0,0,0,30,0,214,0,139,0,44,0,99,0,0,0,66,0,219,0,0,0,200,0,200,0,229,0,0,0,210,0,30,0,0,0,0,0,2,0,105,0,48,0,0,0,111,0,119,0,0,0,137,0,0,0,0,0,206,0,45,0,2,0,130,0,218,0,63,0,110,0,248,0,235,0,0,0,240,0,248,0,184,0,242,0,209,0,216,0,176,0,0,0,240,0,170,0,178,0,4,0,254,0,59,0,0,0,103,0,204,0,239,0,169,0,147,0,42,0,92,0,160,0,98,0,0,0,0,0,3,0,15,0,77,0,173,0,0,0,0,0,148,0,204,0,242,0,0,0,197,0,206,0,233,0,118,0,237,0,16,0,83,0,240,0,116,0,0,0,20,0,80,0,98,0,230,0,0,0,0,0,64,0,125,0,59,0,0,0,44,0,183,0,104,0,229,0,161,0,242,0,211,0,0,0,245,0,0,0,63,0,16,0,162,0,122,0,66,0,159,0,146,0,0,0,16,0,145,0,104,0,43,0,55,0,0,0,124,0,250,0,0,0,182,0,191,0,0,0,23,0,1,0,64,0,132,0,98,0,242,0,0,0,25,0,224,0,146,0,0,0,0,0,26,0,173,0,0,0,136,0,245,0,36,0,113,0,0,0,146,0,28,0,0,0,55,0,126,0,49,0,211,0,164,0,61,0,197,0,217,0,0,0,211,0,66,0,187,0,140,0,93,0,110,0,137,0,96,0,34,0,22,0,243,0,253,0,142,0,29,0,95,0,246,0,1,0,0,0,220,0,23,0,188,0,0,0,0,0,44,0,50,0,170,0,133,0,88,0,162,0,20,0,71,0,155,0,169,0,234,0,0,0,64,0,186,0,68,0,204,0,227,0,15,0,0,0,134,0,168,0,20,0,106,0,74,0,96,0,0,0,0,0,0,0,97,0,85,0,14,0,0,0,218,0,0,0,0,0,0,0,0,0,93,0,30,0,116,0,207,0,16,0,242,0,0,0,195,0,0,0,170,0,0,0,0,0,187,0,214,0,40,0,23,0,0,0,24,0,208,0,188,0,165,0,254,0,37,0,0,0,102,0,188,0,242,0,145,0,7,0,0,0,146,0,0,0,154,0,0,0,40,0,128,0,244,0,153,0,203,0,69,0,96,0,205,0,0,0,188,0,36,0,239,0,107,0,92,0,27,0,138,0,56,0,14,0,156,0,31,0,191,0,18,0,33,0,219,0,199,0,20,0,241,0,0,0,56,0,226,0,0,0,0,0,57,0,67,0,0,0,127,0,250,0,35,0,223,0,79,0,64,0,0,0,53,0,23,0,88,0,136,0,2,0,52,0,61,0,222,0,169,0,123,0,46,0,34,0,0,0,98,0,0,0,173,0,199,0,230,0,48,0,209,0,54,0,111,0,252,0,230,0,79,0,9,0,149,0,0,0,113,0,138,0,233,0,50,0,101,0,0,0,175,0,22,0,0,0,213,0,228,0,97,0,16,0,170,0,105,0,233,0,229,0,0,0,197,0,0,0,0,0,157,0,113,0,24,0,52,0,78,0,172,0,102,0,40,0,0,0,127,0,222,0,0,0,25,0,172,0,154,0,230,0,0,0,176,0,0,0,166,0,38,0,134,0,11,0,188,0,53,0,137,0,91,0,112,0,123,0,195,0,181,0,147,0,160,0,140,0,156,0,80,0,0,0,0,0,170,0,183,0,113,0,0,0,32,0,25,0,19,0,202,0,61,0,149,0,52,0,0,0,159,0,12,0,182,0,218,0,199,0,55,0,18,0,234,0,154,0,106,0,220,0,128,0,178,0,0,0,67,0,0,0,215,0,86,0,169,0,139,0,108,0,4,0,0,0,0,0,133,0,36,0,0,0,0,0,0,0,154,0,2,0,0,0,98,0,0,0,214,0,0,0,0,0,164,0,107,0,66,0,0,0,189,0,150,0,13,0,129,0,0,0,105,0,164,0,178,0,0,0,46,0,19,0,152,0,138,0,252,0,161,0,150,0,0,0,31,0,91,0,213,0,126,0,0,0,28,0,80,0,31,0,0,0,201,0,83,0,61,0,129,0,170,0,0,0,182,0,94,0,45,0,197,0,44,0,234,0,247,0,64,0,33,0,51,0,0,0,0,0,118,0,0,0,222,0,182,0,0,0,0,0,239,0,0,0,66,0,99,0,0,0,207,0,51,0,0,0,232,0,117,0,0,0,5,0,0,0,220,0,85,0,108,0,0,0,186,0,148,0,137,0,204,0,0,0,175,0,193,0,16,0,36,0,207,0,235,0,0,0,91,0,83,0,0,0,118,0,108,0,232,0,0,0,154,0,125,0,85,0,191,0,53,0,73,0,213,0,0,0,0,0,243,0,0,0,160,0,92,0,69,0,231,0,209,0,157,0,70,0,194,0,126,0,247,0,0,0,139,0,135,0,35,0,159,0,52,0,245,0,24,0,0,0,28,0,0,0,53,0,182,0,72,0,35,0,218,0,57,0,1,0,140,0,126,0,19,0,204,0,33,0,72,0,174,0,156,0,0,0,114,0,88,0,34,0,0,0,62,0,0,0,2,0,0,0,0,0,0,0,103,0,0,0,57,0,242,0,25,0,231,0,31,0,139,0,251,0,114,0,0,0,0,0,6,0,48,0,0,0,251,0,140,0,82,0,207,0,99,0,118,0,0,0,0,0,227,0,142,0,71,0,207,0,89,0,0,0,119,0,106,0,72,0,66,0,0,0,239,0,138,0,101,0,136,0,210,0,238,0,0,0,124,0,0,0,88,0,111,0,1,0,228,0,198,0,0,0,248,0,173,0,0,0,92,0,22,0,75,0,0,0,193,0,89,0,0,0,0,0,154,0,0,0,89,0,0,0,67,0,153,0,209,0,174,0,243,0,7,0,238,0,201,0,37,0,1,0,144,0,93,0,66,0,175,0,228,0,0,0,104,0,219,0,78,0,0,0,233,0,38,0,144,0,121,0,0,0,11,0,97,0,205,0,59,0,50,0,218,0,145,0,240,0,0,0,0,0,169,0,255,0,149,0,15,0,64,0,94,0,75,0,34,0,0,0,107,0,9,0,54,0,252,0,56,0,0,0,223,0,238,0,161,0,36,0,48,0,5,0,184,0,171,0,18,0,20,0,40,0,114,0,0,0,187,0,123,0,113,0,182,0,109,0,0,0,178,0,0,0,135,0,158,0,241,0,168,0,14,0,0,0,0,0,0,0,79,0,0,0,2,0,41,0,181,0,23,0,56,0,196,0,187,0,0,0,74,0,129,0,0,0,217,0,139,0,182,0,188,0,109,0,3,0,0,0,236,0,22,0,146,0,156,0,0,0,0,0,9,0,122,0,205,0,45,0,60,0,246,0,73,0,130,0,177,0,183,0,0,0);
signal scenario_full  : scenario_type := (111,31,186,31,233,31,77,31,197,31,197,30,174,31,240,31,57,31,57,30,148,31,137,31,4,31,182,31,7,31,7,30,15,31,135,31,145,31,71,31,67,31,62,31,62,31,4,31,4,30,64,31,241,31,241,30,134,31,34,31,83,31,83,30,192,31,97,31,178,31,57,31,163,31,159,31,71,31,71,30,46,31,138,31,126,31,174,31,255,31,135,31,2,31,2,30,148,31,148,30,148,29,148,28,8,31,8,30,228,31,22,31,22,30,165,31,122,31,76,31,116,31,88,31,111,31,101,31,63,31,63,30,185,31,185,30,185,29,185,28,185,27,185,26,106,31,84,31,84,30,30,31,214,31,139,31,44,31,99,31,99,30,66,31,219,31,219,30,200,31,200,31,229,31,229,30,210,31,30,31,30,30,30,29,2,31,105,31,48,31,48,30,111,31,119,31,119,30,137,31,137,30,137,29,206,31,45,31,2,31,130,31,218,31,63,31,110,31,248,31,235,31,235,30,240,31,248,31,184,31,242,31,209,31,216,31,176,31,176,30,240,31,170,31,178,31,4,31,254,31,59,31,59,30,103,31,204,31,239,31,169,31,147,31,42,31,92,31,160,31,98,31,98,30,98,29,3,31,15,31,77,31,173,31,173,30,173,29,148,31,204,31,242,31,242,30,197,31,206,31,233,31,118,31,237,31,16,31,83,31,240,31,116,31,116,30,20,31,80,31,98,31,230,31,230,30,230,29,64,31,125,31,59,31,59,30,44,31,183,31,104,31,229,31,161,31,242,31,211,31,211,30,245,31,245,30,63,31,16,31,162,31,122,31,66,31,159,31,146,31,146,30,16,31,145,31,104,31,43,31,55,31,55,30,124,31,250,31,250,30,182,31,191,31,191,30,23,31,1,31,64,31,132,31,98,31,242,31,242,30,25,31,224,31,146,31,146,30,146,29,26,31,173,31,173,30,136,31,245,31,36,31,113,31,113,30,146,31,28,31,28,30,55,31,126,31,49,31,211,31,164,31,61,31,197,31,217,31,217,30,211,31,66,31,187,31,140,31,93,31,110,31,137,31,96,31,34,31,22,31,243,31,253,31,142,31,29,31,95,31,246,31,1,31,1,30,220,31,23,31,188,31,188,30,188,29,44,31,50,31,170,31,133,31,88,31,162,31,20,31,71,31,155,31,169,31,234,31,234,30,64,31,186,31,68,31,204,31,227,31,15,31,15,30,134,31,168,31,20,31,106,31,74,31,96,31,96,30,96,29,96,28,97,31,85,31,14,31,14,30,218,31,218,30,218,29,218,28,218,27,93,31,30,31,116,31,207,31,16,31,242,31,242,30,195,31,195,30,170,31,170,30,170,29,187,31,214,31,40,31,23,31,23,30,24,31,208,31,188,31,165,31,254,31,37,31,37,30,102,31,188,31,242,31,145,31,7,31,7,30,146,31,146,30,154,31,154,30,40,31,128,31,244,31,153,31,203,31,69,31,96,31,205,31,205,30,188,31,36,31,239,31,107,31,92,31,27,31,138,31,56,31,14,31,156,31,31,31,191,31,18,31,33,31,219,31,199,31,20,31,241,31,241,30,56,31,226,31,226,30,226,29,57,31,67,31,67,30,127,31,250,31,35,31,223,31,79,31,64,31,64,30,53,31,23,31,88,31,136,31,2,31,52,31,61,31,222,31,169,31,123,31,46,31,34,31,34,30,98,31,98,30,173,31,199,31,230,31,48,31,209,31,54,31,111,31,252,31,230,31,79,31,9,31,149,31,149,30,113,31,138,31,233,31,50,31,101,31,101,30,175,31,22,31,22,30,213,31,228,31,97,31,16,31,170,31,105,31,233,31,229,31,229,30,197,31,197,30,197,29,157,31,113,31,24,31,52,31,78,31,172,31,102,31,40,31,40,30,127,31,222,31,222,30,25,31,172,31,154,31,230,31,230,30,176,31,176,30,166,31,38,31,134,31,11,31,188,31,53,31,137,31,91,31,112,31,123,31,195,31,181,31,147,31,160,31,140,31,156,31,80,31,80,30,80,29,170,31,183,31,113,31,113,30,32,31,25,31,19,31,202,31,61,31,149,31,52,31,52,30,159,31,12,31,182,31,218,31,199,31,55,31,18,31,234,31,154,31,106,31,220,31,128,31,178,31,178,30,67,31,67,30,215,31,86,31,169,31,139,31,108,31,4,31,4,30,4,29,133,31,36,31,36,30,36,29,36,28,154,31,2,31,2,30,98,31,98,30,214,31,214,30,214,29,164,31,107,31,66,31,66,30,189,31,150,31,13,31,129,31,129,30,105,31,164,31,178,31,178,30,46,31,19,31,152,31,138,31,252,31,161,31,150,31,150,30,31,31,91,31,213,31,126,31,126,30,28,31,80,31,31,31,31,30,201,31,83,31,61,31,129,31,170,31,170,30,182,31,94,31,45,31,197,31,44,31,234,31,247,31,64,31,33,31,51,31,51,30,51,29,118,31,118,30,222,31,182,31,182,30,182,29,239,31,239,30,66,31,99,31,99,30,207,31,51,31,51,30,232,31,117,31,117,30,5,31,5,30,220,31,85,31,108,31,108,30,186,31,148,31,137,31,204,31,204,30,175,31,193,31,16,31,36,31,207,31,235,31,235,30,91,31,83,31,83,30,118,31,108,31,232,31,232,30,154,31,125,31,85,31,191,31,53,31,73,31,213,31,213,30,213,29,243,31,243,30,160,31,92,31,69,31,231,31,209,31,157,31,70,31,194,31,126,31,247,31,247,30,139,31,135,31,35,31,159,31,52,31,245,31,24,31,24,30,28,31,28,30,53,31,182,31,72,31,35,31,218,31,57,31,1,31,140,31,126,31,19,31,204,31,33,31,72,31,174,31,156,31,156,30,114,31,88,31,34,31,34,30,62,31,62,30,2,31,2,30,2,29,2,28,103,31,103,30,57,31,242,31,25,31,231,31,31,31,139,31,251,31,114,31,114,30,114,29,6,31,48,31,48,30,251,31,140,31,82,31,207,31,99,31,118,31,118,30,118,29,227,31,142,31,71,31,207,31,89,31,89,30,119,31,106,31,72,31,66,31,66,30,239,31,138,31,101,31,136,31,210,31,238,31,238,30,124,31,124,30,88,31,111,31,1,31,228,31,198,31,198,30,248,31,173,31,173,30,92,31,22,31,75,31,75,30,193,31,89,31,89,30,89,29,154,31,154,30,89,31,89,30,67,31,153,31,209,31,174,31,243,31,7,31,238,31,201,31,37,31,1,31,144,31,93,31,66,31,175,31,228,31,228,30,104,31,219,31,78,31,78,30,233,31,38,31,144,31,121,31,121,30,11,31,97,31,205,31,59,31,50,31,218,31,145,31,240,31,240,30,240,29,169,31,255,31,149,31,15,31,64,31,94,31,75,31,34,31,34,30,107,31,9,31,54,31,252,31,56,31,56,30,223,31,238,31,161,31,36,31,48,31,5,31,184,31,171,31,18,31,20,31,40,31,114,31,114,30,187,31,123,31,113,31,182,31,109,31,109,30,178,31,178,30,135,31,158,31,241,31,168,31,14,31,14,30,14,29,14,28,79,31,79,30,2,31,41,31,181,31,23,31,56,31,196,31,187,31,187,30,74,31,129,31,129,30,217,31,139,31,182,31,188,31,109,31,3,31,3,30,236,31,22,31,146,31,156,31,156,30,156,29,9,31,122,31,205,31,45,31,60,31,246,31,73,31,130,31,177,31,183,31,183,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
