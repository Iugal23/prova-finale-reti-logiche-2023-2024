-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_711 is
end project_tb_711;

architecture project_tb_arch_711 of project_tb_711 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 506;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (79,0,68,0,193,0,26,0,0,0,223,0,240,0,91,0,179,0,92,0,51,0,9,0,81,0,112,0,147,0,248,0,221,0,93,0,159,0,72,0,0,0,24,0,98,0,0,0,108,0,45,0,134,0,183,0,54,0,0,0,104,0,206,0,168,0,213,0,148,0,0,0,147,0,0,0,0,0,69,0,93,0,93,0,30,0,253,0,210,0,0,0,72,0,83,0,78,0,183,0,33,0,220,0,226,0,0,0,0,0,0,0,0,0,77,0,174,0,0,0,236,0,0,0,0,0,229,0,86,0,11,0,106,0,55,0,188,0,34,0,47,0,103,0,96,0,148,0,0,0,85,0,33,0,55,0,242,0,0,0,232,0,171,0,0,0,73,0,0,0,85,0,0,0,98,0,35,0,175,0,46,0,0,0,242,0,146,0,18,0,23,0,244,0,27,0,196,0,82,0,105,0,0,0,60,0,241,0,2,0,206,0,0,0,119,0,147,0,205,0,48,0,242,0,30,0,46,0,119,0,203,0,0,0,29,0,94,0,6,0,246,0,0,0,211,0,0,0,13,0,0,0,4,0,34,0,0,0,65,0,32,0,40,0,135,0,240,0,164,0,50,0,83,0,0,0,131,0,229,0,0,0,0,0,20,0,83,0,161,0,246,0,186,0,97,0,210,0,185,0,177,0,250,0,0,0,164,0,0,0,86,0,214,0,117,0,18,0,218,0,0,0,0,0,214,0,57,0,0,0,180,0,155,0,177,0,0,0,179,0,136,0,0,0,0,0,0,0,0,0,0,0,164,0,0,0,68,0,205,0,0,0,241,0,229,0,78,0,15,0,0,0,165,0,160,0,228,0,208,0,89,0,17,0,228,0,158,0,0,0,208,0,0,0,129,0,68,0,197,0,83,0,39,0,194,0,0,0,82,0,0,0,155,0,148,0,243,0,56,0,36,0,34,0,238,0,0,0,77,0,54,0,245,0,64,0,0,0,0,0,232,0,0,0,38,0,246,0,0,0,0,0,163,0,68,0,65,0,51,0,194,0,247,0,172,0,73,0,0,0,0,0,108,0,121,0,85,0,190,0,0,0,248,0,247,0,128,0,0,0,0,0,167,0,230,0,0,0,181,0,59,0,122,0,144,0,154,0,229,0,63,0,114,0,173,0,221,0,128,0,56,0,0,0,255,0,207,0,214,0,47,0,0,0,241,0,207,0,113,0,168,0,244,0,180,0,119,0,29,0,24,0,6,0,50,0,139,0,218,0,0,0,97,0,138,0,236,0,162,0,0,0,49,0,60,0,24,0,0,0,30,0,164,0,0,0,30,0,4,0,255,0,101,0,110,0,84,0,239,0,47,0,0,0,0,0,130,0,0,0,240,0,54,0,127,0,11,0,215,0,112,0,91,0,0,0,0,0,139,0,100,0,0,0,0,0,91,0,242,0,127,0,200,0,0,0,20,0,230,0,32,0,22,0,127,0,197,0,10,0,54,0,227,0,3,0,91,0,58,0,51,0,113,0,194,0,108,0,152,0,180,0,234,0,252,0,172,0,231,0,146,0,68,0,248,0,0,0,6,0,0,0,0,0,89,0,246,0,212,0,180,0,243,0,184,0,0,0,175,0,80,0,44,0,248,0,126,0,146,0,1,0,84,0,99,0,0,0,196,0,212,0,186,0,143,0,25,0,133,0,109,0,184,0,136,0,134,0,0,0,138,0,62,0,92,0,197,0,204,0,0,0,66,0,58,0,89,0,173,0,174,0,0,0,154,0,0,0,184,0,191,0,198,0,96,0,68,0,0,0,115,0,148,0,0,0,18,0,8,0,231,0,81,0,0,0,192,0,99,0,93,0,0,0,114,0,108,0,149,0,159,0,66,0,125,0,205,0,230,0,7,0,63,0,14,0,73,0,108,0,182,0,226,0,68,0,148,0,0,0,38,0,23,0,0,0,143,0,139,0,7,0,104,0,0,0,207,0,0,0,108,0,0,0,58,0,52,0,0,0,0,0,154,0,218,0,242,0,36,0,3,0,46,0,0,0,42,0,0,0,8,0,0,0,82,0,119,0,0,0,184,0,181,0,218,0,97,0,110,0,246,0,212,0,237,0,59,0,70,0,39,0,152,0,96,0,186,0,0,0,97,0,0,0,0,0,0,0,106,0,136,0,0,0,57,0,142,0,147,0,245,0,12,0,81,0,172,0,26,0,0,0,226,0,192,0,240,0,29,0,96,0,30,0,67,0,203,0,71,0,0,0,0,0,109,0,138,0,0,0,204,0);
signal scenario_full  : scenario_type := (79,31,68,31,193,31,26,31,26,30,223,31,240,31,91,31,179,31,92,31,51,31,9,31,81,31,112,31,147,31,248,31,221,31,93,31,159,31,72,31,72,30,24,31,98,31,98,30,108,31,45,31,134,31,183,31,54,31,54,30,104,31,206,31,168,31,213,31,148,31,148,30,147,31,147,30,147,29,69,31,93,31,93,31,30,31,253,31,210,31,210,30,72,31,83,31,78,31,183,31,33,31,220,31,226,31,226,30,226,29,226,28,226,27,77,31,174,31,174,30,236,31,236,30,236,29,229,31,86,31,11,31,106,31,55,31,188,31,34,31,47,31,103,31,96,31,148,31,148,30,85,31,33,31,55,31,242,31,242,30,232,31,171,31,171,30,73,31,73,30,85,31,85,30,98,31,35,31,175,31,46,31,46,30,242,31,146,31,18,31,23,31,244,31,27,31,196,31,82,31,105,31,105,30,60,31,241,31,2,31,206,31,206,30,119,31,147,31,205,31,48,31,242,31,30,31,46,31,119,31,203,31,203,30,29,31,94,31,6,31,246,31,246,30,211,31,211,30,13,31,13,30,4,31,34,31,34,30,65,31,32,31,40,31,135,31,240,31,164,31,50,31,83,31,83,30,131,31,229,31,229,30,229,29,20,31,83,31,161,31,246,31,186,31,97,31,210,31,185,31,177,31,250,31,250,30,164,31,164,30,86,31,214,31,117,31,18,31,218,31,218,30,218,29,214,31,57,31,57,30,180,31,155,31,177,31,177,30,179,31,136,31,136,30,136,29,136,28,136,27,136,26,164,31,164,30,68,31,205,31,205,30,241,31,229,31,78,31,15,31,15,30,165,31,160,31,228,31,208,31,89,31,17,31,228,31,158,31,158,30,208,31,208,30,129,31,68,31,197,31,83,31,39,31,194,31,194,30,82,31,82,30,155,31,148,31,243,31,56,31,36,31,34,31,238,31,238,30,77,31,54,31,245,31,64,31,64,30,64,29,232,31,232,30,38,31,246,31,246,30,246,29,163,31,68,31,65,31,51,31,194,31,247,31,172,31,73,31,73,30,73,29,108,31,121,31,85,31,190,31,190,30,248,31,247,31,128,31,128,30,128,29,167,31,230,31,230,30,181,31,59,31,122,31,144,31,154,31,229,31,63,31,114,31,173,31,221,31,128,31,56,31,56,30,255,31,207,31,214,31,47,31,47,30,241,31,207,31,113,31,168,31,244,31,180,31,119,31,29,31,24,31,6,31,50,31,139,31,218,31,218,30,97,31,138,31,236,31,162,31,162,30,49,31,60,31,24,31,24,30,30,31,164,31,164,30,30,31,4,31,255,31,101,31,110,31,84,31,239,31,47,31,47,30,47,29,130,31,130,30,240,31,54,31,127,31,11,31,215,31,112,31,91,31,91,30,91,29,139,31,100,31,100,30,100,29,91,31,242,31,127,31,200,31,200,30,20,31,230,31,32,31,22,31,127,31,197,31,10,31,54,31,227,31,3,31,91,31,58,31,51,31,113,31,194,31,108,31,152,31,180,31,234,31,252,31,172,31,231,31,146,31,68,31,248,31,248,30,6,31,6,30,6,29,89,31,246,31,212,31,180,31,243,31,184,31,184,30,175,31,80,31,44,31,248,31,126,31,146,31,1,31,84,31,99,31,99,30,196,31,212,31,186,31,143,31,25,31,133,31,109,31,184,31,136,31,134,31,134,30,138,31,62,31,92,31,197,31,204,31,204,30,66,31,58,31,89,31,173,31,174,31,174,30,154,31,154,30,184,31,191,31,198,31,96,31,68,31,68,30,115,31,148,31,148,30,18,31,8,31,231,31,81,31,81,30,192,31,99,31,93,31,93,30,114,31,108,31,149,31,159,31,66,31,125,31,205,31,230,31,7,31,63,31,14,31,73,31,108,31,182,31,226,31,68,31,148,31,148,30,38,31,23,31,23,30,143,31,139,31,7,31,104,31,104,30,207,31,207,30,108,31,108,30,58,31,52,31,52,30,52,29,154,31,218,31,242,31,36,31,3,31,46,31,46,30,42,31,42,30,8,31,8,30,82,31,119,31,119,30,184,31,181,31,218,31,97,31,110,31,246,31,212,31,237,31,59,31,70,31,39,31,152,31,96,31,186,31,186,30,97,31,97,30,97,29,97,28,106,31,136,31,136,30,57,31,142,31,147,31,245,31,12,31,81,31,172,31,26,31,26,30,226,31,192,31,240,31,29,31,96,31,30,31,67,31,203,31,71,31,71,30,71,29,109,31,138,31,138,30,204,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
