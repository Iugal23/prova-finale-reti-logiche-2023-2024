-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_691 is
end project_tb_691;

architecture project_tb_arch_691 of project_tb_691 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 520;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (237,0,16,0,230,0,119,0,148,0,23,0,212,0,82,0,179,0,0,0,145,0,169,0,97,0,233,0,138,0,103,0,0,0,141,0,154,0,155,0,143,0,52,0,220,0,0,0,68,0,0,0,13,0,205,0,0,0,0,0,185,0,204,0,34,0,202,0,103,0,61,0,248,0,0,0,204,0,0,0,0,0,0,0,0,0,211,0,156,0,133,0,93,0,0,0,223,0,123,0,0,0,65,0,229,0,0,0,136,0,225,0,206,0,237,0,189,0,88,0,54,0,0,0,227,0,167,0,192,0,216,0,107,0,181,0,225,0,61,0,147,0,213,0,27,0,141,0,0,0,91,0,135,0,165,0,171,0,145,0,41,0,105,0,132,0,64,0,189,0,38,0,0,0,248,0,220,0,0,0,88,0,105,0,121,0,247,0,246,0,113,0,32,0,166,0,146,0,227,0,86,0,172,0,214,0,0,0,173,0,82,0,93,0,0,0,0,0,0,0,0,0,225,0,72,0,233,0,91,0,69,0,41,0,0,0,175,0,0,0,133,0,162,0,22,0,214,0,113,0,18,0,27,0,237,0,161,0,162,0,0,0,195,0,118,0,225,0,190,0,43,0,138,0,0,0,0,0,96,0,239,0,230,0,185,0,225,0,212,0,200,0,49,0,205,0,160,0,0,0,66,0,83,0,181,0,63,0,182,0,167,0,0,0,199,0,10,0,156,0,175,0,0,0,12,0,85,0,103,0,192,0,70,0,184,0,240,0,133,0,0,0,0,0,0,0,199,0,0,0,28,0,236,0,22,0,126,0,0,0,0,0,82,0,98,0,240,0,161,0,176,0,0,0,82,0,86,0,77,0,218,0,136,0,0,0,212,0,178,0,215,0,90,0,246,0,182,0,254,0,9,0,0,0,13,0,32,0,147,0,58,0,163,0,92,0,0,0,0,0,204,0,71,0,0,0,229,0,255,0,0,0,158,0,148,0,250,0,142,0,230,0,0,0,30,0,143,0,255,0,0,0,218,0,123,0,0,0,1,0,177,0,0,0,70,0,255,0,121,0,145,0,215,0,224,0,217,0,192,0,175,0,13,0,201,0,42,0,222,0,97,0,10,0,0,0,77,0,135,0,123,0,137,0,0,0,48,0,59,0,0,0,98,0,169,0,134,0,85,0,220,0,53,0,235,0,182,0,129,0,180,0,24,0,57,0,0,0,206,0,114,0,166,0,191,0,15,0,0,0,89,0,168,0,29,0,183,0,127,0,53,0,243,0,118,0,172,0,0,0,106,0,25,0,88,0,0,0,71,0,166,0,0,0,237,0,0,0,252,0,238,0,0,0,64,0,59,0,123,0,197,0,44,0,56,0,64,0,205,0,0,0,5,0,86,0,114,0,73,0,0,0,51,0,244,0,0,0,244,0,172,0,181,0,42,0,65,0,215,0,0,0,214,0,210,0,85,0,152,0,113,0,217,0,88,0,249,0,81,0,167,0,103,0,102,0,0,0,0,0,190,0,142,0,9,0,71,0,161,0,31,0,170,0,90,0,204,0,204,0,139,0,178,0,253,0,21,0,213,0,0,0,68,0,120,0,48,0,10,0,239,0,0,0,0,0,45,0,0,0,111,0,187,0,85,0,198,0,189,0,27,0,46,0,53,0,0,0,0,0,9,0,124,0,0,0,93,0,166,0,130,0,95,0,0,0,0,0,202,0,235,0,0,0,112,0,37,0,222,0,188,0,0,0,3,0,255,0,0,0,0,0,34,0,0,0,0,0,117,0,0,0,0,0,0,0,206,0,217,0,0,0,46,0,21,0,216,0,137,0,90,0,0,0,201,0,210,0,0,0,42,0,145,0,0,0,125,0,0,0,17,0,0,0,27,0,210,0,24,0,133,0,0,0,56,0,154,0,198,0,25,0,136,0,85,0,82,0,48,0,154,0,174,0,192,0,56,0,133,0,0,0,219,0,215,0,206,0,148,0,244,0,237,0,110,0,109,0,0,0,173,0,139,0,194,0,0,0,216,0,25,0,0,0,127,0,183,0,213,0,42,0,0,0,12,0,145,0,172,0,138,0,185,0,49,0,98,0,174,0,184,0,150,0,175,0,59,0,0,0,0,0,39,0,75,0,0,0,0,0,190,0,100,0,242,0,177,0,39,0,0,0,0,0,0,0,0,0,0,0,227,0,214,0,0,0,14,0,172,0,175,0,42,0,201,0,77,0,250,0,55,0,0,0,83,0,238,0,112,0,191,0,253,0,174,0,0,0,33,0,0,0,103,0,0,0,202,0,0,0,10,0,0,0,141,0,122,0,118,0,187,0,121,0,200,0,0,0,30,0);
signal scenario_full  : scenario_type := (237,31,16,31,230,31,119,31,148,31,23,31,212,31,82,31,179,31,179,30,145,31,169,31,97,31,233,31,138,31,103,31,103,30,141,31,154,31,155,31,143,31,52,31,220,31,220,30,68,31,68,30,13,31,205,31,205,30,205,29,185,31,204,31,34,31,202,31,103,31,61,31,248,31,248,30,204,31,204,30,204,29,204,28,204,27,211,31,156,31,133,31,93,31,93,30,223,31,123,31,123,30,65,31,229,31,229,30,136,31,225,31,206,31,237,31,189,31,88,31,54,31,54,30,227,31,167,31,192,31,216,31,107,31,181,31,225,31,61,31,147,31,213,31,27,31,141,31,141,30,91,31,135,31,165,31,171,31,145,31,41,31,105,31,132,31,64,31,189,31,38,31,38,30,248,31,220,31,220,30,88,31,105,31,121,31,247,31,246,31,113,31,32,31,166,31,146,31,227,31,86,31,172,31,214,31,214,30,173,31,82,31,93,31,93,30,93,29,93,28,93,27,225,31,72,31,233,31,91,31,69,31,41,31,41,30,175,31,175,30,133,31,162,31,22,31,214,31,113,31,18,31,27,31,237,31,161,31,162,31,162,30,195,31,118,31,225,31,190,31,43,31,138,31,138,30,138,29,96,31,239,31,230,31,185,31,225,31,212,31,200,31,49,31,205,31,160,31,160,30,66,31,83,31,181,31,63,31,182,31,167,31,167,30,199,31,10,31,156,31,175,31,175,30,12,31,85,31,103,31,192,31,70,31,184,31,240,31,133,31,133,30,133,29,133,28,199,31,199,30,28,31,236,31,22,31,126,31,126,30,126,29,82,31,98,31,240,31,161,31,176,31,176,30,82,31,86,31,77,31,218,31,136,31,136,30,212,31,178,31,215,31,90,31,246,31,182,31,254,31,9,31,9,30,13,31,32,31,147,31,58,31,163,31,92,31,92,30,92,29,204,31,71,31,71,30,229,31,255,31,255,30,158,31,148,31,250,31,142,31,230,31,230,30,30,31,143,31,255,31,255,30,218,31,123,31,123,30,1,31,177,31,177,30,70,31,255,31,121,31,145,31,215,31,224,31,217,31,192,31,175,31,13,31,201,31,42,31,222,31,97,31,10,31,10,30,77,31,135,31,123,31,137,31,137,30,48,31,59,31,59,30,98,31,169,31,134,31,85,31,220,31,53,31,235,31,182,31,129,31,180,31,24,31,57,31,57,30,206,31,114,31,166,31,191,31,15,31,15,30,89,31,168,31,29,31,183,31,127,31,53,31,243,31,118,31,172,31,172,30,106,31,25,31,88,31,88,30,71,31,166,31,166,30,237,31,237,30,252,31,238,31,238,30,64,31,59,31,123,31,197,31,44,31,56,31,64,31,205,31,205,30,5,31,86,31,114,31,73,31,73,30,51,31,244,31,244,30,244,31,172,31,181,31,42,31,65,31,215,31,215,30,214,31,210,31,85,31,152,31,113,31,217,31,88,31,249,31,81,31,167,31,103,31,102,31,102,30,102,29,190,31,142,31,9,31,71,31,161,31,31,31,170,31,90,31,204,31,204,31,139,31,178,31,253,31,21,31,213,31,213,30,68,31,120,31,48,31,10,31,239,31,239,30,239,29,45,31,45,30,111,31,187,31,85,31,198,31,189,31,27,31,46,31,53,31,53,30,53,29,9,31,124,31,124,30,93,31,166,31,130,31,95,31,95,30,95,29,202,31,235,31,235,30,112,31,37,31,222,31,188,31,188,30,3,31,255,31,255,30,255,29,34,31,34,30,34,29,117,31,117,30,117,29,117,28,206,31,217,31,217,30,46,31,21,31,216,31,137,31,90,31,90,30,201,31,210,31,210,30,42,31,145,31,145,30,125,31,125,30,17,31,17,30,27,31,210,31,24,31,133,31,133,30,56,31,154,31,198,31,25,31,136,31,85,31,82,31,48,31,154,31,174,31,192,31,56,31,133,31,133,30,219,31,215,31,206,31,148,31,244,31,237,31,110,31,109,31,109,30,173,31,139,31,194,31,194,30,216,31,25,31,25,30,127,31,183,31,213,31,42,31,42,30,12,31,145,31,172,31,138,31,185,31,49,31,98,31,174,31,184,31,150,31,175,31,59,31,59,30,59,29,39,31,75,31,75,30,75,29,190,31,100,31,242,31,177,31,39,31,39,30,39,29,39,28,39,27,39,26,227,31,214,31,214,30,14,31,172,31,175,31,42,31,201,31,77,31,250,31,55,31,55,30,83,31,238,31,112,31,191,31,253,31,174,31,174,30,33,31,33,30,103,31,103,30,202,31,202,30,10,31,10,30,141,31,122,31,118,31,187,31,121,31,200,31,200,30,30,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
