-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_681 is
end project_tb_681;

architecture project_tb_arch_681 of project_tb_681 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 673;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (147,0,0,0,114,0,0,0,0,0,70,0,0,0,24,0,0,0,21,0,14,0,187,0,0,0,27,0,111,0,54,0,21,0,74,0,238,0,0,0,76,0,28,0,122,0,185,0,175,0,0,0,19,0,84,0,211,0,160,0,134,0,0,0,17,0,0,0,4,0,86,0,243,0,178,0,152,0,175,0,52,0,118,0,29,0,210,0,118,0,35,0,244,0,0,0,184,0,154,0,35,0,0,0,115,0,0,0,175,0,106,0,191,0,18,0,188,0,112,0,7,0,46,0,121,0,255,0,206,0,76,0,197,0,0,0,53,0,0,0,173,0,0,0,252,0,0,0,133,0,30,0,169,0,101,0,113,0,42,0,228,0,0,0,0,0,52,0,220,0,0,0,246,0,0,0,144,0,70,0,187,0,192,0,228,0,139,0,225,0,13,0,247,0,114,0,18,0,182,0,0,0,61,0,0,0,192,0,43,0,199,0,227,0,86,0,0,0,221,0,193,0,96,0,191,0,54,0,45,0,0,0,7,0,0,0,76,0,0,0,36,0,200,0,0,0,0,0,113,0,250,0,67,0,67,0,178,0,0,0,191,0,25,0,0,0,0,0,43,0,0,0,122,0,203,0,48,0,119,0,248,0,153,0,168,0,0,0,0,0,0,0,71,0,220,0,244,0,59,0,72,0,0,0,160,0,35,0,239,0,0,0,197,0,77,0,0,0,246,0,114,0,203,0,180,0,65,0,177,0,0,0,248,0,64,0,21,0,156,0,209,0,0,0,0,0,35,0,183,0,0,0,0,0,86,0,152,0,191,0,106,0,212,0,159,0,228,0,100,0,0,0,4,0,166,0,0,0,186,0,215,0,184,0,133,0,48,0,246,0,71,0,185,0,5,0,24,0,254,0,68,0,107,0,78,0,134,0,79,0,253,0,198,0,175,0,96,0,148,0,190,0,247,0,111,0,80,0,103,0,178,0,0,0,76,0,0,0,0,0,0,0,96,0,242,0,0,0,0,0,134,0,226,0,119,0,109,0,38,0,126,0,134,0,4,0,206,0,162,0,210,0,248,0,239,0,108,0,209,0,56,0,27,0,189,0,119,0,56,0,53,0,169,0,237,0,89,0,116,0,231,0,0,0,183,0,6,0,213,0,0,0,117,0,181,0,37,0,97,0,0,0,22,0,168,0,90,0,0,0,229,0,136,0,32,0,230,0,98,0,148,0,78,0,0,0,97,0,223,0,159,0,0,0,0,0,60,0,85,0,55,0,41,0,0,0,0,0,0,0,0,0,182,0,79,0,151,0,0,0,161,0,151,0,209,0,43,0,213,0,250,0,0,0,243,0,100,0,88,0,185,0,139,0,34,0,112,0,0,0,188,0,0,0,170,0,179,0,4,0,197,0,141,0,185,0,201,0,43,0,182,0,0,0,0,0,163,0,0,0,199,0,148,0,126,0,194,0,0,0,194,0,14,0,0,0,140,0,68,0,164,0,109,0,0,0,0,0,0,0,2,0,138,0,17,0,0,0,143,0,251,0,47,0,154,0,27,0,253,0,255,0,166,0,180,0,16,0,197,0,241,0,6,0,0,0,81,0,131,0,68,0,51,0,0,0,166,0,173,0,0,0,0,0,111,0,226,0,0,0,18,0,68,0,174,0,163,0,106,0,50,0,124,0,212,0,115,0,44,0,171,0,51,0,218,0,250,0,224,0,0,0,69,0,146,0,0,0,179,0,73,0,0,0,208,0,179,0,0,0,18,0,229,0,162,0,0,0,42,0,126,0,52,0,74,0,214,0,254,0,127,0,201,0,149,0,0,0,0,0,247,0,0,0,174,0,69,0,40,0,57,0,71,0,4,0,0,0,31,0,75,0,58,0,0,0,101,0,90,0,16,0,148,0,0,0,131,0,128,0,234,0,198,0,139,0,69,0,130,0,102,0,0,0,2,0,112,0,43,0,213,0,149,0,160,0,193,0,52,0,149,0,0,0,85,0,194,0,131,0,200,0,190,0,139,0,39,0,0,0,127,0,210,0,0,0,157,0,98,0,227,0,80,0,206,0,0,0,128,0,11,0,37,0,9,0,112,0,139,0,0,0,137,0,21,0,97,0,202,0,109,0,95,0,208,0,132,0,41,0,123,0,31,0,58,0,171,0,78,0,243,0,0,0,28,0,97,0,0,0,18,0,109,0,37,0,214,0,68,0,12,0,234,0,235,0,0,0,118,0,16,0,250,0,0,0,218,0,79,0,172,0,185,0,173,0,130,0,82,0,247,0,0,0,93,0,0,0,0,0,36,0,182,0,92,0,89,0,248,0,37,0,61,0,0,0,27,0,25,0,4,0,153,0,0,0,122,0,30,0,192,0,97,0,0,0,63,0,65,0,46,0,210,0,201,0,120,0,34,0,14,0,185,0,138,0,178,0,0,0,58,0,130,0,255,0,0,0,219,0,179,0,166,0,79,0,179,0,194,0,78,0,164,0,178,0,57,0,58,0,128,0,120,0,120,0,229,0,0,0,16,0,58,0,7,0,85,0,175,0,52,0,38,0,138,0,126,0,205,0,121,0,0,0,143,0,30,0,47,0,0,0,182,0,0,0,199,0,239,0,86,0,0,0,144,0,191,0,0,0,0,0,103,0,13,0,4,0,31,0,178,0,238,0,226,0,0,0,230,0,0,0,69,0,254,0,0,0,22,0,0,0,245,0,185,0,21,0,0,0,10,0,45,0,238,0,41,0,0,0,0,0,140,0,99,0,0,0,132,0,23,0,70,0,237,0,104,0,0,0,0,0,136,0,159,0,115,0,63,0,36,0,235,0,32,0,248,0,105,0,78,0,192,0,0,0,34,0,221,0,160,0,176,0,202,0,210,0,189,0,202,0,222,0,194,0,0,0,215,0,113,0,126,0,167,0,28,0,61,0,138,0,26,0,205,0,0,0,87,0,1,0,31,0,252,0,0,0,0,0,227,0,102,0,247,0,163,0,192,0,0,0,106,0,47,0,144,0,181,0,58,0,92,0,209,0);
signal scenario_full  : scenario_type := (147,31,147,30,114,31,114,30,114,29,70,31,70,30,24,31,24,30,21,31,14,31,187,31,187,30,27,31,111,31,54,31,21,31,74,31,238,31,238,30,76,31,28,31,122,31,185,31,175,31,175,30,19,31,84,31,211,31,160,31,134,31,134,30,17,31,17,30,4,31,86,31,243,31,178,31,152,31,175,31,52,31,118,31,29,31,210,31,118,31,35,31,244,31,244,30,184,31,154,31,35,31,35,30,115,31,115,30,175,31,106,31,191,31,18,31,188,31,112,31,7,31,46,31,121,31,255,31,206,31,76,31,197,31,197,30,53,31,53,30,173,31,173,30,252,31,252,30,133,31,30,31,169,31,101,31,113,31,42,31,228,31,228,30,228,29,52,31,220,31,220,30,246,31,246,30,144,31,70,31,187,31,192,31,228,31,139,31,225,31,13,31,247,31,114,31,18,31,182,31,182,30,61,31,61,30,192,31,43,31,199,31,227,31,86,31,86,30,221,31,193,31,96,31,191,31,54,31,45,31,45,30,7,31,7,30,76,31,76,30,36,31,200,31,200,30,200,29,113,31,250,31,67,31,67,31,178,31,178,30,191,31,25,31,25,30,25,29,43,31,43,30,122,31,203,31,48,31,119,31,248,31,153,31,168,31,168,30,168,29,168,28,71,31,220,31,244,31,59,31,72,31,72,30,160,31,35,31,239,31,239,30,197,31,77,31,77,30,246,31,114,31,203,31,180,31,65,31,177,31,177,30,248,31,64,31,21,31,156,31,209,31,209,30,209,29,35,31,183,31,183,30,183,29,86,31,152,31,191,31,106,31,212,31,159,31,228,31,100,31,100,30,4,31,166,31,166,30,186,31,215,31,184,31,133,31,48,31,246,31,71,31,185,31,5,31,24,31,254,31,68,31,107,31,78,31,134,31,79,31,253,31,198,31,175,31,96,31,148,31,190,31,247,31,111,31,80,31,103,31,178,31,178,30,76,31,76,30,76,29,76,28,96,31,242,31,242,30,242,29,134,31,226,31,119,31,109,31,38,31,126,31,134,31,4,31,206,31,162,31,210,31,248,31,239,31,108,31,209,31,56,31,27,31,189,31,119,31,56,31,53,31,169,31,237,31,89,31,116,31,231,31,231,30,183,31,6,31,213,31,213,30,117,31,181,31,37,31,97,31,97,30,22,31,168,31,90,31,90,30,229,31,136,31,32,31,230,31,98,31,148,31,78,31,78,30,97,31,223,31,159,31,159,30,159,29,60,31,85,31,55,31,41,31,41,30,41,29,41,28,41,27,182,31,79,31,151,31,151,30,161,31,151,31,209,31,43,31,213,31,250,31,250,30,243,31,100,31,88,31,185,31,139,31,34,31,112,31,112,30,188,31,188,30,170,31,179,31,4,31,197,31,141,31,185,31,201,31,43,31,182,31,182,30,182,29,163,31,163,30,199,31,148,31,126,31,194,31,194,30,194,31,14,31,14,30,140,31,68,31,164,31,109,31,109,30,109,29,109,28,2,31,138,31,17,31,17,30,143,31,251,31,47,31,154,31,27,31,253,31,255,31,166,31,180,31,16,31,197,31,241,31,6,31,6,30,81,31,131,31,68,31,51,31,51,30,166,31,173,31,173,30,173,29,111,31,226,31,226,30,18,31,68,31,174,31,163,31,106,31,50,31,124,31,212,31,115,31,44,31,171,31,51,31,218,31,250,31,224,31,224,30,69,31,146,31,146,30,179,31,73,31,73,30,208,31,179,31,179,30,18,31,229,31,162,31,162,30,42,31,126,31,52,31,74,31,214,31,254,31,127,31,201,31,149,31,149,30,149,29,247,31,247,30,174,31,69,31,40,31,57,31,71,31,4,31,4,30,31,31,75,31,58,31,58,30,101,31,90,31,16,31,148,31,148,30,131,31,128,31,234,31,198,31,139,31,69,31,130,31,102,31,102,30,2,31,112,31,43,31,213,31,149,31,160,31,193,31,52,31,149,31,149,30,85,31,194,31,131,31,200,31,190,31,139,31,39,31,39,30,127,31,210,31,210,30,157,31,98,31,227,31,80,31,206,31,206,30,128,31,11,31,37,31,9,31,112,31,139,31,139,30,137,31,21,31,97,31,202,31,109,31,95,31,208,31,132,31,41,31,123,31,31,31,58,31,171,31,78,31,243,31,243,30,28,31,97,31,97,30,18,31,109,31,37,31,214,31,68,31,12,31,234,31,235,31,235,30,118,31,16,31,250,31,250,30,218,31,79,31,172,31,185,31,173,31,130,31,82,31,247,31,247,30,93,31,93,30,93,29,36,31,182,31,92,31,89,31,248,31,37,31,61,31,61,30,27,31,25,31,4,31,153,31,153,30,122,31,30,31,192,31,97,31,97,30,63,31,65,31,46,31,210,31,201,31,120,31,34,31,14,31,185,31,138,31,178,31,178,30,58,31,130,31,255,31,255,30,219,31,179,31,166,31,79,31,179,31,194,31,78,31,164,31,178,31,57,31,58,31,128,31,120,31,120,31,229,31,229,30,16,31,58,31,7,31,85,31,175,31,52,31,38,31,138,31,126,31,205,31,121,31,121,30,143,31,30,31,47,31,47,30,182,31,182,30,199,31,239,31,86,31,86,30,144,31,191,31,191,30,191,29,103,31,13,31,4,31,31,31,178,31,238,31,226,31,226,30,230,31,230,30,69,31,254,31,254,30,22,31,22,30,245,31,185,31,21,31,21,30,10,31,45,31,238,31,41,31,41,30,41,29,140,31,99,31,99,30,132,31,23,31,70,31,237,31,104,31,104,30,104,29,136,31,159,31,115,31,63,31,36,31,235,31,32,31,248,31,105,31,78,31,192,31,192,30,34,31,221,31,160,31,176,31,202,31,210,31,189,31,202,31,222,31,194,31,194,30,215,31,113,31,126,31,167,31,28,31,61,31,138,31,26,31,205,31,205,30,87,31,1,31,31,31,252,31,252,30,252,29,227,31,102,31,247,31,163,31,192,31,192,30,106,31,47,31,144,31,181,31,58,31,92,31,209,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
