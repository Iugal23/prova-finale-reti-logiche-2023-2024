-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_224 is
end project_tb_224;

architecture project_tb_arch_224 of project_tb_224 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 426;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,160,0,48,0,217,0,0,0,47,0,57,0,180,0,86,0,68,0,0,0,169,0,151,0,110,0,0,0,0,0,132,0,234,0,123,0,0,0,0,0,0,0,21,0,217,0,242,0,188,0,5,0,167,0,33,0,71,0,0,0,214,0,253,0,187,0,248,0,0,0,150,0,0,0,86,0,139,0,64,0,172,0,108,0,205,0,226,0,72,0,176,0,201,0,134,0,115,0,212,0,0,0,115,0,198,0,0,0,219,0,168,0,218,0,72,0,210,0,97,0,0,0,164,0,246,0,0,0,0,0,4,0,149,0,98,0,102,0,218,0,13,0,99,0,123,0,28,0,2,0,170,0,211,0,79,0,186,0,220,0,191,0,44,0,55,0,1,0,220,0,230,0,180,0,108,0,7,0,251,0,113,0,64,0,242,0,179,0,115,0,158,0,45,0,155,0,212,0,22,0,122,0,45,0,20,0,0,0,158,0,54,0,0,0,0,0,189,0,173,0,29,0,39,0,87,0,120,0,203,0,75,0,233,0,244,0,154,0,0,0,29,0,131,0,34,0,235,0,225,0,98,0,108,0,65,0,19,0,171,0,204,0,94,0,0,0,18,0,147,0,102,0,171,0,226,0,0,0,0,0,0,0,112,0,199,0,139,0,185,0,104,0,0,0,183,0,2,0,115,0,0,0,133,0,78,0,0,0,128,0,169,0,74,0,135,0,9,0,0,0,114,0,220,0,98,0,35,0,23,0,77,0,111,0,0,0,141,0,47,0,0,0,243,0,18,0,225,0,63,0,168,0,211,0,217,0,138,0,0,0,186,0,37,0,0,0,45,0,215,0,234,0,68,0,182,0,50,0,173,0,65,0,0,0,12,0,22,0,215,0,43,0,62,0,133,0,8,0,183,0,0,0,0,0,0,0,58,0,28,0,182,0,191,0,254,0,61,0,132,0,246,0,160,0,119,0,23,0,24,0,115,0,151,0,37,0,158,0,15,0,211,0,238,0,215,0,213,0,60,0,0,0,153,0,2,0,160,0,191,0,40,0,93,0,0,0,0,0,228,0,140,0,48,0,226,0,73,0,101,0,186,0,247,0,187,0,148,0,63,0,93,0,128,0,84,0,206,0,242,0,220,0,224,0,221,0,48,0,113,0,230,0,244,0,186,0,210,0,0,0,77,0,226,0,0,0,148,0,0,0,163,0,72,0,9,0,211,0,78,0,31,0,0,0,185,0,163,0,173,0,128,0,0,0,11,0,109,0,12,0,49,0,84,0,25,0,0,0,31,0,115,0,175,0,61,0,0,0,94,0,119,0,53,0,106,0,7,0,248,0,137,0,1,0,115,0,249,0,86,0,13,0,5,0,74,0,35,0,245,0,183,0,56,0,122,0,159,0,69,0,47,0,203,0,0,0,169,0,50,0,211,0,0,0,130,0,0,0,0,0,0,0,253,0,10,0,181,0,10,0,181,0,0,0,0,0,0,0,169,0,80,0,0,0,227,0,0,0,0,0,96,0,251,0,255,0,212,0,221,0,2,0,195,0,72,0,0,0,11,0,180,0,218,0,83,0,183,0,254,0,108,0,224,0,0,0,202,0,225,0,236,0,0,0,93,0,168,0,3,0,76,0,185,0,97,0,188,0,184,0,150,0,206,0,171,0,144,0,181,0,224,0,0,0,119,0,248,0,106,0,181,0,92,0,53,0,150,0,177,0,168,0,196,0,149,0,90,0,131,0,0,0,82,0,230,0,245,0,97,0,159,0,173,0,26,0,71,0,56,0,0,0,209,0,226,0,48,0,70,0,0,0,79,0,98,0,149,0,10,0,0,0,186,0,199,0,64,0,154,0,206,0,0,0,228,0,179,0,0,0,117,0,178,0,0,0,243,0,50,0,253,0,176,0,25,0,11,0,0,0);
signal scenario_full  : scenario_type := (0,0,160,31,48,31,217,31,217,30,47,31,57,31,180,31,86,31,68,31,68,30,169,31,151,31,110,31,110,30,110,29,132,31,234,31,123,31,123,30,123,29,123,28,21,31,217,31,242,31,188,31,5,31,167,31,33,31,71,31,71,30,214,31,253,31,187,31,248,31,248,30,150,31,150,30,86,31,139,31,64,31,172,31,108,31,205,31,226,31,72,31,176,31,201,31,134,31,115,31,212,31,212,30,115,31,198,31,198,30,219,31,168,31,218,31,72,31,210,31,97,31,97,30,164,31,246,31,246,30,246,29,4,31,149,31,98,31,102,31,218,31,13,31,99,31,123,31,28,31,2,31,170,31,211,31,79,31,186,31,220,31,191,31,44,31,55,31,1,31,220,31,230,31,180,31,108,31,7,31,251,31,113,31,64,31,242,31,179,31,115,31,158,31,45,31,155,31,212,31,22,31,122,31,45,31,20,31,20,30,158,31,54,31,54,30,54,29,189,31,173,31,29,31,39,31,87,31,120,31,203,31,75,31,233,31,244,31,154,31,154,30,29,31,131,31,34,31,235,31,225,31,98,31,108,31,65,31,19,31,171,31,204,31,94,31,94,30,18,31,147,31,102,31,171,31,226,31,226,30,226,29,226,28,112,31,199,31,139,31,185,31,104,31,104,30,183,31,2,31,115,31,115,30,133,31,78,31,78,30,128,31,169,31,74,31,135,31,9,31,9,30,114,31,220,31,98,31,35,31,23,31,77,31,111,31,111,30,141,31,47,31,47,30,243,31,18,31,225,31,63,31,168,31,211,31,217,31,138,31,138,30,186,31,37,31,37,30,45,31,215,31,234,31,68,31,182,31,50,31,173,31,65,31,65,30,12,31,22,31,215,31,43,31,62,31,133,31,8,31,183,31,183,30,183,29,183,28,58,31,28,31,182,31,191,31,254,31,61,31,132,31,246,31,160,31,119,31,23,31,24,31,115,31,151,31,37,31,158,31,15,31,211,31,238,31,215,31,213,31,60,31,60,30,153,31,2,31,160,31,191,31,40,31,93,31,93,30,93,29,228,31,140,31,48,31,226,31,73,31,101,31,186,31,247,31,187,31,148,31,63,31,93,31,128,31,84,31,206,31,242,31,220,31,224,31,221,31,48,31,113,31,230,31,244,31,186,31,210,31,210,30,77,31,226,31,226,30,148,31,148,30,163,31,72,31,9,31,211,31,78,31,31,31,31,30,185,31,163,31,173,31,128,31,128,30,11,31,109,31,12,31,49,31,84,31,25,31,25,30,31,31,115,31,175,31,61,31,61,30,94,31,119,31,53,31,106,31,7,31,248,31,137,31,1,31,115,31,249,31,86,31,13,31,5,31,74,31,35,31,245,31,183,31,56,31,122,31,159,31,69,31,47,31,203,31,203,30,169,31,50,31,211,31,211,30,130,31,130,30,130,29,130,28,253,31,10,31,181,31,10,31,181,31,181,30,181,29,181,28,169,31,80,31,80,30,227,31,227,30,227,29,96,31,251,31,255,31,212,31,221,31,2,31,195,31,72,31,72,30,11,31,180,31,218,31,83,31,183,31,254,31,108,31,224,31,224,30,202,31,225,31,236,31,236,30,93,31,168,31,3,31,76,31,185,31,97,31,188,31,184,31,150,31,206,31,171,31,144,31,181,31,224,31,224,30,119,31,248,31,106,31,181,31,92,31,53,31,150,31,177,31,168,31,196,31,149,31,90,31,131,31,131,30,82,31,230,31,245,31,97,31,159,31,173,31,26,31,71,31,56,31,56,30,209,31,226,31,48,31,70,31,70,30,79,31,98,31,149,31,10,31,10,30,186,31,199,31,64,31,154,31,206,31,206,30,228,31,179,31,179,30,117,31,178,31,178,30,243,31,50,31,253,31,176,31,25,31,11,31,11,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
