-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 909;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,23,0,125,0,218,0,0,0,142,0,83,0,145,0,0,0,13,0,160,0,241,0,143,0,245,0,183,0,181,0,53,0,0,0,197,0,134,0,150,0,202,0,132,0,137,0,74,0,14,0,170,0,0,0,0,0,123,0,194,0,41,0,153,0,4,0,85,0,110,0,209,0,246,0,242,0,0,0,95,0,229,0,232,0,75,0,177,0,63,0,98,0,0,0,0,0,88,0,152,0,45,0,193,0,118,0,151,0,63,0,60,0,0,0,4,0,0,0,170,0,210,0,0,0,160,0,243,0,16,0,102,0,45,0,0,0,87,0,183,0,209,0,136,0,204,0,10,0,0,0,0,0,113,0,237,0,152,0,204,0,9,0,41,0,205,0,0,0,188,0,70,0,234,0,1,0,69,0,60,0,0,0,163,0,0,0,227,0,11,0,134,0,127,0,84,0,0,0,225,0,244,0,254,0,179,0,2,0,13,0,181,0,190,0,0,0,207,0,33,0,41,0,73,0,36,0,133,0,26,0,57,0,42,0,244,0,221,0,13,0,235,0,100,0,83,0,230,0,138,0,0,0,54,0,48,0,0,0,42,0,52,0,182,0,109,0,236,0,252,0,162,0,175,0,63,0,26,0,20,0,70,0,7,0,0,0,162,0,89,0,112,0,74,0,1,0,173,0,225,0,197,0,31,0,68,0,209,0,176,0,52,0,0,0,181,0,52,0,79,0,59,0,128,0,236,0,195,0,102,0,0,0,105,0,130,0,237,0,0,0,42,0,51,0,180,0,144,0,194,0,139,0,0,0,6,0,0,0,185,0,0,0,73,0,40,0,63,0,93,0,52,0,248,0,230,0,47,0,167,0,239,0,0,0,113,0,124,0,0,0,0,0,0,0,133,0,0,0,71,0,144,0,161,0,0,0,32,0,249,0,0,0,201,0,91,0,199,0,95,0,217,0,231,0,41,0,1,0,184,0,216,0,206,0,0,0,7,0,66,0,99,0,175,0,160,0,44,0,44,0,0,0,8,0,118,0,93,0,121,0,0,0,233,0,57,0,119,0,49,0,233,0,32,0,0,0,52,0,204,0,124,0,131,0,51,0,0,0,205,0,26,0,191,0,89,0,84,0,0,0,115,0,23,0,192,0,0,0,151,0,82,0,162,0,212,0,145,0,100,0,171,0,136,0,105,0,77,0,153,0,9,0,168,0,168,0,237,0,0,0,125,0,0,0,241,0,57,0,235,0,125,0,0,0,14,0,119,0,0,0,249,0,163,0,216,0,62,0,26,0,0,0,51,0,34,0,213,0,0,0,0,0,221,0,253,0,33,0,150,0,133,0,104,0,73,0,29,0,250,0,0,0,183,0,170,0,227,0,138,0,199,0,0,0,74,0,0,0,248,0,59,0,174,0,201,0,0,0,0,0,118,0,110,0,145,0,114,0,85,0,99,0,207,0,89,0,97,0,89,0,88,0,122,0,150,0,152,0,34,0,59,0,91,0,0,0,0,0,193,0,106,0,0,0,164,0,226,0,192,0,54,0,219,0,0,0,211,0,198,0,64,0,3,0,67,0,190,0,0,0,26,0,0,0,79,0,4,0,245,0,144,0,23,0,46,0,59,0,0,0,30,0,210,0,88,0,48,0,0,0,170,0,216,0,223,0,182,0,210,0,226,0,168,0,0,0,157,0,120,0,208,0,63,0,215,0,120,0,253,0,250,0,159,0,44,0,0,0,242,0,237,0,194,0,72,0,188,0,215,0,0,0,0,0,99,0,0,0,0,0,200,0,107,0,0,0,0,0,0,0,121,0,89,0,0,0,0,0,0,0,0,0,196,0,43,0,32,0,158,0,58,0,118,0,99,0,113,0,111,0,180,0,112,0,167,0,0,0,40,0,177,0,223,0,59,0,0,0,46,0,82,0,0,0,128,0,228,0,46,0,27,0,218,0,113,0,0,0,210,0,0,0,106,0,73,0,142,0,216,0,145,0,0,0,164,0,116,0,0,0,13,0,142,0,136,0,140,0,88,0,160,0,159,0,240,0,104,0,209,0,184,0,0,0,169,0,0,0,109,0,143,0,30,0,0,0,186,0,121,0,185,0,0,0,41,0,88,0,189,0,139,0,200,0,7,0,233,0,104,0,0,0,208,0,208,0,0,0,197,0,94,0,0,0,242,0,230,0,0,0,68,0,0,0,0,0,236,0,233,0,201,0,0,0,0,0,146,0,67,0,185,0,0,0,30,0,0,0,162,0,227,0,236,0,0,0,29,0,124,0,209,0,163,0,97,0,8,0,0,0,146,0,152,0,186,0,191,0,72,0,152,0,198,0,169,0,206,0,59,0,23,0,153,0,159,0,0,0,178,0,38,0,86,0,152,0,151,0,14,0,104,0,0,0,45,0,101,0,51,0,69,0,91,0,0,0,180,0,101,0,19,0,0,0,49,0,242,0,0,0,42,0,165,0,235,0,238,0,67,0,150,0,16,0,66,0,0,0,140,0,56,0,36,0,133,0,82,0,184,0,88,0,0,0,0,0,226,0,57,0,173,0,65,0,184,0,0,0,112,0,117,0,151,0,19,0,78,0,0,0,162,0,0,0,178,0,40,0,102,0,238,0,59,0,226,0,26,0,47,0,222,0,43,0,168,0,202,0,92,0,91,0,137,0,209,0,146,0,176,0,0,0,198,0,203,0,222,0,190,0,0,0,55,0,48,0,96,0,234,0,180,0,118,0,234,0,38,0,0,0,214,0,177,0,177,0,146,0,0,0,37,0,139,0,255,0,72,0,0,0,166,0,0,0,244,0,0,0,187,0,0,0,194,0,167,0,35,0,77,0,97,0,0,0,62,0,0,0,169,0,100,0,0,0,0,0,170,0,44,0,196,0,211,0,0,0,219,0,171,0,0,0,0,0,0,0,0,0,248,0,204,0,190,0,9,0,165,0,160,0,232,0,0,0,0,0,61,0,129,0,209,0,0,0,211,0,0,0,101,0,37,0,78,0,0,0,251,0,25,0,79,0,157,0,60,0,5,0,128,0,116,0,222,0,124,0,158,0,185,0,0,0,122,0,221,0,32,0,98,0,0,0,0,0,161,0,207,0,0,0,174,0,109,0,118,0,200,0,0,0,47,0,104,0,103,0,198,0,127,0,0,0,216,0,0,0,111,0,76,0,40,0,247,0,3,0,0,0,188,0,131,0,0,0,0,0,130,0,0,0,197,0,0,0,0,0,255,0,61,0,233,0,223,0,137,0,121,0,114,0,177,0,181,0,0,0,144,0,104,0,242,0,0,0,73,0,64,0,117,0,223,0,0,0,0,0,0,0,0,0,43,0,0,0,209,0,76,0,0,0,122,0,206,0,140,0,106,0,0,0,143,0,48,0,128,0,255,0,0,0,223,0,55,0,5,0,2,0,164,0,146,0,170,0,60,0,201,0,0,0,164,0,152,0,117,0,205,0,101,0,113,0,0,0,83,0,75,0,176,0,128,0,34,0,209,0,87,0,206,0,246,0,135,0,192,0,115,0,145,0,246,0,10,0,179,0,0,0,0,0,6,0,130,0,43,0,0,0,252,0,130,0,209,0,50,0,0,0,123,0,216,0,0,0,216,0,25,0,0,0,68,0,19,0,182,0,217,0,102,0,244,0,63,0,93,0,0,0,222,0,230,0,20,0,3,0,11,0,0,0,147,0,85,0,168,0,0,0,78,0,0,0,0,0,17,0,230,0,45,0,144,0,30,0,254,0,144,0,84,0,0,0,7,0,183,0,169,0,178,0,239,0,68,0,49,0,181,0,21,0,116,0,250,0,126,0,49,0,0,0,0,0,219,0,183,0,109,0,36,0,113,0,202,0,67,0,191,0,133,0,180,0,0,0,0,0,218,0,229,0,212,0,148,0,237,0,0,0,109,0,254,0,40,0,0,0,217,0,0,0,216,0,238,0,15,0,142,0,228,0,33,0,0,0,21,0,26,0,244,0,0,0,117,0,29,0,93,0,170,0,133,0,0,0,6,0,253,0,0,0,124,0,107,0,226,0,189,0,0,0,168,0,249,0,204,0,255,0,149,0,80,0,132,0,175,0);
signal scenario_full  : scenario_type := (0,0,23,31,125,31,218,31,218,30,142,31,83,31,145,31,145,30,13,31,160,31,241,31,143,31,245,31,183,31,181,31,53,31,53,30,197,31,134,31,150,31,202,31,132,31,137,31,74,31,14,31,170,31,170,30,170,29,123,31,194,31,41,31,153,31,4,31,85,31,110,31,209,31,246,31,242,31,242,30,95,31,229,31,232,31,75,31,177,31,63,31,98,31,98,30,98,29,88,31,152,31,45,31,193,31,118,31,151,31,63,31,60,31,60,30,4,31,4,30,170,31,210,31,210,30,160,31,243,31,16,31,102,31,45,31,45,30,87,31,183,31,209,31,136,31,204,31,10,31,10,30,10,29,113,31,237,31,152,31,204,31,9,31,41,31,205,31,205,30,188,31,70,31,234,31,1,31,69,31,60,31,60,30,163,31,163,30,227,31,11,31,134,31,127,31,84,31,84,30,225,31,244,31,254,31,179,31,2,31,13,31,181,31,190,31,190,30,207,31,33,31,41,31,73,31,36,31,133,31,26,31,57,31,42,31,244,31,221,31,13,31,235,31,100,31,83,31,230,31,138,31,138,30,54,31,48,31,48,30,42,31,52,31,182,31,109,31,236,31,252,31,162,31,175,31,63,31,26,31,20,31,70,31,7,31,7,30,162,31,89,31,112,31,74,31,1,31,173,31,225,31,197,31,31,31,68,31,209,31,176,31,52,31,52,30,181,31,52,31,79,31,59,31,128,31,236,31,195,31,102,31,102,30,105,31,130,31,237,31,237,30,42,31,51,31,180,31,144,31,194,31,139,31,139,30,6,31,6,30,185,31,185,30,73,31,40,31,63,31,93,31,52,31,248,31,230,31,47,31,167,31,239,31,239,30,113,31,124,31,124,30,124,29,124,28,133,31,133,30,71,31,144,31,161,31,161,30,32,31,249,31,249,30,201,31,91,31,199,31,95,31,217,31,231,31,41,31,1,31,184,31,216,31,206,31,206,30,7,31,66,31,99,31,175,31,160,31,44,31,44,31,44,30,8,31,118,31,93,31,121,31,121,30,233,31,57,31,119,31,49,31,233,31,32,31,32,30,52,31,204,31,124,31,131,31,51,31,51,30,205,31,26,31,191,31,89,31,84,31,84,30,115,31,23,31,192,31,192,30,151,31,82,31,162,31,212,31,145,31,100,31,171,31,136,31,105,31,77,31,153,31,9,31,168,31,168,31,237,31,237,30,125,31,125,30,241,31,57,31,235,31,125,31,125,30,14,31,119,31,119,30,249,31,163,31,216,31,62,31,26,31,26,30,51,31,34,31,213,31,213,30,213,29,221,31,253,31,33,31,150,31,133,31,104,31,73,31,29,31,250,31,250,30,183,31,170,31,227,31,138,31,199,31,199,30,74,31,74,30,248,31,59,31,174,31,201,31,201,30,201,29,118,31,110,31,145,31,114,31,85,31,99,31,207,31,89,31,97,31,89,31,88,31,122,31,150,31,152,31,34,31,59,31,91,31,91,30,91,29,193,31,106,31,106,30,164,31,226,31,192,31,54,31,219,31,219,30,211,31,198,31,64,31,3,31,67,31,190,31,190,30,26,31,26,30,79,31,4,31,245,31,144,31,23,31,46,31,59,31,59,30,30,31,210,31,88,31,48,31,48,30,170,31,216,31,223,31,182,31,210,31,226,31,168,31,168,30,157,31,120,31,208,31,63,31,215,31,120,31,253,31,250,31,159,31,44,31,44,30,242,31,237,31,194,31,72,31,188,31,215,31,215,30,215,29,99,31,99,30,99,29,200,31,107,31,107,30,107,29,107,28,121,31,89,31,89,30,89,29,89,28,89,27,196,31,43,31,32,31,158,31,58,31,118,31,99,31,113,31,111,31,180,31,112,31,167,31,167,30,40,31,177,31,223,31,59,31,59,30,46,31,82,31,82,30,128,31,228,31,46,31,27,31,218,31,113,31,113,30,210,31,210,30,106,31,73,31,142,31,216,31,145,31,145,30,164,31,116,31,116,30,13,31,142,31,136,31,140,31,88,31,160,31,159,31,240,31,104,31,209,31,184,31,184,30,169,31,169,30,109,31,143,31,30,31,30,30,186,31,121,31,185,31,185,30,41,31,88,31,189,31,139,31,200,31,7,31,233,31,104,31,104,30,208,31,208,31,208,30,197,31,94,31,94,30,242,31,230,31,230,30,68,31,68,30,68,29,236,31,233,31,201,31,201,30,201,29,146,31,67,31,185,31,185,30,30,31,30,30,162,31,227,31,236,31,236,30,29,31,124,31,209,31,163,31,97,31,8,31,8,30,146,31,152,31,186,31,191,31,72,31,152,31,198,31,169,31,206,31,59,31,23,31,153,31,159,31,159,30,178,31,38,31,86,31,152,31,151,31,14,31,104,31,104,30,45,31,101,31,51,31,69,31,91,31,91,30,180,31,101,31,19,31,19,30,49,31,242,31,242,30,42,31,165,31,235,31,238,31,67,31,150,31,16,31,66,31,66,30,140,31,56,31,36,31,133,31,82,31,184,31,88,31,88,30,88,29,226,31,57,31,173,31,65,31,184,31,184,30,112,31,117,31,151,31,19,31,78,31,78,30,162,31,162,30,178,31,40,31,102,31,238,31,59,31,226,31,26,31,47,31,222,31,43,31,168,31,202,31,92,31,91,31,137,31,209,31,146,31,176,31,176,30,198,31,203,31,222,31,190,31,190,30,55,31,48,31,96,31,234,31,180,31,118,31,234,31,38,31,38,30,214,31,177,31,177,31,146,31,146,30,37,31,139,31,255,31,72,31,72,30,166,31,166,30,244,31,244,30,187,31,187,30,194,31,167,31,35,31,77,31,97,31,97,30,62,31,62,30,169,31,100,31,100,30,100,29,170,31,44,31,196,31,211,31,211,30,219,31,171,31,171,30,171,29,171,28,171,27,248,31,204,31,190,31,9,31,165,31,160,31,232,31,232,30,232,29,61,31,129,31,209,31,209,30,211,31,211,30,101,31,37,31,78,31,78,30,251,31,25,31,79,31,157,31,60,31,5,31,128,31,116,31,222,31,124,31,158,31,185,31,185,30,122,31,221,31,32,31,98,31,98,30,98,29,161,31,207,31,207,30,174,31,109,31,118,31,200,31,200,30,47,31,104,31,103,31,198,31,127,31,127,30,216,31,216,30,111,31,76,31,40,31,247,31,3,31,3,30,188,31,131,31,131,30,131,29,130,31,130,30,197,31,197,30,197,29,255,31,61,31,233,31,223,31,137,31,121,31,114,31,177,31,181,31,181,30,144,31,104,31,242,31,242,30,73,31,64,31,117,31,223,31,223,30,223,29,223,28,223,27,43,31,43,30,209,31,76,31,76,30,122,31,206,31,140,31,106,31,106,30,143,31,48,31,128,31,255,31,255,30,223,31,55,31,5,31,2,31,164,31,146,31,170,31,60,31,201,31,201,30,164,31,152,31,117,31,205,31,101,31,113,31,113,30,83,31,75,31,176,31,128,31,34,31,209,31,87,31,206,31,246,31,135,31,192,31,115,31,145,31,246,31,10,31,179,31,179,30,179,29,6,31,130,31,43,31,43,30,252,31,130,31,209,31,50,31,50,30,123,31,216,31,216,30,216,31,25,31,25,30,68,31,19,31,182,31,217,31,102,31,244,31,63,31,93,31,93,30,222,31,230,31,20,31,3,31,11,31,11,30,147,31,85,31,168,31,168,30,78,31,78,30,78,29,17,31,230,31,45,31,144,31,30,31,254,31,144,31,84,31,84,30,7,31,183,31,169,31,178,31,239,31,68,31,49,31,181,31,21,31,116,31,250,31,126,31,49,31,49,30,49,29,219,31,183,31,109,31,36,31,113,31,202,31,67,31,191,31,133,31,180,31,180,30,180,29,218,31,229,31,212,31,148,31,237,31,237,30,109,31,254,31,40,31,40,30,217,31,217,30,216,31,238,31,15,31,142,31,228,31,33,31,33,30,21,31,26,31,244,31,244,30,117,31,29,31,93,31,170,31,133,31,133,30,6,31,253,31,253,30,124,31,107,31,226,31,189,31,189,30,168,31,249,31,204,31,255,31,149,31,80,31,132,31,175,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
