-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 355;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (29,0,124,0,183,0,134,0,1,0,11,0,170,0,0,0,49,0,112,0,26,0,43,0,0,0,189,0,192,0,200,0,0,0,211,0,117,0,83,0,0,0,0,0,100,0,0,0,197,0,245,0,108,0,0,0,179,0,0,0,0,0,152,0,86,0,0,0,72,0,164,0,0,0,33,0,254,0,0,0,176,0,254,0,0,0,181,0,2,0,228,0,0,0,137,0,28,0,33,0,187,0,0,0,24,0,0,0,36,0,140,0,46,0,0,0,237,0,30,0,243,0,197,0,178,0,173,0,207,0,0,0,254,0,0,0,245,0,220,0,244,0,0,0,4,0,0,0,197,0,0,0,219,0,193,0,0,0,71,0,7,0,0,0,237,0,0,0,159,0,0,0,178,0,109,0,248,0,36,0,18,0,241,0,17,0,11,0,0,0,0,0,217,0,79,0,0,0,197,0,0,0,14,0,0,0,19,0,10,0,72,0,205,0,72,0,209,0,6,0,229,0,39,0,211,0,36,0,140,0,198,0,0,0,115,0,183,0,33,0,85,0,158,0,0,0,0,0,123,0,93,0,0,0,18,0,18,0,0,0,125,0,94,0,235,0,150,0,196,0,10,0,37,0,28,0,247,0,9,0,140,0,0,0,0,0,196,0,122,0,42,0,0,0,99,0,250,0,42,0,160,0,113,0,151,0,194,0,0,0,44,0,186,0,250,0,60,0,159,0,238,0,0,0,0,0,53,0,113,0,146,0,56,0,63,0,0,0,128,0,4,0,0,0,150,0,79,0,13,0,188,0,216,0,24,0,244,0,0,0,63,0,55,0,154,0,33,0,254,0,19,0,192,0,242,0,156,0,0,0,169,0,206,0,162,0,137,0,244,0,125,0,176,0,80,0,13,0,107,0,0,0,207,0,196,0,0,0,1,0,0,0,127,0,181,0,145,0,76,0,33,0,151,0,178,0,169,0,183,0,135,0,190,0,126,0,48,0,219,0,233,0,0,0,149,0,63,0,221,0,53,0,250,0,246,0,0,0,83,0,0,0,152,0,216,0,26,0,192,0,220,0,97,0,150,0,130,0,234,0,152,0,253,0,57,0,0,0,211,0,115,0,236,0,45,0,225,0,41,0,115,0,252,0,128,0,184,0,187,0,249,0,189,0,79,0,224,0,75,0,52,0,6,0,246,0,127,0,0,0,131,0,0,0,22,0,217,0,148,0,0,0,8,0,206,0,119,0,52,0,189,0,8,0,0,0,252,0,152,0,209,0,224,0,109,0,0,0,0,0,75,0,0,0,32,0,189,0,37,0,0,0,0,0,12,0,133,0,134,0,0,0,180,0,15,0,58,0,4,0,143,0,18,0,41,0,20,0,198,0,233,0,235,0,0,0,86,0,0,0,0,0,121,0,0,0,64,0,16,0,194,0,202,0,0,0,0,0,226,0,31,0,99,0,73,0,0,0,41,0,136,0,22,0,5,0,44,0,139,0,30,0,194,0,0,0,0,0,0,0,0,0,192,0,0,0,9,0,171,0,207,0,123,0,40,0,197,0,0,0,0,0,173,0,0,0,214,0,133,0,0,0,232,0,166,0,210,0,130,0);
signal scenario_full  : scenario_type := (29,31,124,31,183,31,134,31,1,31,11,31,170,31,170,30,49,31,112,31,26,31,43,31,43,30,189,31,192,31,200,31,200,30,211,31,117,31,83,31,83,30,83,29,100,31,100,30,197,31,245,31,108,31,108,30,179,31,179,30,179,29,152,31,86,31,86,30,72,31,164,31,164,30,33,31,254,31,254,30,176,31,254,31,254,30,181,31,2,31,228,31,228,30,137,31,28,31,33,31,187,31,187,30,24,31,24,30,36,31,140,31,46,31,46,30,237,31,30,31,243,31,197,31,178,31,173,31,207,31,207,30,254,31,254,30,245,31,220,31,244,31,244,30,4,31,4,30,197,31,197,30,219,31,193,31,193,30,71,31,7,31,7,30,237,31,237,30,159,31,159,30,178,31,109,31,248,31,36,31,18,31,241,31,17,31,11,31,11,30,11,29,217,31,79,31,79,30,197,31,197,30,14,31,14,30,19,31,10,31,72,31,205,31,72,31,209,31,6,31,229,31,39,31,211,31,36,31,140,31,198,31,198,30,115,31,183,31,33,31,85,31,158,31,158,30,158,29,123,31,93,31,93,30,18,31,18,31,18,30,125,31,94,31,235,31,150,31,196,31,10,31,37,31,28,31,247,31,9,31,140,31,140,30,140,29,196,31,122,31,42,31,42,30,99,31,250,31,42,31,160,31,113,31,151,31,194,31,194,30,44,31,186,31,250,31,60,31,159,31,238,31,238,30,238,29,53,31,113,31,146,31,56,31,63,31,63,30,128,31,4,31,4,30,150,31,79,31,13,31,188,31,216,31,24,31,244,31,244,30,63,31,55,31,154,31,33,31,254,31,19,31,192,31,242,31,156,31,156,30,169,31,206,31,162,31,137,31,244,31,125,31,176,31,80,31,13,31,107,31,107,30,207,31,196,31,196,30,1,31,1,30,127,31,181,31,145,31,76,31,33,31,151,31,178,31,169,31,183,31,135,31,190,31,126,31,48,31,219,31,233,31,233,30,149,31,63,31,221,31,53,31,250,31,246,31,246,30,83,31,83,30,152,31,216,31,26,31,192,31,220,31,97,31,150,31,130,31,234,31,152,31,253,31,57,31,57,30,211,31,115,31,236,31,45,31,225,31,41,31,115,31,252,31,128,31,184,31,187,31,249,31,189,31,79,31,224,31,75,31,52,31,6,31,246,31,127,31,127,30,131,31,131,30,22,31,217,31,148,31,148,30,8,31,206,31,119,31,52,31,189,31,8,31,8,30,252,31,152,31,209,31,224,31,109,31,109,30,109,29,75,31,75,30,32,31,189,31,37,31,37,30,37,29,12,31,133,31,134,31,134,30,180,31,15,31,58,31,4,31,143,31,18,31,41,31,20,31,198,31,233,31,235,31,235,30,86,31,86,30,86,29,121,31,121,30,64,31,16,31,194,31,202,31,202,30,202,29,226,31,31,31,99,31,73,31,73,30,41,31,136,31,22,31,5,31,44,31,139,31,30,31,194,31,194,30,194,29,194,28,194,27,192,31,192,30,9,31,171,31,207,31,123,31,40,31,197,31,197,30,197,29,173,31,173,30,214,31,133,31,133,30,232,31,166,31,210,31,130,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
