-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 999;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (210,0,224,0,241,0,23,0,204,0,0,0,162,0,44,0,17,0,174,0,53,0,81,0,15,0,227,0,0,0,45,0,106,0,150,0,184,0,127,0,179,0,142,0,40,0,247,0,31,0,39,0,214,0,118,0,2,0,19,0,244,0,0,0,241,0,18,0,211,0,48,0,158,0,33,0,249,0,8,0,34,0,84,0,0,0,19,0,177,0,0,0,61,0,88,0,229,0,248,0,0,0,39,0,30,0,114,0,232,0,0,0,0,0,221,0,135,0,2,0,0,0,0,0,192,0,149,0,17,0,37,0,58,0,33,0,50,0,100,0,144,0,0,0,0,0,0,0,252,0,65,0,13,0,124,0,176,0,15,0,132,0,0,0,176,0,251,0,177,0,72,0,51,0,241,0,73,0,197,0,77,0,131,0,45,0,33,0,0,0,83,0,251,0,0,0,0,0,0,0,149,0,108,0,76,0,190,0,0,0,99,0,120,0,126,0,198,0,152,0,38,0,204,0,109,0,141,0,0,0,0,0,40,0,0,0,102,0,145,0,0,0,39,0,169,0,93,0,250,0,144,0,2,0,0,0,174,0,167,0,180,0,187,0,99,0,63,0,40,0,41,0,35,0,201,0,170,0,55,0,167,0,79,0,62,0,249,0,213,0,222,0,80,0,123,0,98,0,163,0,110,0,0,0,85,0,21,0,118,0,193,0,0,0,9,0,161,0,119,0,177,0,0,0,43,0,41,0,87,0,234,0,94,0,244,0,20,0,231,0,16,0,215,0,0,0,107,0,0,0,0,0,175,0,174,0,84,0,10,0,0,0,255,0,0,0,247,0,7,0,72,0,14,0,46,0,195,0,110,0,157,0,86,0,25,0,244,0,250,0,171,0,3,0,225,0,231,0,199,0,189,0,147,0,95,0,0,0,14,0,60,0,50,0,208,0,246,0,160,0,19,0,223,0,215,0,219,0,78,0,0,0,32,0,72,0,1,0,0,0,0,0,79,0,35,0,181,0,118,0,51,0,194,0,163,0,149,0,28,0,223,0,78,0,138,0,141,0,29,0,0,0,140,0,68,0,238,0,0,0,191,0,222,0,197,0,64,0,200,0,56,0,225,0,0,0,0,0,0,0,132,0,93,0,0,0,44,0,8,0,0,0,1,0,0,0,12,0,0,0,249,0,212,0,187,0,80,0,122,0,109,0,221,0,228,0,203,0,162,0,13,0,94,0,48,0,15,0,45,0,97,0,198,0,169,0,0,0,228,0,119,0,45,0,244,0,123,0,60,0,154,0,146,0,0,0,31,0,0,0,102,0,199,0,120,0,103,0,93,0,0,0,0,0,0,0,59,0,33,0,234,0,57,0,0,0,8,0,209,0,42,0,213,0,0,0,103,0,0,0,0,0,37,0,7,0,106,0,109,0,68,0,198,0,221,0,169,0,123,0,94,0,134,0,0,0,58,0,55,0,111,0,73,0,254,0,220,0,26,0,30,0,238,0,107,0,0,0,175,0,43,0,4,0,0,0,85,0,0,0,103,0,53,0,213,0,141,0,0,0,43,0,236,0,0,0,144,0,92,0,104,0,84,0,64,0,141,0,196,0,233,0,190,0,250,0,190,0,148,0,80,0,208,0,31,0,173,0,243,0,202,0,0,0,193,0,136,0,0,0,168,0,0,0,50,0,0,0,111,0,0,0,212,0,75,0,49,0,162,0,97,0,96,0,133,0,156,0,126,0,0,0,71,0,110,0,254,0,190,0,222,0,97,0,199,0,123,0,133,0,130,0,59,0,132,0,185,0,0,0,228,0,172,0,25,0,78,0,166,0,93,0,5,0,185,0,44,0,196,0,232,0,59,0,92,0,15,0,9,0,0,0,0,0,0,0,233,0,0,0,0,0,0,0,66,0,44,0,201,0,198,0,166,0,0,0,21,0,26,0,0,0,200,0,59,0,0,0,201,0,0,0,176,0,0,0,3,0,121,0,0,0,0,0,249,0,172,0,0,0,7,0,11,0,220,0,32,0,248,0,0,0,253,0,0,0,75,0,70,0,119,0,63,0,71,0,0,0,17,0,20,0,252,0,218,0,0,0,0,0,111,0,0,0,7,0,216,0,13,0,0,0,247,0,219,0,170,0,0,0,120,0,0,0,44,0,0,0,0,0,223,0,24,0,156,0,66,0,177,0,216,0,241,0,222,0,46,0,138,0,127,0,108,0,234,0,0,0,75,0,190,0,85,0,253,0,173,0,9,0,0,0,4,0,199,0,164,0,155,0,148,0,146,0,105,0,215,0,48,0,172,0,251,0,119,0,150,0,146,0,73,0,35,0,0,0,248,0,0,0,0,0,0,0,195,0,213,0,0,0,0,0,251,0,221,0,23,0,161,0,0,0,77,0,226,0,8,0,3,0,0,0,184,0,137,0,252,0,67,0,142,0,118,0,8,0,41,0,242,0,225,0,160,0,38,0,76,0,64,0,0,0,128,0,124,0,209,0,162,0,149,0,176,0,8,0,11,0,199,0,223,0,122,0,140,0,0,0,70,0,196,0,0,0,44,0,4,0,0,0,0,0,10,0,243,0,24,0,208,0,232,0,237,0,63,0,11,0,232,0,118,0,52,0,106,0,0,0,206,0,170,0,0,0,0,0,116,0,156,0,144,0,69,0,216,0,89,0,32,0,0,0,0,0,69,0,85,0,0,0,0,0,177,0,0,0,174,0,194,0,191,0,196,0,220,0,0,0,0,0,33,0,103,0,202,0,178,0,0,0,0,0,111,0,188,0,194,0,43,0,59,0,87,0,189,0,150,0,43,0,0,0,185,0,95,0,233,0,184,0,57,0,9,0,72,0,153,0,109,0,127,0,43,0,140,0,0,0,182,0,185,0,108,0,142,0,175,0,37,0,66,0,203,0,0,0,53,0,0,0,22,0,156,0,0,0,137,0,92,0,186,0,150,0,216,0,229,0,94,0,171,0,0,0,6,0,138,0,107,0,112,0,0,0,0,0,252,0,142,0,108,0,235,0,131,0,199,0,225,0,0,0,77,0,152,0,16,0,198,0,159,0,87,0,21,0,0,0,114,0,102,0,178,0,185,0,154,0,0,0,69,0,141,0,15,0,125,0,121,0,0,0,104,0,230,0,0,0,136,0,216,0,0,0,173,0,0,0,144,0,150,0,51,0,107,0,0,0,202,0,0,0,0,0,0,0,255,0,177,0,16,0,231,0,0,0,0,0,203,0,0,0,187,0,213,0,142,0,0,0,0,0,125,0,221,0,43,0,98,0,130,0,0,0,28,0,10,0,0,0,148,0,169,0,175,0,0,0,9,0,69,0,194,0,51,0,0,0,39,0,110,0,231,0,0,0,110,0,108,0,145,0,96,0,0,0,22,0,0,0,0,0,187,0,92,0,175,0,0,0,246,0,19,0,96,0,0,0,239,0,60,0,226,0,173,0,76,0,0,0,104,0,119,0,0,0,91,0,14,0,0,0,97,0,0,0,77,0,242,0,121,0,98,0,54,0,0,0,59,0,48,0,192,0,95,0,45,0,55,0,0,0,55,0,0,0,0,0,94,0,197,0,0,0,148,0,48,0,141,0,95,0,224,0,120,0,0,0,46,0,0,0,45,0,193,0,103,0,147,0,138,0,208,0,152,0,3,0,58,0,0,0,18,0,0,0,179,0,0,0,223,0,34,0,23,0,12,0,71,0,174,0,134,0,23,0,226,0,244,0,222,0,9,0,0,0,62,0,102,0,176,0,0,0,43,0,122,0,14,0,138,0,114,0,163,0,0,0,168,0,0,0,158,0,126,0,246,0,28,0,82,0,22,0,74,0,116,0,0,0,251,0,199,0,212,0,13,0,74,0,52,0,206,0,0,0,0,0,193,0,0,0,0,0,144,0,48,0,195,0,76,0,13,0,115,0,42,0,30,0,97,0,85,0,50,0,1,0,141,0,64,0,138,0,4,0,41,0,215,0,76,0,0,0,0,0,110,0,251,0,0,0,0,0,250,0,128,0,223,0,38,0,0,0,142,0,37,0,224,0,62,0,207,0,0,0,29,0,122,0,165,0,147,0,247,0,96,0,178,0,0,0,75,0,213,0,0,0,53,0,138,0,0,0,13,0,62,0,169,0,237,0,108,0,152,0,224,0,0,0,0,0,0,0,97,0,67,0,201,0,0,0,164,0,24,0,229,0,174,0,217,0,29,0,216,0,0,0,158,0,212,0,45,0,0,0,92,0,178,0,252,0,106,0,49,0,0,0,0,0,60,0,45,0,25,0,66,0,188,0,84,0,127,0,0,0,132,0,45,0,92,0,12,0,120,0,0,0,179,0,0,0,233,0,177,0,126,0,191,0,11,0,212,0,154,0,73,0,102,0,0,0,183,0,231,0,22,0,49,0,63,0,76,0,44,0,0,0,33,0,223,0,20,0,0,0,145,0,0,0,238,0,141,0,4,0,163,0,0,0,243,0,99,0,217,0,126,0);
signal scenario_full  : scenario_type := (210,31,224,31,241,31,23,31,204,31,204,30,162,31,44,31,17,31,174,31,53,31,81,31,15,31,227,31,227,30,45,31,106,31,150,31,184,31,127,31,179,31,142,31,40,31,247,31,31,31,39,31,214,31,118,31,2,31,19,31,244,31,244,30,241,31,18,31,211,31,48,31,158,31,33,31,249,31,8,31,34,31,84,31,84,30,19,31,177,31,177,30,61,31,88,31,229,31,248,31,248,30,39,31,30,31,114,31,232,31,232,30,232,29,221,31,135,31,2,31,2,30,2,29,192,31,149,31,17,31,37,31,58,31,33,31,50,31,100,31,144,31,144,30,144,29,144,28,252,31,65,31,13,31,124,31,176,31,15,31,132,31,132,30,176,31,251,31,177,31,72,31,51,31,241,31,73,31,197,31,77,31,131,31,45,31,33,31,33,30,83,31,251,31,251,30,251,29,251,28,149,31,108,31,76,31,190,31,190,30,99,31,120,31,126,31,198,31,152,31,38,31,204,31,109,31,141,31,141,30,141,29,40,31,40,30,102,31,145,31,145,30,39,31,169,31,93,31,250,31,144,31,2,31,2,30,174,31,167,31,180,31,187,31,99,31,63,31,40,31,41,31,35,31,201,31,170,31,55,31,167,31,79,31,62,31,249,31,213,31,222,31,80,31,123,31,98,31,163,31,110,31,110,30,85,31,21,31,118,31,193,31,193,30,9,31,161,31,119,31,177,31,177,30,43,31,41,31,87,31,234,31,94,31,244,31,20,31,231,31,16,31,215,31,215,30,107,31,107,30,107,29,175,31,174,31,84,31,10,31,10,30,255,31,255,30,247,31,7,31,72,31,14,31,46,31,195,31,110,31,157,31,86,31,25,31,244,31,250,31,171,31,3,31,225,31,231,31,199,31,189,31,147,31,95,31,95,30,14,31,60,31,50,31,208,31,246,31,160,31,19,31,223,31,215,31,219,31,78,31,78,30,32,31,72,31,1,31,1,30,1,29,79,31,35,31,181,31,118,31,51,31,194,31,163,31,149,31,28,31,223,31,78,31,138,31,141,31,29,31,29,30,140,31,68,31,238,31,238,30,191,31,222,31,197,31,64,31,200,31,56,31,225,31,225,30,225,29,225,28,132,31,93,31,93,30,44,31,8,31,8,30,1,31,1,30,12,31,12,30,249,31,212,31,187,31,80,31,122,31,109,31,221,31,228,31,203,31,162,31,13,31,94,31,48,31,15,31,45,31,97,31,198,31,169,31,169,30,228,31,119,31,45,31,244,31,123,31,60,31,154,31,146,31,146,30,31,31,31,30,102,31,199,31,120,31,103,31,93,31,93,30,93,29,93,28,59,31,33,31,234,31,57,31,57,30,8,31,209,31,42,31,213,31,213,30,103,31,103,30,103,29,37,31,7,31,106,31,109,31,68,31,198,31,221,31,169,31,123,31,94,31,134,31,134,30,58,31,55,31,111,31,73,31,254,31,220,31,26,31,30,31,238,31,107,31,107,30,175,31,43,31,4,31,4,30,85,31,85,30,103,31,53,31,213,31,141,31,141,30,43,31,236,31,236,30,144,31,92,31,104,31,84,31,64,31,141,31,196,31,233,31,190,31,250,31,190,31,148,31,80,31,208,31,31,31,173,31,243,31,202,31,202,30,193,31,136,31,136,30,168,31,168,30,50,31,50,30,111,31,111,30,212,31,75,31,49,31,162,31,97,31,96,31,133,31,156,31,126,31,126,30,71,31,110,31,254,31,190,31,222,31,97,31,199,31,123,31,133,31,130,31,59,31,132,31,185,31,185,30,228,31,172,31,25,31,78,31,166,31,93,31,5,31,185,31,44,31,196,31,232,31,59,31,92,31,15,31,9,31,9,30,9,29,9,28,233,31,233,30,233,29,233,28,66,31,44,31,201,31,198,31,166,31,166,30,21,31,26,31,26,30,200,31,59,31,59,30,201,31,201,30,176,31,176,30,3,31,121,31,121,30,121,29,249,31,172,31,172,30,7,31,11,31,220,31,32,31,248,31,248,30,253,31,253,30,75,31,70,31,119,31,63,31,71,31,71,30,17,31,20,31,252,31,218,31,218,30,218,29,111,31,111,30,7,31,216,31,13,31,13,30,247,31,219,31,170,31,170,30,120,31,120,30,44,31,44,30,44,29,223,31,24,31,156,31,66,31,177,31,216,31,241,31,222,31,46,31,138,31,127,31,108,31,234,31,234,30,75,31,190,31,85,31,253,31,173,31,9,31,9,30,4,31,199,31,164,31,155,31,148,31,146,31,105,31,215,31,48,31,172,31,251,31,119,31,150,31,146,31,73,31,35,31,35,30,248,31,248,30,248,29,248,28,195,31,213,31,213,30,213,29,251,31,221,31,23,31,161,31,161,30,77,31,226,31,8,31,3,31,3,30,184,31,137,31,252,31,67,31,142,31,118,31,8,31,41,31,242,31,225,31,160,31,38,31,76,31,64,31,64,30,128,31,124,31,209,31,162,31,149,31,176,31,8,31,11,31,199,31,223,31,122,31,140,31,140,30,70,31,196,31,196,30,44,31,4,31,4,30,4,29,10,31,243,31,24,31,208,31,232,31,237,31,63,31,11,31,232,31,118,31,52,31,106,31,106,30,206,31,170,31,170,30,170,29,116,31,156,31,144,31,69,31,216,31,89,31,32,31,32,30,32,29,69,31,85,31,85,30,85,29,177,31,177,30,174,31,194,31,191,31,196,31,220,31,220,30,220,29,33,31,103,31,202,31,178,31,178,30,178,29,111,31,188,31,194,31,43,31,59,31,87,31,189,31,150,31,43,31,43,30,185,31,95,31,233,31,184,31,57,31,9,31,72,31,153,31,109,31,127,31,43,31,140,31,140,30,182,31,185,31,108,31,142,31,175,31,37,31,66,31,203,31,203,30,53,31,53,30,22,31,156,31,156,30,137,31,92,31,186,31,150,31,216,31,229,31,94,31,171,31,171,30,6,31,138,31,107,31,112,31,112,30,112,29,252,31,142,31,108,31,235,31,131,31,199,31,225,31,225,30,77,31,152,31,16,31,198,31,159,31,87,31,21,31,21,30,114,31,102,31,178,31,185,31,154,31,154,30,69,31,141,31,15,31,125,31,121,31,121,30,104,31,230,31,230,30,136,31,216,31,216,30,173,31,173,30,144,31,150,31,51,31,107,31,107,30,202,31,202,30,202,29,202,28,255,31,177,31,16,31,231,31,231,30,231,29,203,31,203,30,187,31,213,31,142,31,142,30,142,29,125,31,221,31,43,31,98,31,130,31,130,30,28,31,10,31,10,30,148,31,169,31,175,31,175,30,9,31,69,31,194,31,51,31,51,30,39,31,110,31,231,31,231,30,110,31,108,31,145,31,96,31,96,30,22,31,22,30,22,29,187,31,92,31,175,31,175,30,246,31,19,31,96,31,96,30,239,31,60,31,226,31,173,31,76,31,76,30,104,31,119,31,119,30,91,31,14,31,14,30,97,31,97,30,77,31,242,31,121,31,98,31,54,31,54,30,59,31,48,31,192,31,95,31,45,31,55,31,55,30,55,31,55,30,55,29,94,31,197,31,197,30,148,31,48,31,141,31,95,31,224,31,120,31,120,30,46,31,46,30,45,31,193,31,103,31,147,31,138,31,208,31,152,31,3,31,58,31,58,30,18,31,18,30,179,31,179,30,223,31,34,31,23,31,12,31,71,31,174,31,134,31,23,31,226,31,244,31,222,31,9,31,9,30,62,31,102,31,176,31,176,30,43,31,122,31,14,31,138,31,114,31,163,31,163,30,168,31,168,30,158,31,126,31,246,31,28,31,82,31,22,31,74,31,116,31,116,30,251,31,199,31,212,31,13,31,74,31,52,31,206,31,206,30,206,29,193,31,193,30,193,29,144,31,48,31,195,31,76,31,13,31,115,31,42,31,30,31,97,31,85,31,50,31,1,31,141,31,64,31,138,31,4,31,41,31,215,31,76,31,76,30,76,29,110,31,251,31,251,30,251,29,250,31,128,31,223,31,38,31,38,30,142,31,37,31,224,31,62,31,207,31,207,30,29,31,122,31,165,31,147,31,247,31,96,31,178,31,178,30,75,31,213,31,213,30,53,31,138,31,138,30,13,31,62,31,169,31,237,31,108,31,152,31,224,31,224,30,224,29,224,28,97,31,67,31,201,31,201,30,164,31,24,31,229,31,174,31,217,31,29,31,216,31,216,30,158,31,212,31,45,31,45,30,92,31,178,31,252,31,106,31,49,31,49,30,49,29,60,31,45,31,25,31,66,31,188,31,84,31,127,31,127,30,132,31,45,31,92,31,12,31,120,31,120,30,179,31,179,30,233,31,177,31,126,31,191,31,11,31,212,31,154,31,73,31,102,31,102,30,183,31,231,31,22,31,49,31,63,31,76,31,44,31,44,30,33,31,223,31,20,31,20,30,145,31,145,30,238,31,141,31,4,31,163,31,163,30,243,31,99,31,217,31,126,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
