-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 204;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (144,0,0,0,209,0,83,0,182,0,114,0,195,0,0,0,0,0,55,0,147,0,126,0,0,0,39,0,141,0,16,0,219,0,27,0,46,0,215,0,7,0,116,0,73,0,175,0,159,0,232,0,235,0,0,0,74,0,57,0,47,0,0,0,138,0,0,0,85,0,0,0,206,0,175,0,0,0,27,0,0,0,147,0,169,0,154,0,203,0,31,0,78,0,211,0,0,0,170,0,225,0,69,0,33,0,66,0,112,0,65,0,68,0,0,0,216,0,0,0,213,0,239,0,0,0,237,0,46,0,0,0,191,0,54,0,103,0,78,0,31,0,54,0,143,0,25,0,135,0,220,0,13,0,79,0,47,0,200,0,0,0,93,0,0,0,120,0,151,0,12,0,82,0,116,0,0,0,192,0,0,0,0,0,54,0,0,0,141,0,184,0,167,0,0,0,0,0,0,0,0,0,94,0,63,0,45,0,20,0,1,0,0,0,30,0,26,0,7,0,35,0,46,0,113,0,241,0,253,0,0,0,0,0,166,0,240,0,247,0,47,0,233,0,38,0,156,0,81,0,127,0,0,0,58,0,4,0,169,0,142,0,83,0,181,0,7,0,45,0,0,0,30,0,90,0,220,0,163,0,0,0,139,0,0,0,88,0,228,0,35,0,191,0,88,0,233,0,0,0,61,0,74,0,0,0,59,0,46,0,78,0,88,0,15,0,146,0,0,0,123,0,244,0,120,0,198,0,200,0,4,0,0,0,22,0,55,0,0,0,112,0,209,0,174,0,224,0,93,0,0,0,155,0,124,0,85,0,144,0,31,0,71,0,64,0,3,0,3,0,124,0,104,0,98,0,0,0,145,0,0,0,91,0,83,0,160,0,61,0,106,0,59,0,13,0,83,0,0,0,101,0,166,0,65,0,226,0);
signal scenario_full  : scenario_type := (144,31,144,30,209,31,83,31,182,31,114,31,195,31,195,30,195,29,55,31,147,31,126,31,126,30,39,31,141,31,16,31,219,31,27,31,46,31,215,31,7,31,116,31,73,31,175,31,159,31,232,31,235,31,235,30,74,31,57,31,47,31,47,30,138,31,138,30,85,31,85,30,206,31,175,31,175,30,27,31,27,30,147,31,169,31,154,31,203,31,31,31,78,31,211,31,211,30,170,31,225,31,69,31,33,31,66,31,112,31,65,31,68,31,68,30,216,31,216,30,213,31,239,31,239,30,237,31,46,31,46,30,191,31,54,31,103,31,78,31,31,31,54,31,143,31,25,31,135,31,220,31,13,31,79,31,47,31,200,31,200,30,93,31,93,30,120,31,151,31,12,31,82,31,116,31,116,30,192,31,192,30,192,29,54,31,54,30,141,31,184,31,167,31,167,30,167,29,167,28,167,27,94,31,63,31,45,31,20,31,1,31,1,30,30,31,26,31,7,31,35,31,46,31,113,31,241,31,253,31,253,30,253,29,166,31,240,31,247,31,47,31,233,31,38,31,156,31,81,31,127,31,127,30,58,31,4,31,169,31,142,31,83,31,181,31,7,31,45,31,45,30,30,31,90,31,220,31,163,31,163,30,139,31,139,30,88,31,228,31,35,31,191,31,88,31,233,31,233,30,61,31,74,31,74,30,59,31,46,31,78,31,88,31,15,31,146,31,146,30,123,31,244,31,120,31,198,31,200,31,4,31,4,30,22,31,55,31,55,30,112,31,209,31,174,31,224,31,93,31,93,30,155,31,124,31,85,31,144,31,31,31,71,31,64,31,3,31,3,31,124,31,104,31,98,31,98,30,145,31,145,30,91,31,83,31,160,31,61,31,106,31,59,31,13,31,83,31,83,30,101,31,166,31,65,31,226,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
