-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 974;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (2,0,117,0,230,0,215,0,112,0,17,0,122,0,0,0,104,0,239,0,46,0,12,0,74,0,22,0,156,0,52,0,0,0,67,0,246,0,45,0,6,0,66,0,0,0,62,0,0,0,51,0,144,0,0,0,105,0,0,0,0,0,231,0,67,0,57,0,247,0,242,0,0,0,29,0,232,0,140,0,0,0,0,0,60,0,68,0,223,0,162,0,0,0,244,0,0,0,108,0,0,0,233,0,231,0,3,0,179,0,139,0,64,0,0,0,233,0,96,0,68,0,190,0,0,0,132,0,59,0,47,0,236,0,242,0,162,0,0,0,182,0,57,0,179,0,0,0,0,0,224,0,0,0,171,0,0,0,9,0,237,0,0,0,0,0,129,0,0,0,4,0,163,0,183,0,182,0,0,0,215,0,34,0,215,0,0,0,18,0,133,0,0,0,134,0,103,0,240,0,220,0,223,0,225,0,210,0,207,0,70,0,0,0,0,0,130,0,147,0,0,0,154,0,137,0,13,0,176,0,121,0,221,0,170,0,145,0,237,0,212,0,0,0,97,0,239,0,229,0,198,0,239,0,0,0,101,0,107,0,236,0,44,0,123,0,110,0,0,0,0,0,254,0,202,0,104,0,156,0,0,0,0,0,25,0,52,0,0,0,31,0,227,0,90,0,93,0,9,0,190,0,84,0,254,0,0,0,225,0,157,0,58,0,0,0,228,0,137,0,26,0,0,0,31,0,0,0,0,0,190,0,250,0,96,0,26,0,45,0,62,0,171,0,76,0,65,0,0,0,0,0,245,0,100,0,19,0,80,0,190,0,14,0,148,0,228,0,19,0,85,0,208,0,0,0,211,0,241,0,0,0,111,0,150,0,65,0,97,0,118,0,135,0,241,0,123,0,217,0,229,0,145,0,162,0,247,0,51,0,0,0,0,0,0,0,114,0,147,0,213,0,178,0,218,0,17,0,66,0,80,0,211,0,252,0,107,0,232,0,58,0,254,0,108,0,133,0,79,0,211,0,80,0,0,0,197,0,39,0,167,0,53,0,125,0,28,0,41,0,96,0,130,0,246,0,83,0,93,0,150,0,134,0,26,0,33,0,95,0,90,0,39,0,221,0,159,0,103,0,42,0,212,0,207,0,0,0,0,0,0,0,0,0,226,0,6,0,246,0,110,0,240,0,0,0,0,0,84,0,129,0,102,0,36,0,0,0,24,0,38,0,101,0,0,0,0,0,187,0,30,0,207,0,102,0,172,0,101,0,120,0,104,0,0,0,212,0,31,0,0,0,177,0,237,0,208,0,0,0,111,0,174,0,51,0,0,0,49,0,69,0,0,0,224,0,213,0,99,0,199,0,239,0,242,0,54,0,0,0,191,0,0,0,145,0,220,0,186,0,68,0,40,0,163,0,0,0,213,0,118,0,93,0,0,0,232,0,185,0,167,0,46,0,183,0,160,0,61,0,159,0,252,0,139,0,245,0,176,0,0,0,167,0,0,0,97,0,0,0,0,0,166,0,0,0,100,0,241,0,0,0,170,0,149,0,162,0,195,0,101,0,222,0,121,0,171,0,239,0,215,0,88,0,191,0,48,0,98,0,177,0,0,0,47,0,174,0,95,0,164,0,144,0,164,0,140,0,29,0,0,0,225,0,109,0,210,0,19,0,184,0,112,0,218,0,66,0,247,0,237,0,243,0,158,0,171,0,4,0,40,0,79,0,0,0,177,0,123,0,0,0,194,0,245,0,6,0,0,0,140,0,0,0,127,0,36,0,2,0,182,0,196,0,0,0,25,0,0,0,0,0,138,0,9,0,116,0,123,0,37,0,85,0,194,0,0,0,0,0,50,0,19,0,0,0,180,0,0,0,158,0,5,0,113,0,130,0,3,0,40,0,130,0,41,0,3,0,0,0,134,0,220,0,0,0,232,0,57,0,0,0,0,0,74,0,200,0,168,0,0,0,175,0,63,0,0,0,91,0,0,0,165,0,255,0,69,0,240,0,223,0,69,0,96,0,0,0,0,0,0,0,136,0,128,0,23,0,11,0,240,0,88,0,156,0,144,0,53,0,52,0,152,0,110,0,184,0,168,0,186,0,76,0,218,0,62,0,148,0,126,0,206,0,177,0,117,0,157,0,254,0,152,0,241,0,58,0,0,0,66,0,36,0,140,0,66,0,146,0,245,0,170,0,0,0,0,0,0,0,9,0,102,0,76,0,67,0,0,0,65,0,187,0,0,0,64,0,57,0,183,0,87,0,12,0,245,0,228,0,34,0,67,0,0,0,0,0,59,0,0,0,0,0,0,0,57,0,125,0,0,0,37,0,173,0,116,0,230,0,210,0,12,0,8,0,24,0,162,0,137,0,112,0,148,0,0,0,72,0,5,0,237,0,245,0,68,0,55,0,115,0,0,0,95,0,226,0,99,0,0,0,191,0,226,0,78,0,0,0,155,0,171,0,251,0,85,0,156,0,143,0,55,0,145,0,0,0,28,0,168,0,163,0,148,0,41,0,51,0,13,0,35,0,99,0,242,0,37,0,113,0,116,0,0,0,0,0,105,0,203,0,245,0,13,0,222,0,196,0,9,0,107,0,208,0,168,0,141,0,254,0,188,0,0,0,185,0,80,0,45,0,126,0,232,0,239,0,182,0,0,0,0,0,0,0,139,0,248,0,0,0,255,0,44,0,0,0,97,0,255,0,190,0,169,0,0,0,154,0,254,0,118,0,0,0,92,0,230,0,41,0,33,0,59,0,76,0,0,0,89,0,213,0,95,0,249,0,221,0,14,0,0,0,98,0,0,0,22,0,229,0,162,0,0,0,228,0,136,0,49,0,22,0,5,0,28,0,35,0,73,0,0,0,67,0,133,0,251,0,183,0,0,0,0,0,239,0,174,0,0,0,159,0,205,0,117,0,98,0,0,0,227,0,255,0,73,0,0,0,23,0,99,0,51,0,240,0,3,0,87,0,245,0,50,0,165,0,184,0,0,0,186,0,0,0,62,0,37,0,208,0,0,0,162,0,131,0,85,0,35,0,80,0,0,0,0,0,179,0,133,0,0,0,241,0,92,0,0,0,113,0,60,0,243,0,45,0,0,0,186,0,167,0,206,0,53,0,0,0,0,0,131,0,167,0,0,0,121,0,0,0,227,0,0,0,30,0,0,0,0,0,196,0,159,0,0,0,15,0,75,0,12,0,127,0,70,0,0,0,0,0,197,0,10,0,244,0,227,0,192,0,10,0,255,0,101,0,127,0,56,0,233,0,247,0,158,0,56,0,165,0,0,0,51,0,253,0,200,0,133,0,0,0,0,0,38,0,192,0,0,0,224,0,17,0,190,0,0,0,150,0,71,0,243,0,0,0,248,0,0,0,204,0,0,0,28,0,0,0,161,0,63,0,229,0,235,0,162,0,27,0,147,0,0,0,43,0,235,0,224,0,177,0,80,0,0,0,143,0,151,0,251,0,28,0,157,0,184,0,142,0,98,0,158,0,14,0,38,0,19,0,0,0,0,0,0,0,155,0,0,0,2,0,28,0,64,0,38,0,0,0,108,0,104,0,0,0,42,0,158,0,229,0,105,0,0,0,67,0,0,0,67,0,145,0,126,0,47,0,0,0,53,0,0,0,0,0,0,0,0,0,117,0,0,0,112,0,169,0,0,0,252,0,28,0,45,0,76,0,102,0,0,0,166,0,214,0,127,0,167,0,212,0,0,0,178,0,133,0,144,0,200,0,45,0,15,0,37,0,0,0,57,0,0,0,54,0,148,0,230,0,87,0,200,0,0,0,0,0,27,0,0,0,76,0,237,0,116,0,0,0,0,0,0,0,209,0,122,0,28,0,32,0,15,0,206,0,217,0,73,0,198,0,121,0,0,0,186,0,130,0,0,0,6,0,86,0,225,0,1,0,106,0,211,0,130,0,56,0,0,0,205,0,247,0,92,0,103,0,202,0,204,0,237,0,108,0,167,0,13,0,51,0,79,0,26,0,222,0,55,0,213,0,0,0,145,0,159,0,212,0,118,0,0,0,42,0,189,0,0,0,192,0,122,0,183,0,250,0,50,0,140,0,0,0,28,0,64,0,142,0,110,0,137,0,124,0,0,0,66,0,216,0,83,0,250,0,0,0,0,0,251,0,0,0,63,0,133,0,79,0,49,0,100,0,0,0,0,0,34,0,148,0,247,0,235,0,107,0,29,0,80,0,0,0,230,0,62,0,209,0,26,0,123,0,93,0,127,0,246,0,69,0,138,0,135,0,70,0,138,0,0,0,218,0,0,0,110,0,140,0,0,0,234,0,141,0,208,0,97,0,163,0,118,0,67,0,69,0,0,0,122,0,172,0,142,0,114,0,85,0,0,0,207,0,174,0);
signal scenario_full  : scenario_type := (2,31,117,31,230,31,215,31,112,31,17,31,122,31,122,30,104,31,239,31,46,31,12,31,74,31,22,31,156,31,52,31,52,30,67,31,246,31,45,31,6,31,66,31,66,30,62,31,62,30,51,31,144,31,144,30,105,31,105,30,105,29,231,31,67,31,57,31,247,31,242,31,242,30,29,31,232,31,140,31,140,30,140,29,60,31,68,31,223,31,162,31,162,30,244,31,244,30,108,31,108,30,233,31,231,31,3,31,179,31,139,31,64,31,64,30,233,31,96,31,68,31,190,31,190,30,132,31,59,31,47,31,236,31,242,31,162,31,162,30,182,31,57,31,179,31,179,30,179,29,224,31,224,30,171,31,171,30,9,31,237,31,237,30,237,29,129,31,129,30,4,31,163,31,183,31,182,31,182,30,215,31,34,31,215,31,215,30,18,31,133,31,133,30,134,31,103,31,240,31,220,31,223,31,225,31,210,31,207,31,70,31,70,30,70,29,130,31,147,31,147,30,154,31,137,31,13,31,176,31,121,31,221,31,170,31,145,31,237,31,212,31,212,30,97,31,239,31,229,31,198,31,239,31,239,30,101,31,107,31,236,31,44,31,123,31,110,31,110,30,110,29,254,31,202,31,104,31,156,31,156,30,156,29,25,31,52,31,52,30,31,31,227,31,90,31,93,31,9,31,190,31,84,31,254,31,254,30,225,31,157,31,58,31,58,30,228,31,137,31,26,31,26,30,31,31,31,30,31,29,190,31,250,31,96,31,26,31,45,31,62,31,171,31,76,31,65,31,65,30,65,29,245,31,100,31,19,31,80,31,190,31,14,31,148,31,228,31,19,31,85,31,208,31,208,30,211,31,241,31,241,30,111,31,150,31,65,31,97,31,118,31,135,31,241,31,123,31,217,31,229,31,145,31,162,31,247,31,51,31,51,30,51,29,51,28,114,31,147,31,213,31,178,31,218,31,17,31,66,31,80,31,211,31,252,31,107,31,232,31,58,31,254,31,108,31,133,31,79,31,211,31,80,31,80,30,197,31,39,31,167,31,53,31,125,31,28,31,41,31,96,31,130,31,246,31,83,31,93,31,150,31,134,31,26,31,33,31,95,31,90,31,39,31,221,31,159,31,103,31,42,31,212,31,207,31,207,30,207,29,207,28,207,27,226,31,6,31,246,31,110,31,240,31,240,30,240,29,84,31,129,31,102,31,36,31,36,30,24,31,38,31,101,31,101,30,101,29,187,31,30,31,207,31,102,31,172,31,101,31,120,31,104,31,104,30,212,31,31,31,31,30,177,31,237,31,208,31,208,30,111,31,174,31,51,31,51,30,49,31,69,31,69,30,224,31,213,31,99,31,199,31,239,31,242,31,54,31,54,30,191,31,191,30,145,31,220,31,186,31,68,31,40,31,163,31,163,30,213,31,118,31,93,31,93,30,232,31,185,31,167,31,46,31,183,31,160,31,61,31,159,31,252,31,139,31,245,31,176,31,176,30,167,31,167,30,97,31,97,30,97,29,166,31,166,30,100,31,241,31,241,30,170,31,149,31,162,31,195,31,101,31,222,31,121,31,171,31,239,31,215,31,88,31,191,31,48,31,98,31,177,31,177,30,47,31,174,31,95,31,164,31,144,31,164,31,140,31,29,31,29,30,225,31,109,31,210,31,19,31,184,31,112,31,218,31,66,31,247,31,237,31,243,31,158,31,171,31,4,31,40,31,79,31,79,30,177,31,123,31,123,30,194,31,245,31,6,31,6,30,140,31,140,30,127,31,36,31,2,31,182,31,196,31,196,30,25,31,25,30,25,29,138,31,9,31,116,31,123,31,37,31,85,31,194,31,194,30,194,29,50,31,19,31,19,30,180,31,180,30,158,31,5,31,113,31,130,31,3,31,40,31,130,31,41,31,3,31,3,30,134,31,220,31,220,30,232,31,57,31,57,30,57,29,74,31,200,31,168,31,168,30,175,31,63,31,63,30,91,31,91,30,165,31,255,31,69,31,240,31,223,31,69,31,96,31,96,30,96,29,96,28,136,31,128,31,23,31,11,31,240,31,88,31,156,31,144,31,53,31,52,31,152,31,110,31,184,31,168,31,186,31,76,31,218,31,62,31,148,31,126,31,206,31,177,31,117,31,157,31,254,31,152,31,241,31,58,31,58,30,66,31,36,31,140,31,66,31,146,31,245,31,170,31,170,30,170,29,170,28,9,31,102,31,76,31,67,31,67,30,65,31,187,31,187,30,64,31,57,31,183,31,87,31,12,31,245,31,228,31,34,31,67,31,67,30,67,29,59,31,59,30,59,29,59,28,57,31,125,31,125,30,37,31,173,31,116,31,230,31,210,31,12,31,8,31,24,31,162,31,137,31,112,31,148,31,148,30,72,31,5,31,237,31,245,31,68,31,55,31,115,31,115,30,95,31,226,31,99,31,99,30,191,31,226,31,78,31,78,30,155,31,171,31,251,31,85,31,156,31,143,31,55,31,145,31,145,30,28,31,168,31,163,31,148,31,41,31,51,31,13,31,35,31,99,31,242,31,37,31,113,31,116,31,116,30,116,29,105,31,203,31,245,31,13,31,222,31,196,31,9,31,107,31,208,31,168,31,141,31,254,31,188,31,188,30,185,31,80,31,45,31,126,31,232,31,239,31,182,31,182,30,182,29,182,28,139,31,248,31,248,30,255,31,44,31,44,30,97,31,255,31,190,31,169,31,169,30,154,31,254,31,118,31,118,30,92,31,230,31,41,31,33,31,59,31,76,31,76,30,89,31,213,31,95,31,249,31,221,31,14,31,14,30,98,31,98,30,22,31,229,31,162,31,162,30,228,31,136,31,49,31,22,31,5,31,28,31,35,31,73,31,73,30,67,31,133,31,251,31,183,31,183,30,183,29,239,31,174,31,174,30,159,31,205,31,117,31,98,31,98,30,227,31,255,31,73,31,73,30,23,31,99,31,51,31,240,31,3,31,87,31,245,31,50,31,165,31,184,31,184,30,186,31,186,30,62,31,37,31,208,31,208,30,162,31,131,31,85,31,35,31,80,31,80,30,80,29,179,31,133,31,133,30,241,31,92,31,92,30,113,31,60,31,243,31,45,31,45,30,186,31,167,31,206,31,53,31,53,30,53,29,131,31,167,31,167,30,121,31,121,30,227,31,227,30,30,31,30,30,30,29,196,31,159,31,159,30,15,31,75,31,12,31,127,31,70,31,70,30,70,29,197,31,10,31,244,31,227,31,192,31,10,31,255,31,101,31,127,31,56,31,233,31,247,31,158,31,56,31,165,31,165,30,51,31,253,31,200,31,133,31,133,30,133,29,38,31,192,31,192,30,224,31,17,31,190,31,190,30,150,31,71,31,243,31,243,30,248,31,248,30,204,31,204,30,28,31,28,30,161,31,63,31,229,31,235,31,162,31,27,31,147,31,147,30,43,31,235,31,224,31,177,31,80,31,80,30,143,31,151,31,251,31,28,31,157,31,184,31,142,31,98,31,158,31,14,31,38,31,19,31,19,30,19,29,19,28,155,31,155,30,2,31,28,31,64,31,38,31,38,30,108,31,104,31,104,30,42,31,158,31,229,31,105,31,105,30,67,31,67,30,67,31,145,31,126,31,47,31,47,30,53,31,53,30,53,29,53,28,53,27,117,31,117,30,112,31,169,31,169,30,252,31,28,31,45,31,76,31,102,31,102,30,166,31,214,31,127,31,167,31,212,31,212,30,178,31,133,31,144,31,200,31,45,31,15,31,37,31,37,30,57,31,57,30,54,31,148,31,230,31,87,31,200,31,200,30,200,29,27,31,27,30,76,31,237,31,116,31,116,30,116,29,116,28,209,31,122,31,28,31,32,31,15,31,206,31,217,31,73,31,198,31,121,31,121,30,186,31,130,31,130,30,6,31,86,31,225,31,1,31,106,31,211,31,130,31,56,31,56,30,205,31,247,31,92,31,103,31,202,31,204,31,237,31,108,31,167,31,13,31,51,31,79,31,26,31,222,31,55,31,213,31,213,30,145,31,159,31,212,31,118,31,118,30,42,31,189,31,189,30,192,31,122,31,183,31,250,31,50,31,140,31,140,30,28,31,64,31,142,31,110,31,137,31,124,31,124,30,66,31,216,31,83,31,250,31,250,30,250,29,251,31,251,30,63,31,133,31,79,31,49,31,100,31,100,30,100,29,34,31,148,31,247,31,235,31,107,31,29,31,80,31,80,30,230,31,62,31,209,31,26,31,123,31,93,31,127,31,246,31,69,31,138,31,135,31,70,31,138,31,138,30,218,31,218,30,110,31,140,31,140,30,234,31,141,31,208,31,97,31,163,31,118,31,67,31,69,31,69,30,122,31,172,31,142,31,114,31,85,31,85,30,207,31,174,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
