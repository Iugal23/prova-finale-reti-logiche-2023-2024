-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_530 is
end project_tb_530;

architecture project_tb_arch_530 of project_tb_530 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 696;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (111,0,73,0,235,0,36,0,69,0,251,0,160,0,170,0,23,0,82,0,152,0,0,0,97,0,60,0,98,0,0,0,97,0,0,0,0,0,51,0,192,0,0,0,154,0,196,0,0,0,151,0,37,0,147,0,0,0,148,0,101,0,0,0,0,0,163,0,117,0,41,0,234,0,0,0,0,0,0,0,238,0,11,0,0,0,51,0,0,0,183,0,67,0,86,0,0,0,104,0,0,0,178,0,187,0,86,0,217,0,23,0,197,0,217,0,0,0,12,0,134,0,178,0,0,0,0,0,15,0,131,0,69,0,97,0,173,0,201,0,92,0,35,0,80,0,27,0,198,0,76,0,146,0,0,0,60,0,0,0,79,0,57,0,147,0,196,0,48,0,179,0,255,0,178,0,216,0,123,0,254,0,16,0,26,0,178,0,148,0,3,0,245,0,0,0,0,0,68,0,247,0,22,0,14,0,60,0,250,0,135,0,0,0,230,0,41,0,22,0,199,0,0,0,42,0,169,0,92,0,93,0,131,0,0,0,2,0,140,0,114,0,5,0,89,0,160,0,120,0,19,0,84,0,234,0,161,0,180,0,239,0,0,0,0,0,77,0,0,0,26,0,207,0,53,0,248,0,26,0,129,0,49,0,153,0,0,0,195,0,72,0,109,0,204,0,138,0,138,0,125,0,134,0,50,0,244,0,175,0,145,0,83,0,73,0,42,0,0,0,27,0,105,0,0,0,39,0,235,0,243,0,203,0,251,0,130,0,243,0,23,0,14,0,129,0,72,0,0,0,94,0,21,0,81,0,53,0,75,0,0,0,0,0,202,0,45,0,39,0,0,0,0,0,148,0,248,0,90,0,136,0,122,0,234,0,203,0,42,0,188,0,219,0,184,0,0,0,251,0,121,0,23,0,244,0,164,0,185,0,0,0,0,0,248,0,0,0,237,0,253,0,227,0,0,0,9,0,0,0,0,0,20,0,65,0,255,0,221,0,86,0,0,0,0,0,122,0,167,0,76,0,83,0,64,0,67,0,0,0,215,0,107,0,81,0,10,0,155,0,85,0,137,0,26,0,0,0,214,0,0,0,1,0,0,0,0,0,70,0,0,0,8,0,5,0,77,0,89,0,230,0,0,0,208,0,4,0,124,0,0,0,78,0,121,0,246,0,0,0,62,0,228,0,155,0,103,0,255,0,223,0,165,0,93,0,125,0,138,0,66,0,3,0,0,0,115,0,221,0,36,0,113,0,211,0,4,0,33,0,242,0,33,0,0,0,0,0,0,0,13,0,135,0,0,0,92,0,221,0,172,0,238,0,245,0,100,0,200,0,96,0,53,0,0,0,80,0,191,0,135,0,131,0,203,0,82,0,0,0,136,0,13,0,220,0,53,0,129,0,240,0,0,0,218,0,166,0,47,0,124,0,22,0,203,0,24,0,243,0,0,0,70,0,12,0,78,0,9,0,214,0,159,0,71,0,11,0,0,0,0,0,97,0,238,0,0,0,229,0,0,0,0,0,0,0,0,0,126,0,121,0,65,0,58,0,0,0,50,0,0,0,150,0,8,0,0,0,40,0,86,0,0,0,37,0,216,0,73,0,133,0,68,0,0,0,79,0,247,0,223,0,169,0,1,0,0,0,94,0,0,0,80,0,0,0,243,0,215,0,206,0,247,0,70,0,42,0,0,0,72,0,0,0,191,0,0,0,0,0,217,0,1,0,70,0,130,0,65,0,45,0,0,0,5,0,107,0,161,0,0,0,34,0,104,0,125,0,56,0,0,0,127,0,0,0,0,0,126,0,200,0,236,0,162,0,213,0,245,0,122,0,221,0,169,0,145,0,22,0,0,0,201,0,166,0,36,0,158,0,143,0,97,0,234,0,0,0,133,0,179,0,220,0,107,0,3,0,0,0,32,0,203,0,116,0,0,0,55,0,37,0,0,0,179,0,247,0,1,0,52,0,71,0,0,0,29,0,31,0,245,0,148,0,222,0,154,0,155,0,41,0,119,0,11,0,184,0,12,0,0,0,0,0,254,0,96,0,180,0,0,0,0,0,218,0,63,0,210,0,104,0,5,0,248,0,163,0,149,0,0,0,0,0,168,0,173,0,0,0,91,0,0,0,162,0,177,0,176,0,199,0,137,0,11,0,4,0,9,0,105,0,107,0,184,0,11,0,92,0,73,0,50,0,219,0,245,0,255,0,37,0,202,0,123,0,8,0,46,0,0,0,20,0,0,0,204,0,176,0,33,0,232,0,67,0,4,0,43,0,74,0,170,0,43,0,33,0,118,0,0,0,139,0,241,0,82,0,142,0,0,0,46,0,145,0,134,0,147,0,184,0,27,0,134,0,199,0,120,0,0,0,196,0,63,0,182,0,61,0,0,0,247,0,94,0,0,0,0,0,71,0,196,0,98,0,130,0,119,0,189,0,14,0,110,0,81,0,34,0,38,0,0,0,105,0,241,0,64,0,209,0,103,0,20,0,0,0,92,0,0,0,118,0,155,0,0,0,200,0,55,0,0,0,112,0,146,0,154,0,0,0,104,0,50,0,67,0,0,0,181,0,123,0,81,0,154,0,60,0,171,0,160,0,116,0,212,0,0,0,221,0,184,0,93,0,0,0,68,0,0,0,108,0,254,0,187,0,218,0,134,0,0,0,152,0,105,0,170,0,0,0,0,0,108,0,215,0,18,0,199,0,236,0,153,0,33,0,52,0,58,0,39,0,37,0,135,0,33,0,0,0,133,0,173,0,92,0,0,0,0,0,138,0,123,0,3,0,150,0,171,0,88,0,0,0,31,0,49,0,160,0,253,0,81,0,16,0,181,0,247,0,194,0,202,0,198,0,0,0,118,0,244,0,193,0,146,0,245,0,138,0,6,0,201,0,0,0,232,0,0,0,13,0,236,0,9,0,201,0,128,0,186,0,84,0,108,0,227,0,70,0,0,0,78,0,0,0,0,0,203,0,29,0,98,0,146,0,106,0,133,0,221,0,255,0,238,0,102,0,74,0,216,0,252,0,104,0,153,0,60,0,209,0,234,0,0,0,0,0,0,0,106,0,164,0,239,0,138,0,96,0,226,0,243,0,0,0,75,0,0,0,52,0,53,0,66,0,207,0,154,0);
signal scenario_full  : scenario_type := (111,31,73,31,235,31,36,31,69,31,251,31,160,31,170,31,23,31,82,31,152,31,152,30,97,31,60,31,98,31,98,30,97,31,97,30,97,29,51,31,192,31,192,30,154,31,196,31,196,30,151,31,37,31,147,31,147,30,148,31,101,31,101,30,101,29,163,31,117,31,41,31,234,31,234,30,234,29,234,28,238,31,11,31,11,30,51,31,51,30,183,31,67,31,86,31,86,30,104,31,104,30,178,31,187,31,86,31,217,31,23,31,197,31,217,31,217,30,12,31,134,31,178,31,178,30,178,29,15,31,131,31,69,31,97,31,173,31,201,31,92,31,35,31,80,31,27,31,198,31,76,31,146,31,146,30,60,31,60,30,79,31,57,31,147,31,196,31,48,31,179,31,255,31,178,31,216,31,123,31,254,31,16,31,26,31,178,31,148,31,3,31,245,31,245,30,245,29,68,31,247,31,22,31,14,31,60,31,250,31,135,31,135,30,230,31,41,31,22,31,199,31,199,30,42,31,169,31,92,31,93,31,131,31,131,30,2,31,140,31,114,31,5,31,89,31,160,31,120,31,19,31,84,31,234,31,161,31,180,31,239,31,239,30,239,29,77,31,77,30,26,31,207,31,53,31,248,31,26,31,129,31,49,31,153,31,153,30,195,31,72,31,109,31,204,31,138,31,138,31,125,31,134,31,50,31,244,31,175,31,145,31,83,31,73,31,42,31,42,30,27,31,105,31,105,30,39,31,235,31,243,31,203,31,251,31,130,31,243,31,23,31,14,31,129,31,72,31,72,30,94,31,21,31,81,31,53,31,75,31,75,30,75,29,202,31,45,31,39,31,39,30,39,29,148,31,248,31,90,31,136,31,122,31,234,31,203,31,42,31,188,31,219,31,184,31,184,30,251,31,121,31,23,31,244,31,164,31,185,31,185,30,185,29,248,31,248,30,237,31,253,31,227,31,227,30,9,31,9,30,9,29,20,31,65,31,255,31,221,31,86,31,86,30,86,29,122,31,167,31,76,31,83,31,64,31,67,31,67,30,215,31,107,31,81,31,10,31,155,31,85,31,137,31,26,31,26,30,214,31,214,30,1,31,1,30,1,29,70,31,70,30,8,31,5,31,77,31,89,31,230,31,230,30,208,31,4,31,124,31,124,30,78,31,121,31,246,31,246,30,62,31,228,31,155,31,103,31,255,31,223,31,165,31,93,31,125,31,138,31,66,31,3,31,3,30,115,31,221,31,36,31,113,31,211,31,4,31,33,31,242,31,33,31,33,30,33,29,33,28,13,31,135,31,135,30,92,31,221,31,172,31,238,31,245,31,100,31,200,31,96,31,53,31,53,30,80,31,191,31,135,31,131,31,203,31,82,31,82,30,136,31,13,31,220,31,53,31,129,31,240,31,240,30,218,31,166,31,47,31,124,31,22,31,203,31,24,31,243,31,243,30,70,31,12,31,78,31,9,31,214,31,159,31,71,31,11,31,11,30,11,29,97,31,238,31,238,30,229,31,229,30,229,29,229,28,229,27,126,31,121,31,65,31,58,31,58,30,50,31,50,30,150,31,8,31,8,30,40,31,86,31,86,30,37,31,216,31,73,31,133,31,68,31,68,30,79,31,247,31,223,31,169,31,1,31,1,30,94,31,94,30,80,31,80,30,243,31,215,31,206,31,247,31,70,31,42,31,42,30,72,31,72,30,191,31,191,30,191,29,217,31,1,31,70,31,130,31,65,31,45,31,45,30,5,31,107,31,161,31,161,30,34,31,104,31,125,31,56,31,56,30,127,31,127,30,127,29,126,31,200,31,236,31,162,31,213,31,245,31,122,31,221,31,169,31,145,31,22,31,22,30,201,31,166,31,36,31,158,31,143,31,97,31,234,31,234,30,133,31,179,31,220,31,107,31,3,31,3,30,32,31,203,31,116,31,116,30,55,31,37,31,37,30,179,31,247,31,1,31,52,31,71,31,71,30,29,31,31,31,245,31,148,31,222,31,154,31,155,31,41,31,119,31,11,31,184,31,12,31,12,30,12,29,254,31,96,31,180,31,180,30,180,29,218,31,63,31,210,31,104,31,5,31,248,31,163,31,149,31,149,30,149,29,168,31,173,31,173,30,91,31,91,30,162,31,177,31,176,31,199,31,137,31,11,31,4,31,9,31,105,31,107,31,184,31,11,31,92,31,73,31,50,31,219,31,245,31,255,31,37,31,202,31,123,31,8,31,46,31,46,30,20,31,20,30,204,31,176,31,33,31,232,31,67,31,4,31,43,31,74,31,170,31,43,31,33,31,118,31,118,30,139,31,241,31,82,31,142,31,142,30,46,31,145,31,134,31,147,31,184,31,27,31,134,31,199,31,120,31,120,30,196,31,63,31,182,31,61,31,61,30,247,31,94,31,94,30,94,29,71,31,196,31,98,31,130,31,119,31,189,31,14,31,110,31,81,31,34,31,38,31,38,30,105,31,241,31,64,31,209,31,103,31,20,31,20,30,92,31,92,30,118,31,155,31,155,30,200,31,55,31,55,30,112,31,146,31,154,31,154,30,104,31,50,31,67,31,67,30,181,31,123,31,81,31,154,31,60,31,171,31,160,31,116,31,212,31,212,30,221,31,184,31,93,31,93,30,68,31,68,30,108,31,254,31,187,31,218,31,134,31,134,30,152,31,105,31,170,31,170,30,170,29,108,31,215,31,18,31,199,31,236,31,153,31,33,31,52,31,58,31,39,31,37,31,135,31,33,31,33,30,133,31,173,31,92,31,92,30,92,29,138,31,123,31,3,31,150,31,171,31,88,31,88,30,31,31,49,31,160,31,253,31,81,31,16,31,181,31,247,31,194,31,202,31,198,31,198,30,118,31,244,31,193,31,146,31,245,31,138,31,6,31,201,31,201,30,232,31,232,30,13,31,236,31,9,31,201,31,128,31,186,31,84,31,108,31,227,31,70,31,70,30,78,31,78,30,78,29,203,31,29,31,98,31,146,31,106,31,133,31,221,31,255,31,238,31,102,31,74,31,216,31,252,31,104,31,153,31,60,31,209,31,234,31,234,30,234,29,234,28,106,31,164,31,239,31,138,31,96,31,226,31,243,31,243,30,75,31,75,30,52,31,53,31,66,31,207,31,154,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
