-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 695;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (71,0,30,0,113,0,151,0,117,0,228,0,0,0,49,0,172,0,141,0,121,0,198,0,122,0,240,0,179,0,240,0,25,0,46,0,0,0,239,0,97,0,222,0,230,0,247,0,0,0,240,0,64,0,0,0,0,0,147,0,124,0,172,0,139,0,176,0,216,0,200,0,174,0,183,0,12,0,30,0,0,0,5,0,87,0,222,0,0,0,192,0,117,0,217,0,69,0,154,0,0,0,125,0,86,0,137,0,29,0,67,0,252,0,56,0,2,0,244,0,23,0,66,0,0,0,240,0,28,0,116,0,251,0,0,0,62,0,93,0,118,0,0,0,178,0,72,0,0,0,34,0,87,0,200,0,66,0,212,0,60,0,205,0,129,0,39,0,91,0,174,0,222,0,16,0,71,0,21,0,92,0,216,0,240,0,0,0,217,0,151,0,0,0,0,0,62,0,246,0,213,0,100,0,122,0,55,0,122,0,84,0,117,0,179,0,125,0,0,0,131,0,99,0,255,0,136,0,113,0,149,0,36,0,230,0,0,0,226,0,87,0,161,0,0,0,54,0,111,0,40,0,0,0,24,0,0,0,0,0,0,0,154,0,0,0,197,0,0,0,161,0,230,0,0,0,31,0,192,0,0,0,169,0,3,0,199,0,0,0,162,0,218,0,0,0,154,0,40,0,205,0,203,0,212,0,0,0,5,0,6,0,134,0,51,0,116,0,24,0,111,0,178,0,221,0,93,0,0,0,112,0,73,0,0,0,232,0,86,0,0,0,135,0,95,0,0,0,187,0,0,0,162,0,114,0,224,0,117,0,163,0,0,0,99,0,254,0,0,0,0,0,249,0,202,0,133,0,0,0,70,0,0,0,0,0,233,0,0,0,0,0,175,0,0,0,52,0,137,0,238,0,8,0,207,0,107,0,17,0,35,0,209,0,106,0,208,0,130,0,0,0,28,0,0,0,112,0,115,0,173,0,0,0,240,0,0,0,9,0,0,0,124,0,0,0,216,0,0,0,70,0,159,0,120,0,59,0,48,0,14,0,165,0,0,0,180,0,139,0,92,0,236,0,147,0,0,0,200,0,225,0,0,0,20,0,0,0,131,0,9,0,0,0,143,0,40,0,83,0,180,0,81,0,14,0,140,0,250,0,108,0,143,0,154,0,0,0,82,0,224,0,40,0,224,0,228,0,169,0,44,0,0,0,155,0,79,0,183,0,105,0,0,0,192,0,238,0,84,0,220,0,67,0,209,0,0,0,132,0,135,0,0,0,234,0,133,0,128,0,0,0,239,0,0,0,9,0,93,0,95,0,81,0,40,0,114,0,173,0,45,0,0,0,31,0,67,0,8,0,0,0,126,0,133,0,169,0,220,0,134,0,17,0,51,0,197,0,87,0,155,0,186,0,0,0,147,0,2,0,0,0,138,0,168,0,0,0,239,0,139,0,8,0,80,0,149,0,93,0,40,0,224,0,198,0,140,0,223,0,91,0,156,0,0,0,0,0,255,0,63,0,250,0,186,0,58,0,114,0,252,0,0,0,5,0,183,0,0,0,0,0,12,0,0,0,0,0,231,0,67,0,55,0,231,0,0,0,49,0,181,0,0,0,68,0,211,0,122,0,153,0,78,0,42,0,0,0,111,0,11,0,54,0,0,0,125,0,171,0,83,0,213,0,136,0,184,0,109,0,29,0,19,0,84,0,196,0,85,0,234,0,249,0,98,0,206,0,230,0,127,0,44,0,0,0,67,0,180,0,253,0,225,0,0,0,209,0,15,0,3,0,139,0,24,0,0,0,64,0,0,0,162,0,0,0,150,0,0,0,5,0,39,0,32,0,57,0,127,0,173,0,14,0,101,0,132,0,98,0,0,0,249,0,198,0,10,0,146,0,27,0,0,0,0,0,105,0,210,0,110,0,132,0,36,0,78,0,181,0,0,0,250,0,0,0,186,0,176,0,0,0,96,0,114,0,177,0,77,0,5,0,119,0,48,0,173,0,0,0,0,0,200,0,186,0,165,0,197,0,165,0,0,0,100,0,37,0,4,0,219,0,0,0,134,0,125,0,169,0,217,0,103,0,246,0,103,0,28,0,108,0,108,0,0,0,0,0,191,0,104,0,23,0,0,0,239,0,213,0,105,0,4,0,176,0,112,0,103,0,0,0,255,0,211,0,44,0,89,0,105,0,211,0,30,0,158,0,232,0,27,0,60,0,0,0,46,0,106,0,0,0,173,0,58,0,187,0,107,0,0,0,0,0,0,0,91,0,25,0,204,0,0,0,2,0,88,0,46,0,230,0,194,0,17,0,206,0,25,0,114,0,145,0,55,0,0,0,0,0,50,0,80,0,159,0,227,0,95,0,0,0,0,0,75,0,187,0,0,0,19,0,185,0,0,0,121,0,229,0,0,0,118,0,55,0,77,0,78,0,1,0,135,0,106,0,187,0,114,0,0,0,201,0,44,0,0,0,34,0,168,0,132,0,32,0,88,0,246,0,23,0,36,0,97,0,0,0,0,0,109,0,0,0,0,0,175,0,145,0,242,0,88,0,0,0,20,0,220,0,147,0,80,0,84,0,0,0,54,0,207,0,18,0,159,0,0,0,0,0,0,0,0,0,169,0,0,0,38,0,67,0,173,0,0,0,74,0,190,0,12,0,31,0,0,0,191,0,0,0,40,0,27,0,107,0,210,0,158,0,0,0,151,0,233,0,69,0,71,0,239,0,40,0,177,0,42,0,177,0,0,0,134,0,160,0,146,0,17,0,130,0,0,0,166,0,217,0,0,0,0,0,50,0,0,0,102,0,162,0,0,0,0,0,217,0,84,0,28,0,111,0,1,0,188,0,181,0,135,0,91,0,8,0,0,0,128,0,130,0,137,0,0,0,197,0,46,0,0,0,193,0,0,0,64,0,9,0,212,0,0,0,0,0,213,0,0,0,188,0,29,0,232,0,128,0,0,0,98,0,171,0,229,0,0,0,235,0,169,0,222,0,66,0,85,0,0,0,0,0,240,0,5,0,128,0,77,0,101,0,0,0,32,0,28,0,43,0,200,0,156,0,0,0,229,0,43,0,0,0,127,0,52,0,11,0,0,0,183,0,48,0,0,0,47,0,0,0,43,0);
signal scenario_full  : scenario_type := (71,31,30,31,113,31,151,31,117,31,228,31,228,30,49,31,172,31,141,31,121,31,198,31,122,31,240,31,179,31,240,31,25,31,46,31,46,30,239,31,97,31,222,31,230,31,247,31,247,30,240,31,64,31,64,30,64,29,147,31,124,31,172,31,139,31,176,31,216,31,200,31,174,31,183,31,12,31,30,31,30,30,5,31,87,31,222,31,222,30,192,31,117,31,217,31,69,31,154,31,154,30,125,31,86,31,137,31,29,31,67,31,252,31,56,31,2,31,244,31,23,31,66,31,66,30,240,31,28,31,116,31,251,31,251,30,62,31,93,31,118,31,118,30,178,31,72,31,72,30,34,31,87,31,200,31,66,31,212,31,60,31,205,31,129,31,39,31,91,31,174,31,222,31,16,31,71,31,21,31,92,31,216,31,240,31,240,30,217,31,151,31,151,30,151,29,62,31,246,31,213,31,100,31,122,31,55,31,122,31,84,31,117,31,179,31,125,31,125,30,131,31,99,31,255,31,136,31,113,31,149,31,36,31,230,31,230,30,226,31,87,31,161,31,161,30,54,31,111,31,40,31,40,30,24,31,24,30,24,29,24,28,154,31,154,30,197,31,197,30,161,31,230,31,230,30,31,31,192,31,192,30,169,31,3,31,199,31,199,30,162,31,218,31,218,30,154,31,40,31,205,31,203,31,212,31,212,30,5,31,6,31,134,31,51,31,116,31,24,31,111,31,178,31,221,31,93,31,93,30,112,31,73,31,73,30,232,31,86,31,86,30,135,31,95,31,95,30,187,31,187,30,162,31,114,31,224,31,117,31,163,31,163,30,99,31,254,31,254,30,254,29,249,31,202,31,133,31,133,30,70,31,70,30,70,29,233,31,233,30,233,29,175,31,175,30,52,31,137,31,238,31,8,31,207,31,107,31,17,31,35,31,209,31,106,31,208,31,130,31,130,30,28,31,28,30,112,31,115,31,173,31,173,30,240,31,240,30,9,31,9,30,124,31,124,30,216,31,216,30,70,31,159,31,120,31,59,31,48,31,14,31,165,31,165,30,180,31,139,31,92,31,236,31,147,31,147,30,200,31,225,31,225,30,20,31,20,30,131,31,9,31,9,30,143,31,40,31,83,31,180,31,81,31,14,31,140,31,250,31,108,31,143,31,154,31,154,30,82,31,224,31,40,31,224,31,228,31,169,31,44,31,44,30,155,31,79,31,183,31,105,31,105,30,192,31,238,31,84,31,220,31,67,31,209,31,209,30,132,31,135,31,135,30,234,31,133,31,128,31,128,30,239,31,239,30,9,31,93,31,95,31,81,31,40,31,114,31,173,31,45,31,45,30,31,31,67,31,8,31,8,30,126,31,133,31,169,31,220,31,134,31,17,31,51,31,197,31,87,31,155,31,186,31,186,30,147,31,2,31,2,30,138,31,168,31,168,30,239,31,139,31,8,31,80,31,149,31,93,31,40,31,224,31,198,31,140,31,223,31,91,31,156,31,156,30,156,29,255,31,63,31,250,31,186,31,58,31,114,31,252,31,252,30,5,31,183,31,183,30,183,29,12,31,12,30,12,29,231,31,67,31,55,31,231,31,231,30,49,31,181,31,181,30,68,31,211,31,122,31,153,31,78,31,42,31,42,30,111,31,11,31,54,31,54,30,125,31,171,31,83,31,213,31,136,31,184,31,109,31,29,31,19,31,84,31,196,31,85,31,234,31,249,31,98,31,206,31,230,31,127,31,44,31,44,30,67,31,180,31,253,31,225,31,225,30,209,31,15,31,3,31,139,31,24,31,24,30,64,31,64,30,162,31,162,30,150,31,150,30,5,31,39,31,32,31,57,31,127,31,173,31,14,31,101,31,132,31,98,31,98,30,249,31,198,31,10,31,146,31,27,31,27,30,27,29,105,31,210,31,110,31,132,31,36,31,78,31,181,31,181,30,250,31,250,30,186,31,176,31,176,30,96,31,114,31,177,31,77,31,5,31,119,31,48,31,173,31,173,30,173,29,200,31,186,31,165,31,197,31,165,31,165,30,100,31,37,31,4,31,219,31,219,30,134,31,125,31,169,31,217,31,103,31,246,31,103,31,28,31,108,31,108,31,108,30,108,29,191,31,104,31,23,31,23,30,239,31,213,31,105,31,4,31,176,31,112,31,103,31,103,30,255,31,211,31,44,31,89,31,105,31,211,31,30,31,158,31,232,31,27,31,60,31,60,30,46,31,106,31,106,30,173,31,58,31,187,31,107,31,107,30,107,29,107,28,91,31,25,31,204,31,204,30,2,31,88,31,46,31,230,31,194,31,17,31,206,31,25,31,114,31,145,31,55,31,55,30,55,29,50,31,80,31,159,31,227,31,95,31,95,30,95,29,75,31,187,31,187,30,19,31,185,31,185,30,121,31,229,31,229,30,118,31,55,31,77,31,78,31,1,31,135,31,106,31,187,31,114,31,114,30,201,31,44,31,44,30,34,31,168,31,132,31,32,31,88,31,246,31,23,31,36,31,97,31,97,30,97,29,109,31,109,30,109,29,175,31,145,31,242,31,88,31,88,30,20,31,220,31,147,31,80,31,84,31,84,30,54,31,207,31,18,31,159,31,159,30,159,29,159,28,159,27,169,31,169,30,38,31,67,31,173,31,173,30,74,31,190,31,12,31,31,31,31,30,191,31,191,30,40,31,27,31,107,31,210,31,158,31,158,30,151,31,233,31,69,31,71,31,239,31,40,31,177,31,42,31,177,31,177,30,134,31,160,31,146,31,17,31,130,31,130,30,166,31,217,31,217,30,217,29,50,31,50,30,102,31,162,31,162,30,162,29,217,31,84,31,28,31,111,31,1,31,188,31,181,31,135,31,91,31,8,31,8,30,128,31,130,31,137,31,137,30,197,31,46,31,46,30,193,31,193,30,64,31,9,31,212,31,212,30,212,29,213,31,213,30,188,31,29,31,232,31,128,31,128,30,98,31,171,31,229,31,229,30,235,31,169,31,222,31,66,31,85,31,85,30,85,29,240,31,5,31,128,31,77,31,101,31,101,30,32,31,28,31,43,31,200,31,156,31,156,30,229,31,43,31,43,30,127,31,52,31,11,31,11,30,183,31,48,31,48,30,47,31,47,30,43,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
