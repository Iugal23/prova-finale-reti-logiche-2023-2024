-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_153 is
end project_tb_153;

architecture project_tb_arch_153 of project_tb_153 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 808;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (40,0,166,0,0,0,108,0,10,0,0,0,131,0,206,0,120,0,6,0,77,0,16,0,0,0,0,0,148,0,240,0,121,0,77,0,0,0,0,0,147,0,125,0,46,0,0,0,171,0,180,0,154,0,0,0,170,0,210,0,12,0,133,0,45,0,0,0,129,0,189,0,0,0,140,0,79,0,183,0,0,0,164,0,0,0,254,0,80,0,0,0,79,0,172,0,164,0,93,0,0,0,174,0,233,0,243,0,43,0,0,0,168,0,77,0,187,0,234,0,224,0,1,0,0,0,168,0,185,0,151,0,200,0,211,0,135,0,215,0,0,0,0,0,140,0,0,0,32,0,182,0,112,0,248,0,182,0,12,0,207,0,243,0,192,0,254,0,0,0,153,0,191,0,224,0,159,0,63,0,110,0,212,0,101,0,0,0,146,0,114,0,102,0,109,0,198,0,94,0,0,0,55,0,135,0,201,0,176,0,222,0,61,0,36,0,60,0,110,0,193,0,194,0,131,0,114,0,125,0,44,0,0,0,0,0,48,0,94,0,20,0,0,0,124,0,117,0,0,0,123,0,39,0,119,0,221,0,0,0,124,0,106,0,0,0,1,0,163,0,195,0,220,0,172,0,121,0,0,0,0,0,136,0,100,0,0,0,238,0,221,0,244,0,0,0,0,0,254,0,81,0,86,0,0,0,138,0,217,0,0,0,0,0,224,0,160,0,0,0,211,0,45,0,115,0,40,0,175,0,17,0,104,0,0,0,151,0,182,0,162,0,0,0,2,0,0,0,213,0,91,0,129,0,134,0,0,0,137,0,84,0,49,0,0,0,174,0,0,0,201,0,164,0,88,0,97,0,59,0,168,0,0,0,29,0,0,0,241,0,8,0,254,0,40,0,0,0,177,0,16,0,198,0,222,0,0,0,101,0,193,0,191,0,44,0,135,0,0,0,25,0,0,0,0,0,252,0,0,0,224,0,0,0,21,0,218,0,227,0,175,0,66,0,57,0,0,0,0,0,229,0,135,0,0,0,182,0,191,0,140,0,145,0,183,0,70,0,93,0,27,0,117,0,99,0,191,0,219,0,108,0,15,0,0,0,244,0,59,0,137,0,55,0,95,0,18,0,201,0,0,0,0,0,0,0,218,0,30,0,0,0,246,0,239,0,159,0,168,0,134,0,140,0,25,0,158,0,75,0,225,0,125,0,70,0,83,0,170,0,224,0,26,0,111,0,231,0,104,0,219,0,0,0,169,0,183,0,148,0,194,0,47,0,4,0,251,0,215,0,109,0,0,0,242,0,31,0,0,0,0,0,0,0,0,0,194,0,234,0,0,0,0,0,0,0,201,0,0,0,0,0,106,0,37,0,0,0,0,0,94,0,209,0,97,0,126,0,219,0,40,0,184,0,0,0,125,0,87,0,0,0,96,0,245,0,137,0,0,0,251,0,0,0,0,0,161,0,144,0,56,0,223,0,36,0,17,0,145,0,173,0,106,0,217,0,27,0,236,0,72,0,0,0,0,0,41,0,219,0,66,0,0,0,194,0,189,0,0,0,217,0,43,0,117,0,180,0,162,0,118,0,62,0,4,0,128,0,0,0,47,0,77,0,13,0,240,0,255,0,10,0,83,0,0,0,178,0,207,0,221,0,97,0,0,0,67,0,40,0,0,0,182,0,173,0,218,0,29,0,67,0,237,0,0,0,210,0,243,0,10,0,193,0,117,0,14,0,0,0,32,0,211,0,0,0,161,0,52,0,251,0,204,0,91,0,0,0,240,0,74,0,93,0,43,0,248,0,197,0,173,0,214,0,96,0,216,0,0,0,3,0,142,0,136,0,44,0,70,0,103,0,216,0,98,0,0,0,8,0,244,0,172,0,251,0,99,0,221,0,103,0,0,0,137,0,108,0,102,0,140,0,91,0,0,0,91,0,96,0,245,0,99,0,0,0,7,0,161,0,200,0,192,0,155,0,240,0,232,0,43,0,44,0,0,0,0,0,0,0,255,0,29,0,184,0,235,0,20,0,67,0,147,0,102,0,157,0,215,0,43,0,54,0,79,0,137,0,96,0,25,0,45,0,111,0,165,0,0,0,250,0,113,0,0,0,249,0,22,0,117,0,135,0,192,0,21,0,72,0,160,0,134,0,35,0,167,0,48,0,150,0,93,0,220,0,155,0,0,0,6,0,182,0,150,0,191,0,0,0,222,0,0,0,253,0,0,0,221,0,134,0,224,0,0,0,0,0,245,0,243,0,240,0,228,0,151,0,15,0,231,0,93,0,52,0,164,0,205,0,0,0,85,0,22,0,247,0,0,0,43,0,158,0,245,0,114,0,65,0,112,0,251,0,0,0,0,0,234,0,0,0,65,0,28,0,0,0,93,0,12,0,119,0,0,0,64,0,0,0,214,0,41,0,0,0,119,0,168,0,113,0,216,0,48,0,254,0,140,0,132,0,139,0,166,0,249,0,0,0,240,0,0,0,216,0,202,0,195,0,169,0,0,0,56,0,193,0,75,0,235,0,0,0,0,0,204,0,35,0,129,0,102,0,230,0,38,0,0,0,0,0,66,0,0,0,160,0,137,0,221,0,61,0,239,0,0,0,128,0,192,0,0,0,0,0,41,0,0,0,219,0,0,0,73,0,81,0,0,0,0,0,45,0,132,0,32,0,138,0,202,0,198,0,0,0,96,0,77,0,255,0,246,0,0,0,0,0,241,0,53,0,19,0,5,0,131,0,50,0,214,0,0,0,47,0,222,0,0,0,40,0,19,0,85,0,0,0,99,0,77,0,243,0,0,0,235,0,68,0,0,0,190,0,13,0,149,0,0,0,152,0,12,0,12,0,225,0,249,0,22,0,97,0,237,0,49,0,0,0,236,0,0,0,56,0,33,0,146,0,181,0,122,0,220,0,109,0,191,0,252,0,81,0,246,0,0,0,233,0,63,0,122,0,248,0,199,0,0,0,168,0,123,0,215,0,181,0,74,0,159,0,25,0,29,0,200,0,135,0,2,0,156,0,17,0,205,0,200,0,249,0,107,0,79,0,192,0,139,0,254,0,255,0,120,0,111,0,150,0,88,0,134,0,0,0,210,0,0,0,0,0,0,0,0,0,242,0,127,0,231,0,129,0,3,0,65,0,97,0,192,0,71,0,141,0,237,0,0,0,0,0,0,0,18,0,167,0,135,0,0,0,194,0,200,0,111,0,0,0,163,0,254,0,27,0,0,0,0,0,61,0,225,0,49,0,12,0,0,0,39,0,148,0,62,0,145,0,141,0,136,0,35,0,96,0,192,0,67,0,255,0,0,0,154,0,48,0,0,0,216,0,177,0,130,0,158,0,58,0,0,0,242,0,230,0,244,0,106,0,139,0,27,0,57,0,115,0,228,0,28,0,254,0,0,0,186,0,155,0,212,0,222,0,0,0,218,0,89,0,180,0,0,0,247,0,0,0,154,0,158,0,227,0,184,0,12,0,61,0,172,0,98,0,173,0,76,0,0,0,0,0,30,0,129,0,139,0,118,0,229,0,229,0,61,0,0,0,224,0,209,0,209,0,0,0,45,0,0,0,168,0,164,0,16,0,183,0,99,0,218,0,0,0,36,0,164,0,189,0,71,0,173,0,0,0);
signal scenario_full  : scenario_type := (40,31,166,31,166,30,108,31,10,31,10,30,131,31,206,31,120,31,6,31,77,31,16,31,16,30,16,29,148,31,240,31,121,31,77,31,77,30,77,29,147,31,125,31,46,31,46,30,171,31,180,31,154,31,154,30,170,31,210,31,12,31,133,31,45,31,45,30,129,31,189,31,189,30,140,31,79,31,183,31,183,30,164,31,164,30,254,31,80,31,80,30,79,31,172,31,164,31,93,31,93,30,174,31,233,31,243,31,43,31,43,30,168,31,77,31,187,31,234,31,224,31,1,31,1,30,168,31,185,31,151,31,200,31,211,31,135,31,215,31,215,30,215,29,140,31,140,30,32,31,182,31,112,31,248,31,182,31,12,31,207,31,243,31,192,31,254,31,254,30,153,31,191,31,224,31,159,31,63,31,110,31,212,31,101,31,101,30,146,31,114,31,102,31,109,31,198,31,94,31,94,30,55,31,135,31,201,31,176,31,222,31,61,31,36,31,60,31,110,31,193,31,194,31,131,31,114,31,125,31,44,31,44,30,44,29,48,31,94,31,20,31,20,30,124,31,117,31,117,30,123,31,39,31,119,31,221,31,221,30,124,31,106,31,106,30,1,31,163,31,195,31,220,31,172,31,121,31,121,30,121,29,136,31,100,31,100,30,238,31,221,31,244,31,244,30,244,29,254,31,81,31,86,31,86,30,138,31,217,31,217,30,217,29,224,31,160,31,160,30,211,31,45,31,115,31,40,31,175,31,17,31,104,31,104,30,151,31,182,31,162,31,162,30,2,31,2,30,213,31,91,31,129,31,134,31,134,30,137,31,84,31,49,31,49,30,174,31,174,30,201,31,164,31,88,31,97,31,59,31,168,31,168,30,29,31,29,30,241,31,8,31,254,31,40,31,40,30,177,31,16,31,198,31,222,31,222,30,101,31,193,31,191,31,44,31,135,31,135,30,25,31,25,30,25,29,252,31,252,30,224,31,224,30,21,31,218,31,227,31,175,31,66,31,57,31,57,30,57,29,229,31,135,31,135,30,182,31,191,31,140,31,145,31,183,31,70,31,93,31,27,31,117,31,99,31,191,31,219,31,108,31,15,31,15,30,244,31,59,31,137,31,55,31,95,31,18,31,201,31,201,30,201,29,201,28,218,31,30,31,30,30,246,31,239,31,159,31,168,31,134,31,140,31,25,31,158,31,75,31,225,31,125,31,70,31,83,31,170,31,224,31,26,31,111,31,231,31,104,31,219,31,219,30,169,31,183,31,148,31,194,31,47,31,4,31,251,31,215,31,109,31,109,30,242,31,31,31,31,30,31,29,31,28,31,27,194,31,234,31,234,30,234,29,234,28,201,31,201,30,201,29,106,31,37,31,37,30,37,29,94,31,209,31,97,31,126,31,219,31,40,31,184,31,184,30,125,31,87,31,87,30,96,31,245,31,137,31,137,30,251,31,251,30,251,29,161,31,144,31,56,31,223,31,36,31,17,31,145,31,173,31,106,31,217,31,27,31,236,31,72,31,72,30,72,29,41,31,219,31,66,31,66,30,194,31,189,31,189,30,217,31,43,31,117,31,180,31,162,31,118,31,62,31,4,31,128,31,128,30,47,31,77,31,13,31,240,31,255,31,10,31,83,31,83,30,178,31,207,31,221,31,97,31,97,30,67,31,40,31,40,30,182,31,173,31,218,31,29,31,67,31,237,31,237,30,210,31,243,31,10,31,193,31,117,31,14,31,14,30,32,31,211,31,211,30,161,31,52,31,251,31,204,31,91,31,91,30,240,31,74,31,93,31,43,31,248,31,197,31,173,31,214,31,96,31,216,31,216,30,3,31,142,31,136,31,44,31,70,31,103,31,216,31,98,31,98,30,8,31,244,31,172,31,251,31,99,31,221,31,103,31,103,30,137,31,108,31,102,31,140,31,91,31,91,30,91,31,96,31,245,31,99,31,99,30,7,31,161,31,200,31,192,31,155,31,240,31,232,31,43,31,44,31,44,30,44,29,44,28,255,31,29,31,184,31,235,31,20,31,67,31,147,31,102,31,157,31,215,31,43,31,54,31,79,31,137,31,96,31,25,31,45,31,111,31,165,31,165,30,250,31,113,31,113,30,249,31,22,31,117,31,135,31,192,31,21,31,72,31,160,31,134,31,35,31,167,31,48,31,150,31,93,31,220,31,155,31,155,30,6,31,182,31,150,31,191,31,191,30,222,31,222,30,253,31,253,30,221,31,134,31,224,31,224,30,224,29,245,31,243,31,240,31,228,31,151,31,15,31,231,31,93,31,52,31,164,31,205,31,205,30,85,31,22,31,247,31,247,30,43,31,158,31,245,31,114,31,65,31,112,31,251,31,251,30,251,29,234,31,234,30,65,31,28,31,28,30,93,31,12,31,119,31,119,30,64,31,64,30,214,31,41,31,41,30,119,31,168,31,113,31,216,31,48,31,254,31,140,31,132,31,139,31,166,31,249,31,249,30,240,31,240,30,216,31,202,31,195,31,169,31,169,30,56,31,193,31,75,31,235,31,235,30,235,29,204,31,35,31,129,31,102,31,230,31,38,31,38,30,38,29,66,31,66,30,160,31,137,31,221,31,61,31,239,31,239,30,128,31,192,31,192,30,192,29,41,31,41,30,219,31,219,30,73,31,81,31,81,30,81,29,45,31,132,31,32,31,138,31,202,31,198,31,198,30,96,31,77,31,255,31,246,31,246,30,246,29,241,31,53,31,19,31,5,31,131,31,50,31,214,31,214,30,47,31,222,31,222,30,40,31,19,31,85,31,85,30,99,31,77,31,243,31,243,30,235,31,68,31,68,30,190,31,13,31,149,31,149,30,152,31,12,31,12,31,225,31,249,31,22,31,97,31,237,31,49,31,49,30,236,31,236,30,56,31,33,31,146,31,181,31,122,31,220,31,109,31,191,31,252,31,81,31,246,31,246,30,233,31,63,31,122,31,248,31,199,31,199,30,168,31,123,31,215,31,181,31,74,31,159,31,25,31,29,31,200,31,135,31,2,31,156,31,17,31,205,31,200,31,249,31,107,31,79,31,192,31,139,31,254,31,255,31,120,31,111,31,150,31,88,31,134,31,134,30,210,31,210,30,210,29,210,28,210,27,242,31,127,31,231,31,129,31,3,31,65,31,97,31,192,31,71,31,141,31,237,31,237,30,237,29,237,28,18,31,167,31,135,31,135,30,194,31,200,31,111,31,111,30,163,31,254,31,27,31,27,30,27,29,61,31,225,31,49,31,12,31,12,30,39,31,148,31,62,31,145,31,141,31,136,31,35,31,96,31,192,31,67,31,255,31,255,30,154,31,48,31,48,30,216,31,177,31,130,31,158,31,58,31,58,30,242,31,230,31,244,31,106,31,139,31,27,31,57,31,115,31,228,31,28,31,254,31,254,30,186,31,155,31,212,31,222,31,222,30,218,31,89,31,180,31,180,30,247,31,247,30,154,31,158,31,227,31,184,31,12,31,61,31,172,31,98,31,173,31,76,31,76,30,76,29,30,31,129,31,139,31,118,31,229,31,229,31,61,31,61,30,224,31,209,31,209,31,209,30,45,31,45,30,168,31,164,31,16,31,183,31,99,31,218,31,218,30,36,31,164,31,189,31,71,31,173,31,173,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
