-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_516 is
end project_tb_516;

architecture project_tb_arch_516 of project_tb_516 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 300;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (4,0,178,0,0,0,62,0,0,0,149,0,187,0,25,0,123,0,200,0,125,0,154,0,110,0,211,0,0,0,0,0,31,0,21,0,150,0,54,0,192,0,71,0,188,0,97,0,247,0,161,0,0,0,216,0,0,0,0,0,222,0,183,0,89,0,126,0,205,0,141,0,55,0,100,0,146,0,0,0,0,0,66,0,214,0,223,0,135,0,140,0,0,0,185,0,254,0,243,0,0,0,3,0,242,0,183,0,162,0,76,0,112,0,102,0,0,0,96,0,194,0,117,0,96,0,0,0,224,0,131,0,0,0,101,0,29,0,160,0,80,0,126,0,152,0,0,0,0,0,60,0,246,0,176,0,36,0,118,0,43,0,200,0,36,0,153,0,111,0,0,0,55,0,20,0,157,0,0,0,5,0,125,0,250,0,0,0,123,0,192,0,169,0,30,0,44,0,63,0,138,0,60,0,192,0,188,0,232,0,90,0,0,0,250,0,46,0,238,0,238,0,76,0,187,0,217,0,154,0,212,0,238,0,223,0,244,0,50,0,170,0,39,0,179,0,0,0,237,0,42,0,189,0,82,0,174,0,53,0,0,0,235,0,193,0,33,0,142,0,228,0,0,0,0,0,217,0,242,0,236,0,227,0,147,0,45,0,224,0,11,0,106,0,217,0,68,0,0,0,209,0,187,0,180,0,247,0,131,0,0,0,36,0,105,0,49,0,192,0,89,0,147,0,155,0,0,0,44,0,75,0,124,0,21,0,0,0,0,0,39,0,15,0,222,0,0,0,0,0,176,0,119,0,190,0,185,0,0,0,223,0,14,0,95,0,224,0,185,0,0,0,109,0,200,0,0,0,226,0,192,0,203,0,146,0,108,0,183,0,150,0,229,0,0,0,164,0,146,0,0,0,43,0,13,0,0,0,250,0,0,0,0,0,124,0,91,0,102,0,0,0,110,0,44,0,64,0,252,0,44,0,181,0,76,0,24,0,31,0,8,0,0,0,225,0,84,0,31,0,158,0,29,0,130,0,0,0,232,0,176,0,253,0,13,0,103,0,18,0,120,0,162,0,60,0,183,0,181,0,139,0,62,0,108,0,102,0,12,0,47,0,0,0,7,0,123,0,55,0,100,0,0,0,0,0,210,0,138,0,133,0,148,0,131,0,227,0,0,0,0,0,78,0,229,0,96,0,0,0,162,0,193,0,171,0,122,0,0,0,215,0,111,0,243,0,161,0,45,0,225,0,66,0,48,0,20,0,0,0,152,0,74,0,0,0,51,0,66,0,0,0,248,0,0,0,82,0,20,0,0,0,66,0,104,0,208,0,73,0,152,0,152,0,162,0,52,0,214,0);
signal scenario_full  : scenario_type := (4,31,178,31,178,30,62,31,62,30,149,31,187,31,25,31,123,31,200,31,125,31,154,31,110,31,211,31,211,30,211,29,31,31,21,31,150,31,54,31,192,31,71,31,188,31,97,31,247,31,161,31,161,30,216,31,216,30,216,29,222,31,183,31,89,31,126,31,205,31,141,31,55,31,100,31,146,31,146,30,146,29,66,31,214,31,223,31,135,31,140,31,140,30,185,31,254,31,243,31,243,30,3,31,242,31,183,31,162,31,76,31,112,31,102,31,102,30,96,31,194,31,117,31,96,31,96,30,224,31,131,31,131,30,101,31,29,31,160,31,80,31,126,31,152,31,152,30,152,29,60,31,246,31,176,31,36,31,118,31,43,31,200,31,36,31,153,31,111,31,111,30,55,31,20,31,157,31,157,30,5,31,125,31,250,31,250,30,123,31,192,31,169,31,30,31,44,31,63,31,138,31,60,31,192,31,188,31,232,31,90,31,90,30,250,31,46,31,238,31,238,31,76,31,187,31,217,31,154,31,212,31,238,31,223,31,244,31,50,31,170,31,39,31,179,31,179,30,237,31,42,31,189,31,82,31,174,31,53,31,53,30,235,31,193,31,33,31,142,31,228,31,228,30,228,29,217,31,242,31,236,31,227,31,147,31,45,31,224,31,11,31,106,31,217,31,68,31,68,30,209,31,187,31,180,31,247,31,131,31,131,30,36,31,105,31,49,31,192,31,89,31,147,31,155,31,155,30,44,31,75,31,124,31,21,31,21,30,21,29,39,31,15,31,222,31,222,30,222,29,176,31,119,31,190,31,185,31,185,30,223,31,14,31,95,31,224,31,185,31,185,30,109,31,200,31,200,30,226,31,192,31,203,31,146,31,108,31,183,31,150,31,229,31,229,30,164,31,146,31,146,30,43,31,13,31,13,30,250,31,250,30,250,29,124,31,91,31,102,31,102,30,110,31,44,31,64,31,252,31,44,31,181,31,76,31,24,31,31,31,8,31,8,30,225,31,84,31,31,31,158,31,29,31,130,31,130,30,232,31,176,31,253,31,13,31,103,31,18,31,120,31,162,31,60,31,183,31,181,31,139,31,62,31,108,31,102,31,12,31,47,31,47,30,7,31,123,31,55,31,100,31,100,30,100,29,210,31,138,31,133,31,148,31,131,31,227,31,227,30,227,29,78,31,229,31,96,31,96,30,162,31,193,31,171,31,122,31,122,30,215,31,111,31,243,31,161,31,45,31,225,31,66,31,48,31,20,31,20,30,152,31,74,31,74,30,51,31,66,31,66,30,248,31,248,30,82,31,20,31,20,30,66,31,104,31,208,31,73,31,152,31,152,31,162,31,52,31,214,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
