-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 275;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (132,0,251,0,184,0,197,0,207,0,162,0,225,0,188,0,206,0,160,0,246,0,145,0,68,0,185,0,0,0,0,0,252,0,0,0,48,0,195,0,0,0,228,0,209,0,223,0,199,0,216,0,153,0,0,0,56,0,39,0,0,0,0,0,234,0,127,0,133,0,0,0,94,0,207,0,222,0,73,0,139,0,102,0,226,0,110,0,135,0,180,0,234,0,174,0,0,0,242,0,0,0,110,0,0,0,207,0,0,0,118,0,152,0,94,0,197,0,119,0,76,0,0,0,193,0,54,0,223,0,133,0,115,0,0,0,143,0,0,0,253,0,223,0,166,0,0,0,28,0,84,0,237,0,118,0,214,0,200,0,13,0,0,0,0,0,34,0,51,0,140,0,34,0,128,0,92,0,196,0,101,0,0,0,166,0,181,0,164,0,146,0,14,0,0,0,145,0,55,0,0,0,20,0,0,0,118,0,0,0,0,0,0,0,248,0,188,0,0,0,45,0,12,0,88,0,55,0,2,0,56,0,234,0,83,0,116,0,151,0,42,0,252,0,132,0,112,0,122,0,134,0,103,0,0,0,57,0,0,0,0,0,234,0,86,0,0,0,222,0,66,0,195,0,50,0,2,0,0,0,141,0,249,0,110,0,193,0,226,0,82,0,200,0,82,0,225,0,250,0,8,0,132,0,145,0,12,0,47,0,174,0,21,0,250,0,193,0,80,0,235,0,56,0,115,0,189,0,9,0,0,0,0,0,123,0,126,0,198,0,0,0,63,0,219,0,0,0,40,0,22,0,154,0,118,0,76,0,0,0,195,0,51,0,105,0,162,0,154,0,74,0,0,0,188,0,0,0,75,0,253,0,114,0,162,0,0,0,0,0,72,0,2,0,0,0,31,0,193,0,172,0,141,0,89,0,225,0,11,0,154,0,71,0,168,0,82,0,0,0,100,0,187,0,19,0,5,0,185,0,28,0,0,0,15,0,202,0,231,0,226,0,110,0,62,0,227,0,112,0,180,0,0,0,5,0,0,0,127,0,50,0,212,0,144,0,153,0,128,0,71,0,134,0,0,0,33,0,0,0,125,0,71,0,0,0,0,0,64,0,114,0,0,0,165,0,0,0,198,0,132,0,226,0,137,0,65,0,255,0,92,0,0,0,93,0,47,0,148,0,104,0,0,0,30,0,126,0,178,0,0,0,98,0,0,0,155,0,150,0,0,0,92,0,0,0,82,0,159,0);
signal scenario_full  : scenario_type := (132,31,251,31,184,31,197,31,207,31,162,31,225,31,188,31,206,31,160,31,246,31,145,31,68,31,185,31,185,30,185,29,252,31,252,30,48,31,195,31,195,30,228,31,209,31,223,31,199,31,216,31,153,31,153,30,56,31,39,31,39,30,39,29,234,31,127,31,133,31,133,30,94,31,207,31,222,31,73,31,139,31,102,31,226,31,110,31,135,31,180,31,234,31,174,31,174,30,242,31,242,30,110,31,110,30,207,31,207,30,118,31,152,31,94,31,197,31,119,31,76,31,76,30,193,31,54,31,223,31,133,31,115,31,115,30,143,31,143,30,253,31,223,31,166,31,166,30,28,31,84,31,237,31,118,31,214,31,200,31,13,31,13,30,13,29,34,31,51,31,140,31,34,31,128,31,92,31,196,31,101,31,101,30,166,31,181,31,164,31,146,31,14,31,14,30,145,31,55,31,55,30,20,31,20,30,118,31,118,30,118,29,118,28,248,31,188,31,188,30,45,31,12,31,88,31,55,31,2,31,56,31,234,31,83,31,116,31,151,31,42,31,252,31,132,31,112,31,122,31,134,31,103,31,103,30,57,31,57,30,57,29,234,31,86,31,86,30,222,31,66,31,195,31,50,31,2,31,2,30,141,31,249,31,110,31,193,31,226,31,82,31,200,31,82,31,225,31,250,31,8,31,132,31,145,31,12,31,47,31,174,31,21,31,250,31,193,31,80,31,235,31,56,31,115,31,189,31,9,31,9,30,9,29,123,31,126,31,198,31,198,30,63,31,219,31,219,30,40,31,22,31,154,31,118,31,76,31,76,30,195,31,51,31,105,31,162,31,154,31,74,31,74,30,188,31,188,30,75,31,253,31,114,31,162,31,162,30,162,29,72,31,2,31,2,30,31,31,193,31,172,31,141,31,89,31,225,31,11,31,154,31,71,31,168,31,82,31,82,30,100,31,187,31,19,31,5,31,185,31,28,31,28,30,15,31,202,31,231,31,226,31,110,31,62,31,227,31,112,31,180,31,180,30,5,31,5,30,127,31,50,31,212,31,144,31,153,31,128,31,71,31,134,31,134,30,33,31,33,30,125,31,71,31,71,30,71,29,64,31,114,31,114,30,165,31,165,30,198,31,132,31,226,31,137,31,65,31,255,31,92,31,92,30,93,31,47,31,148,31,104,31,104,30,30,31,126,31,178,31,178,30,98,31,98,30,155,31,150,31,150,30,92,31,92,30,82,31,159,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
