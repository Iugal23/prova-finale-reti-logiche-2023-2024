-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_327 is
end project_tb_327;

architecture project_tb_arch_327 of project_tb_327 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 974;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (254,0,65,0,228,0,197,0,204,0,22,0,154,0,146,0,0,0,107,0,196,0,7,0,146,0,0,0,143,0,141,0,180,0,20,0,157,0,20,0,81,0,115,0,45,0,140,0,11,0,229,0,0,0,42,0,19,0,14,0,146,0,0,0,149,0,0,0,118,0,182,0,0,0,157,0,57,0,243,0,150,0,32,0,44,0,222,0,44,0,32,0,161,0,65,0,0,0,0,0,220,0,100,0,183,0,0,0,0,0,0,0,0,0,53,0,53,0,235,0,171,0,72,0,23,0,199,0,0,0,42,0,240,0,0,0,0,0,248,0,62,0,0,0,217,0,9,0,67,0,209,0,80,0,126,0,0,0,12,0,16,0,163,0,161,0,0,0,75,0,236,0,184,0,76,0,11,0,121,0,176,0,119,0,181,0,33,0,226,0,40,0,0,0,246,0,150,0,160,0,199,0,39,0,66,0,21,0,221,0,26,0,141,0,24,0,0,0,192,0,106,0,209,0,107,0,0,0,238,0,0,0,189,0,77,0,184,0,82,0,167,0,235,0,1,0,48,0,208,0,198,0,152,0,243,0,195,0,0,0,140,0,11,0,152,0,156,0,173,0,127,0,96,0,166,0,40,0,0,0,40,0,10,0,128,0,163,0,49,0,230,0,213,0,164,0,0,0,226,0,169,0,144,0,190,0,199,0,156,0,246,0,238,0,0,0,237,0,66,0,0,0,70,0,192,0,71,0,0,0,41,0,126,0,140,0,147,0,130,0,48,0,14,0,172,0,27,0,8,0,195,0,143,0,2,0,46,0,31,0,142,0,175,0,55,0,37,0,100,0,110,0,0,0,142,0,106,0,48,0,43,0,241,0,25,0,156,0,0,0,0,0,0,0,0,0,23,0,220,0,83,0,149,0,4,0,21,0,148,0,47,0,237,0,0,0,0,0,68,0,140,0,165,0,109,0,5,0,38,0,192,0,74,0,9,0,215,0,0,0,168,0,255,0,0,0,0,0,249,0,125,0,88,0,237,0,29,0,0,0,59,0,0,0,253,0,183,0,34,0,251,0,0,0,26,0,85,0,151,0,199,0,0,0,243,0,111,0,66,0,0,0,160,0,225,0,201,0,0,0,156,0,0,0,219,0,6,0,73,0,251,0,113,0,179,0,0,0,175,0,155,0,169,0,162,0,189,0,0,0,168,0,0,0,30,0,67,0,8,0,83,0,0,0,112,0,130,0,73,0,0,0,252,0,101,0,0,0,171,0,103,0,50,0,0,0,0,0,0,0,0,0,180,0,43,0,174,0,162,0,173,0,0,0,176,0,0,0,106,0,184,0,253,0,189,0,0,0,30,0,65,0,214,0,106,0,80,0,151,0,68,0,63,0,0,0,164,0,171,0,34,0,38,0,220,0,132,0,72,0,3,0,52,0,0,0,108,0,80,0,142,0,251,0,79,0,36,0,45,0,111,0,24,0,207,0,240,0,151,0,232,0,0,0,199,0,44,0,134,0,198,0,0,0,168,0,218,0,250,0,75,0,9,0,143,0,241,0,119,0,249,0,219,0,0,0,8,0,243,0,48,0,0,0,216,0,0,0,0,0,227,0,237,0,220,0,209,0,72,0,27,0,31,0,166,0,161,0,15,0,0,0,185,0,212,0,245,0,70,0,236,0,245,0,239,0,0,0,0,0,64,0,94,0,0,0,77,0,224,0,138,0,165,0,30,0,0,0,79,0,76,0,0,0,72,0,172,0,4,0,80,0,80,0,168,0,134,0,10,0,188,0,68,0,220,0,0,0,55,0,57,0,0,0,59,0,67,0,0,0,237,0,60,0,0,0,0,0,30,0,254,0,91,0,135,0,0,0,116,0,235,0,0,0,0,0,220,0,31,0,62,0,169,0,169,0,152,0,6,0,179,0,250,0,175,0,218,0,233,0,54,0,14,0,91,0,148,0,30,0,0,0,140,0,246,0,88,0,0,0,109,0,0,0,0,0,200,0,236,0,123,0,238,0,80,0,202,0,254,0,112,0,138,0,144,0,153,0,61,0,129,0,0,0,61,0,224,0,80,0,16,0,44,0,224,0,111,0,156,0,43,0,252,0,0,0,204,0,36,0,1,0,62,0,243,0,107,0,240,0,0,0,0,0,78,0,182,0,167,0,60,0,14,0,129,0,234,0,100,0,210,0,26,0,132,0,27,0,0,0,10,0,90,0,200,0,15,0,0,0,11,0,142,0,4,0,0,0,0,0,230,0,78,0,89,0,202,0,135,0,50,0,0,0,208,0,215,0,209,0,12,0,17,0,0,0,162,0,47,0,138,0,175,0,185,0,0,0,56,0,35,0,138,0,35,0,120,0,0,0,193,0,57,0,150,0,94,0,92,0,3,0,0,0,96,0,115,0,126,0,4,0,3,0,185,0,240,0,0,0,0,0,93,0,229,0,0,0,14,0,169,0,108,0,138,0,10,0,115,0,9,0,0,0,102,0,104,0,0,0,222,0,95,0,245,0,131,0,112,0,160,0,26,0,0,0,159,0,100,0,0,0,89,0,0,0,0,0,0,0,182,0,84,0,194,0,0,0,109,0,178,0,0,0,219,0,148,0,158,0,26,0,140,0,148,0,43,0,162,0,0,0,155,0,151,0,150,0,157,0,139,0,222,0,35,0,7,0,0,0,159,0,1,0,0,0,144,0,0,0,20,0,36,0,200,0,71,0,151,0,247,0,0,0,39,0,224,0,204,0,197,0,0,0,37,0,31,0,0,0,52,0,91,0,142,0,126,0,82,0,238,0,57,0,102,0,107,0,10,0,0,0,31,0,253,0,13,0,192,0,141,0,0,0,76,0,69,0,0,0,152,0,55,0,0,0,0,0,69,0,46,0,0,0,247,0,0,0,239,0,40,0,195,0,83,0,238,0,206,0,191,0,214,0,0,0,5,0,139,0,222,0,136,0,2,0,138,0,148,0,0,0,0,0,220,0,213,0,51,0,71,0,102,0,0,0,32,0,0,0,199,0,55,0,0,0,80,0,84,0,158,0,164,0,0,0,131,0,235,0,215,0,94,0,3,0,84,0,0,0,0,0,0,0,29,0,0,0,82,0,13,0,174,0,187,0,0,0,96,0,31,0,10,0,0,0,251,0,75,0,226,0,0,0,70,0,41,0,44,0,113,0,183,0,39,0,248,0,210,0,0,0,119,0,247,0,0,0,148,0,0,0,173,0,61,0,0,0,212,0,0,0,77,0,135,0,87,0,126,0,165,0,85,0,0,0,0,0,235,0,138,0,0,0,163,0,105,0,146,0,193,0,182,0,81,0,251,0,139,0,106,0,234,0,12,0,124,0,192,0,11,0,109,0,33,0,185,0,45,0,160,0,30,0,18,0,31,0,143,0,254,0,95,0,0,0,62,0,0,0,106,0,0,0,53,0,0,0,165,0,210,0,0,0,22,0,227,0,9,0,99,0,244,0,69,0,93,0,89,0,41,0,220,0,73,0,200,0,201,0,172,0,103,0,228,0,0,0,146,0,67,0,243,0,22,0,135,0,0,0,48,0,46,0,0,0,128,0,0,0,238,0,0,0,176,0,0,0,99,0,0,0,94,0,233,0,45,0,149,0,139,0,247,0,95,0,75,0,0,0,31,0,28,0,93,0,29,0,37,0,20,0,104,0,0,0,158,0,255,0,233,0,73,0,0,0,133,0,0,0,138,0,0,0,0,0,154,0,79,0,98,0,59,0,237,0,16,0,172,0,232,0,237,0,27,0,14,0,76,0,144,0,119,0,248,0,34,0,140,0,0,0,59,0,238,0,191,0,19,0,143,0,0,0,95,0,59,0,127,0,0,0,223,0,229,0,142,0,209,0,171,0,140,0,228,0,0,0,55,0,109,0,251,0,169,0,0,0,197,0,206,0,0,0,207,0,0,0,23,0,9,0,208,0,185,0,147,0,246,0,0,0,138,0,224,0,48,0,161,0,211,0,155,0,113,0,178,0,51,0,0,0,159,0,7,0,129,0,0,0,0,0,54,0,250,0,152,0,0,0,159,0,1,0,200,0,245,0,248,0,0,0,193,0,255,0,175,0,0,0,252,0,7,0,0,0,47,0,0,0,0,0,103,0,12,0,71,0,65,0,0,0,109,0,61,0,163,0,0,0,85,0,0,0,223,0,165,0,148,0,0,0,86,0,25,0,0,0,163,0,206,0,18,0,35,0,0,0,0,0,36,0,206,0,0,0,169,0,44,0,247,0,76,0,140,0,155,0,103,0,234,0,66,0,87,0,127,0,18,0,108,0,219,0,81,0,0,0,179,0,118,0,17,0,57,0,39,0,0,0,204,0,4,0,144,0,85,0,0,0,237,0,0,0,103,0,206,0);
signal scenario_full  : scenario_type := (254,31,65,31,228,31,197,31,204,31,22,31,154,31,146,31,146,30,107,31,196,31,7,31,146,31,146,30,143,31,141,31,180,31,20,31,157,31,20,31,81,31,115,31,45,31,140,31,11,31,229,31,229,30,42,31,19,31,14,31,146,31,146,30,149,31,149,30,118,31,182,31,182,30,157,31,57,31,243,31,150,31,32,31,44,31,222,31,44,31,32,31,161,31,65,31,65,30,65,29,220,31,100,31,183,31,183,30,183,29,183,28,183,27,53,31,53,31,235,31,171,31,72,31,23,31,199,31,199,30,42,31,240,31,240,30,240,29,248,31,62,31,62,30,217,31,9,31,67,31,209,31,80,31,126,31,126,30,12,31,16,31,163,31,161,31,161,30,75,31,236,31,184,31,76,31,11,31,121,31,176,31,119,31,181,31,33,31,226,31,40,31,40,30,246,31,150,31,160,31,199,31,39,31,66,31,21,31,221,31,26,31,141,31,24,31,24,30,192,31,106,31,209,31,107,31,107,30,238,31,238,30,189,31,77,31,184,31,82,31,167,31,235,31,1,31,48,31,208,31,198,31,152,31,243,31,195,31,195,30,140,31,11,31,152,31,156,31,173,31,127,31,96,31,166,31,40,31,40,30,40,31,10,31,128,31,163,31,49,31,230,31,213,31,164,31,164,30,226,31,169,31,144,31,190,31,199,31,156,31,246,31,238,31,238,30,237,31,66,31,66,30,70,31,192,31,71,31,71,30,41,31,126,31,140,31,147,31,130,31,48,31,14,31,172,31,27,31,8,31,195,31,143,31,2,31,46,31,31,31,142,31,175,31,55,31,37,31,100,31,110,31,110,30,142,31,106,31,48,31,43,31,241,31,25,31,156,31,156,30,156,29,156,28,156,27,23,31,220,31,83,31,149,31,4,31,21,31,148,31,47,31,237,31,237,30,237,29,68,31,140,31,165,31,109,31,5,31,38,31,192,31,74,31,9,31,215,31,215,30,168,31,255,31,255,30,255,29,249,31,125,31,88,31,237,31,29,31,29,30,59,31,59,30,253,31,183,31,34,31,251,31,251,30,26,31,85,31,151,31,199,31,199,30,243,31,111,31,66,31,66,30,160,31,225,31,201,31,201,30,156,31,156,30,219,31,6,31,73,31,251,31,113,31,179,31,179,30,175,31,155,31,169,31,162,31,189,31,189,30,168,31,168,30,30,31,67,31,8,31,83,31,83,30,112,31,130,31,73,31,73,30,252,31,101,31,101,30,171,31,103,31,50,31,50,30,50,29,50,28,50,27,180,31,43,31,174,31,162,31,173,31,173,30,176,31,176,30,106,31,184,31,253,31,189,31,189,30,30,31,65,31,214,31,106,31,80,31,151,31,68,31,63,31,63,30,164,31,171,31,34,31,38,31,220,31,132,31,72,31,3,31,52,31,52,30,108,31,80,31,142,31,251,31,79,31,36,31,45,31,111,31,24,31,207,31,240,31,151,31,232,31,232,30,199,31,44,31,134,31,198,31,198,30,168,31,218,31,250,31,75,31,9,31,143,31,241,31,119,31,249,31,219,31,219,30,8,31,243,31,48,31,48,30,216,31,216,30,216,29,227,31,237,31,220,31,209,31,72,31,27,31,31,31,166,31,161,31,15,31,15,30,185,31,212,31,245,31,70,31,236,31,245,31,239,31,239,30,239,29,64,31,94,31,94,30,77,31,224,31,138,31,165,31,30,31,30,30,79,31,76,31,76,30,72,31,172,31,4,31,80,31,80,31,168,31,134,31,10,31,188,31,68,31,220,31,220,30,55,31,57,31,57,30,59,31,67,31,67,30,237,31,60,31,60,30,60,29,30,31,254,31,91,31,135,31,135,30,116,31,235,31,235,30,235,29,220,31,31,31,62,31,169,31,169,31,152,31,6,31,179,31,250,31,175,31,218,31,233,31,54,31,14,31,91,31,148,31,30,31,30,30,140,31,246,31,88,31,88,30,109,31,109,30,109,29,200,31,236,31,123,31,238,31,80,31,202,31,254,31,112,31,138,31,144,31,153,31,61,31,129,31,129,30,61,31,224,31,80,31,16,31,44,31,224,31,111,31,156,31,43,31,252,31,252,30,204,31,36,31,1,31,62,31,243,31,107,31,240,31,240,30,240,29,78,31,182,31,167,31,60,31,14,31,129,31,234,31,100,31,210,31,26,31,132,31,27,31,27,30,10,31,90,31,200,31,15,31,15,30,11,31,142,31,4,31,4,30,4,29,230,31,78,31,89,31,202,31,135,31,50,31,50,30,208,31,215,31,209,31,12,31,17,31,17,30,162,31,47,31,138,31,175,31,185,31,185,30,56,31,35,31,138,31,35,31,120,31,120,30,193,31,57,31,150,31,94,31,92,31,3,31,3,30,96,31,115,31,126,31,4,31,3,31,185,31,240,31,240,30,240,29,93,31,229,31,229,30,14,31,169,31,108,31,138,31,10,31,115,31,9,31,9,30,102,31,104,31,104,30,222,31,95,31,245,31,131,31,112,31,160,31,26,31,26,30,159,31,100,31,100,30,89,31,89,30,89,29,89,28,182,31,84,31,194,31,194,30,109,31,178,31,178,30,219,31,148,31,158,31,26,31,140,31,148,31,43,31,162,31,162,30,155,31,151,31,150,31,157,31,139,31,222,31,35,31,7,31,7,30,159,31,1,31,1,30,144,31,144,30,20,31,36,31,200,31,71,31,151,31,247,31,247,30,39,31,224,31,204,31,197,31,197,30,37,31,31,31,31,30,52,31,91,31,142,31,126,31,82,31,238,31,57,31,102,31,107,31,10,31,10,30,31,31,253,31,13,31,192,31,141,31,141,30,76,31,69,31,69,30,152,31,55,31,55,30,55,29,69,31,46,31,46,30,247,31,247,30,239,31,40,31,195,31,83,31,238,31,206,31,191,31,214,31,214,30,5,31,139,31,222,31,136,31,2,31,138,31,148,31,148,30,148,29,220,31,213,31,51,31,71,31,102,31,102,30,32,31,32,30,199,31,55,31,55,30,80,31,84,31,158,31,164,31,164,30,131,31,235,31,215,31,94,31,3,31,84,31,84,30,84,29,84,28,29,31,29,30,82,31,13,31,174,31,187,31,187,30,96,31,31,31,10,31,10,30,251,31,75,31,226,31,226,30,70,31,41,31,44,31,113,31,183,31,39,31,248,31,210,31,210,30,119,31,247,31,247,30,148,31,148,30,173,31,61,31,61,30,212,31,212,30,77,31,135,31,87,31,126,31,165,31,85,31,85,30,85,29,235,31,138,31,138,30,163,31,105,31,146,31,193,31,182,31,81,31,251,31,139,31,106,31,234,31,12,31,124,31,192,31,11,31,109,31,33,31,185,31,45,31,160,31,30,31,18,31,31,31,143,31,254,31,95,31,95,30,62,31,62,30,106,31,106,30,53,31,53,30,165,31,210,31,210,30,22,31,227,31,9,31,99,31,244,31,69,31,93,31,89,31,41,31,220,31,73,31,200,31,201,31,172,31,103,31,228,31,228,30,146,31,67,31,243,31,22,31,135,31,135,30,48,31,46,31,46,30,128,31,128,30,238,31,238,30,176,31,176,30,99,31,99,30,94,31,233,31,45,31,149,31,139,31,247,31,95,31,75,31,75,30,31,31,28,31,93,31,29,31,37,31,20,31,104,31,104,30,158,31,255,31,233,31,73,31,73,30,133,31,133,30,138,31,138,30,138,29,154,31,79,31,98,31,59,31,237,31,16,31,172,31,232,31,237,31,27,31,14,31,76,31,144,31,119,31,248,31,34,31,140,31,140,30,59,31,238,31,191,31,19,31,143,31,143,30,95,31,59,31,127,31,127,30,223,31,229,31,142,31,209,31,171,31,140,31,228,31,228,30,55,31,109,31,251,31,169,31,169,30,197,31,206,31,206,30,207,31,207,30,23,31,9,31,208,31,185,31,147,31,246,31,246,30,138,31,224,31,48,31,161,31,211,31,155,31,113,31,178,31,51,31,51,30,159,31,7,31,129,31,129,30,129,29,54,31,250,31,152,31,152,30,159,31,1,31,200,31,245,31,248,31,248,30,193,31,255,31,175,31,175,30,252,31,7,31,7,30,47,31,47,30,47,29,103,31,12,31,71,31,65,31,65,30,109,31,61,31,163,31,163,30,85,31,85,30,223,31,165,31,148,31,148,30,86,31,25,31,25,30,163,31,206,31,18,31,35,31,35,30,35,29,36,31,206,31,206,30,169,31,44,31,247,31,76,31,140,31,155,31,103,31,234,31,66,31,87,31,127,31,18,31,108,31,219,31,81,31,81,30,179,31,118,31,17,31,57,31,39,31,39,30,204,31,4,31,144,31,85,31,85,30,237,31,237,30,103,31,206,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
