-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 922;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (150,0,0,0,199,0,100,0,246,0,21,0,60,0,63,0,0,0,244,0,0,0,207,0,231,0,156,0,0,0,241,0,14,0,0,0,49,0,94,0,97,0,82,0,144,0,34,0,227,0,40,0,0,0,92,0,0,0,218,0,145,0,119,0,245,0,198,0,83,0,195,0,233,0,247,0,45,0,1,0,0,0,222,0,0,0,0,0,102,0,97,0,27,0,97,0,16,0,255,0,86,0,212,0,119,0,88,0,0,0,32,0,153,0,55,0,0,0,62,0,0,0,2,0,24,0,42,0,206,0,0,0,9,0,0,0,0,0,6,0,194,0,31,0,113,0,0,0,20,0,181,0,69,0,52,0,0,0,78,0,27,0,160,0,243,0,101,0,178,0,149,0,35,0,0,0,211,0,154,0,167,0,173,0,126,0,78,0,0,0,220,0,158,0,221,0,117,0,108,0,29,0,250,0,243,0,171,0,201,0,7,0,242,0,0,0,36,0,111,0,0,0,107,0,84,0,4,0,137,0,235,0,24,0,0,0,62,0,0,0,227,0,92,0,0,0,125,0,149,0,0,0,72,0,45,0,0,0,0,0,151,0,152,0,167,0,0,0,121,0,14,0,50,0,10,0,85,0,125,0,130,0,0,0,244,0,167,0,224,0,50,0,95,0,197,0,112,0,82,0,110,0,196,0,11,0,94,0,19,0,0,0,134,0,20,0,149,0,99,0,207,0,0,0,19,0,54,0,31,0,255,0,69,0,0,0,0,0,15,0,58,0,245,0,0,0,171,0,182,0,92,0,0,0,247,0,174,0,144,0,160,0,232,0,171,0,175,0,0,0,11,0,247,0,236,0,0,0,8,0,156,0,144,0,127,0,163,0,0,0,0,0,170,0,190,0,85,0,249,0,114,0,95,0,54,0,0,0,117,0,93,0,0,0,104,0,0,0,58,0,47,0,0,0,4,0,85,0,198,0,165,0,187,0,142,0,46,0,0,0,142,0,144,0,68,0,11,0,203,0,0,0,184,0,0,0,124,0,85,0,238,0,152,0,115,0,21,0,0,0,129,0,179,0,64,0,231,0,169,0,111,0,0,0,93,0,88,0,76,0,235,0,0,0,168,0,211,0,57,0,0,0,235,0,234,0,252,0,62,0,90,0,255,0,0,0,79,0,232,0,9,0,231,0,232,0,0,0,182,0,0,0,0,0,125,0,55,0,0,0,0,0,145,0,59,0,77,0,191,0,193,0,0,0,0,0,0,0,207,0,149,0,70,0,224,0,197,0,25,0,196,0,58,0,0,0,245,0,20,0,40,0,58,0,39,0,118,0,163,0,93,0,16,0,3,0,112,0,0,0,127,0,207,0,97,0,204,0,110,0,252,0,169,0,42,0,87,0,37,0,0,0,148,0,0,0,37,0,40,0,200,0,0,0,0,0,0,0,0,0,0,0,209,0,179,0,22,0,99,0,158,0,243,0,0,0,92,0,209,0,44,0,0,0,0,0,63,0,0,0,100,0,14,0,137,0,49,0,0,0,77,0,189,0,111,0,91,0,146,0,107,0,62,0,0,0,35,0,21,0,141,0,255,0,222,0,0,0,0,0,77,0,83,0,37,0,214,0,71,0,194,0,28,0,218,0,72,0,231,0,191,0,164,0,193,0,193,0,204,0,70,0,89,0,75,0,97,0,0,0,20,0,87,0,0,0,216,0,129,0,226,0,95,0,0,0,0,0,17,0,5,0,48,0,184,0,89,0,0,0,103,0,0,0,14,0,89,0,141,0,29,0,72,0,100,0,128,0,172,0,0,0,223,0,49,0,92,0,103,0,0,0,75,0,137,0,251,0,39,0,0,0,148,0,114,0,214,0,216,0,0,0,250,0,251,0,143,0,33,0,0,0,93,0,0,0,248,0,96,0,0,0,196,0,213,0,149,0,131,0,160,0,132,0,78,0,183,0,227,0,208,0,98,0,0,0,131,0,30,0,204,0,156,0,178,0,23,0,94,0,0,0,223,0,70,0,165,0,220,0,164,0,34,0,36,0,116,0,51,0,0,0,115,0,139,0,161,0,143,0,69,0,153,0,159,0,4,0,82,0,248,0,207,0,22,0,0,0,116,0,197,0,28,0,30,0,0,0,42,0,108,0,42,0,0,0,172,0,194,0,76,0,167,0,245,0,153,0,162,0,0,0,0,0,0,0,0,0,20,0,66,0,143,0,0,0,179,0,236,0,152,0,178,0,93,0,1,0,139,0,230,0,0,0,0,0,81,0,146,0,38,0,255,0,248,0,94,0,125,0,31,0,205,0,213,0,12,0,42,0,193,0,4,0,148,0,199,0,0,0,0,0,107,0,0,0,0,0,0,0,120,0,86,0,198,0,72,0,147,0,210,0,141,0,19,0,204,0,53,0,75,0,0,0,22,0,0,0,148,0,242,0,3,0,186,0,0,0,108,0,96,0,161,0,72,0,3,0,223,0,0,0,243,0,134,0,0,0,0,0,90,0,80,0,97,0,207,0,0,0,0,0,53,0,121,0,62,0,13,0,112,0,240,0,45,0,42,0,50,0,9,0,33,0,244,0,94,0,0,0,225,0,48,0,21,0,203,0,83,0,31,0,201,0,131,0,0,0,222,0,178,0,145,0,0,0,20,0,161,0,158,0,196,0,91,0,137,0,0,0,174,0,145,0,247,0,0,0,241,0,153,0,10,0,30,0,31,0,220,0,0,0,27,0,25,0,161,0,0,0,3,0,0,0,0,0,159,0,0,0,217,0,2,0,230,0,0,0,212,0,190,0,95,0,147,0,176,0,113,0,202,0,130,0,185,0,86,0,110,0,99,0,235,0,96,0,198,0,191,0,207,0,87,0,0,0,135,0,228,0,254,0,179,0,120,0,211,0,231,0,59,0,12,0,53,0,235,0,140,0,10,0,0,0,84,0,0,0,247,0,0,0,0,0,240,0,0,0,140,0,28,0,190,0,214,0,191,0,0,0,0,0,99,0,197,0,57,0,148,0,0,0,132,0,150,0,198,0,25,0,209,0,0,0,0,0,26,0,117,0,0,0,85,0,5,0,18,0,0,0,68,0,127,0,187,0,0,0,210,0,204,0,54,0,214,0,137,0,0,0,205,0,234,0,211,0,183,0,59,0,252,0,40,0,248,0,96,0,130,0,0,0,158,0,0,0,19,0,21,0,47,0,141,0,147,0,108,0,0,0,206,0,25,0,0,0,162,0,0,0,230,0,107,0,108,0,137,0,0,0,148,0,181,0,0,0,85,0,110,0,0,0,238,0,125,0,179,0,56,0,193,0,118,0,82,0,202,0,111,0,252,0,140,0,0,0,7,0,118,0,136,0,124,0,78,0,95,0,147,0,168,0,26,0,5,0,246,0,12,0,41,0,0,0,174,0,86,0,183,0,102,0,242,0,207,0,220,0,87,0,0,0,244,0,225,0,84,0,159,0,6,0,0,0,0,0,198,0,69,0,32,0,71,0,207,0,122,0,230,0,51,0,225,0,173,0,170,0,1,0,186,0,0,0,202,0,202,0,0,0,135,0,204,0,148,0,158,0,45,0,65,0,196,0,216,0,6,0,113,0,249,0,173,0,98,0,0,0,159,0,73,0,241,0,197,0,121,0,140,0,218,0,185,0,103,0,103,0,48,0,178,0,164,0,0,0,113,0,200,0,116,0,229,0,0,0,0,0,0,0,205,0,106,0,148,0,0,0,80,0,180,0,255,0,212,0,234,0,17,0,0,0,173,0,241,0,204,0,119,0,225,0,0,0,135,0,155,0,0,0,224,0,125,0,249,0,107,0,2,0,129,0,204,0,172,0,64,0,101,0,214,0,0,0,166,0,15,0,225,0,199,0,133,0,141,0,182,0,107,0,136,0,27,0,224,0,98,0,0,0,239,0,68,0,93,0,0,0,0,0,0,0,75,0,139,0,124,0,215,0,0,0,56,0,45,0,0,0,180,0,0,0,28,0,134,0,0,0,52,0,135,0,65,0,0,0,140,0,207,0,0,0,202,0,232,0,92,0,193,0,0,0,194,0,0,0,0,0,0,0,79,0,18,0,225,0,232,0,97,0,78,0,0,0,121,0,165,0,0,0,231,0,80,0,39,0,58,0,34,0,107,0,22,0);
signal scenario_full  : scenario_type := (150,31,150,30,199,31,100,31,246,31,21,31,60,31,63,31,63,30,244,31,244,30,207,31,231,31,156,31,156,30,241,31,14,31,14,30,49,31,94,31,97,31,82,31,144,31,34,31,227,31,40,31,40,30,92,31,92,30,218,31,145,31,119,31,245,31,198,31,83,31,195,31,233,31,247,31,45,31,1,31,1,30,222,31,222,30,222,29,102,31,97,31,27,31,97,31,16,31,255,31,86,31,212,31,119,31,88,31,88,30,32,31,153,31,55,31,55,30,62,31,62,30,2,31,24,31,42,31,206,31,206,30,9,31,9,30,9,29,6,31,194,31,31,31,113,31,113,30,20,31,181,31,69,31,52,31,52,30,78,31,27,31,160,31,243,31,101,31,178,31,149,31,35,31,35,30,211,31,154,31,167,31,173,31,126,31,78,31,78,30,220,31,158,31,221,31,117,31,108,31,29,31,250,31,243,31,171,31,201,31,7,31,242,31,242,30,36,31,111,31,111,30,107,31,84,31,4,31,137,31,235,31,24,31,24,30,62,31,62,30,227,31,92,31,92,30,125,31,149,31,149,30,72,31,45,31,45,30,45,29,151,31,152,31,167,31,167,30,121,31,14,31,50,31,10,31,85,31,125,31,130,31,130,30,244,31,167,31,224,31,50,31,95,31,197,31,112,31,82,31,110,31,196,31,11,31,94,31,19,31,19,30,134,31,20,31,149,31,99,31,207,31,207,30,19,31,54,31,31,31,255,31,69,31,69,30,69,29,15,31,58,31,245,31,245,30,171,31,182,31,92,31,92,30,247,31,174,31,144,31,160,31,232,31,171,31,175,31,175,30,11,31,247,31,236,31,236,30,8,31,156,31,144,31,127,31,163,31,163,30,163,29,170,31,190,31,85,31,249,31,114,31,95,31,54,31,54,30,117,31,93,31,93,30,104,31,104,30,58,31,47,31,47,30,4,31,85,31,198,31,165,31,187,31,142,31,46,31,46,30,142,31,144,31,68,31,11,31,203,31,203,30,184,31,184,30,124,31,85,31,238,31,152,31,115,31,21,31,21,30,129,31,179,31,64,31,231,31,169,31,111,31,111,30,93,31,88,31,76,31,235,31,235,30,168,31,211,31,57,31,57,30,235,31,234,31,252,31,62,31,90,31,255,31,255,30,79,31,232,31,9,31,231,31,232,31,232,30,182,31,182,30,182,29,125,31,55,31,55,30,55,29,145,31,59,31,77,31,191,31,193,31,193,30,193,29,193,28,207,31,149,31,70,31,224,31,197,31,25,31,196,31,58,31,58,30,245,31,20,31,40,31,58,31,39,31,118,31,163,31,93,31,16,31,3,31,112,31,112,30,127,31,207,31,97,31,204,31,110,31,252,31,169,31,42,31,87,31,37,31,37,30,148,31,148,30,37,31,40,31,200,31,200,30,200,29,200,28,200,27,200,26,209,31,179,31,22,31,99,31,158,31,243,31,243,30,92,31,209,31,44,31,44,30,44,29,63,31,63,30,100,31,14,31,137,31,49,31,49,30,77,31,189,31,111,31,91,31,146,31,107,31,62,31,62,30,35,31,21,31,141,31,255,31,222,31,222,30,222,29,77,31,83,31,37,31,214,31,71,31,194,31,28,31,218,31,72,31,231,31,191,31,164,31,193,31,193,31,204,31,70,31,89,31,75,31,97,31,97,30,20,31,87,31,87,30,216,31,129,31,226,31,95,31,95,30,95,29,17,31,5,31,48,31,184,31,89,31,89,30,103,31,103,30,14,31,89,31,141,31,29,31,72,31,100,31,128,31,172,31,172,30,223,31,49,31,92,31,103,31,103,30,75,31,137,31,251,31,39,31,39,30,148,31,114,31,214,31,216,31,216,30,250,31,251,31,143,31,33,31,33,30,93,31,93,30,248,31,96,31,96,30,196,31,213,31,149,31,131,31,160,31,132,31,78,31,183,31,227,31,208,31,98,31,98,30,131,31,30,31,204,31,156,31,178,31,23,31,94,31,94,30,223,31,70,31,165,31,220,31,164,31,34,31,36,31,116,31,51,31,51,30,115,31,139,31,161,31,143,31,69,31,153,31,159,31,4,31,82,31,248,31,207,31,22,31,22,30,116,31,197,31,28,31,30,31,30,30,42,31,108,31,42,31,42,30,172,31,194,31,76,31,167,31,245,31,153,31,162,31,162,30,162,29,162,28,162,27,20,31,66,31,143,31,143,30,179,31,236,31,152,31,178,31,93,31,1,31,139,31,230,31,230,30,230,29,81,31,146,31,38,31,255,31,248,31,94,31,125,31,31,31,205,31,213,31,12,31,42,31,193,31,4,31,148,31,199,31,199,30,199,29,107,31,107,30,107,29,107,28,120,31,86,31,198,31,72,31,147,31,210,31,141,31,19,31,204,31,53,31,75,31,75,30,22,31,22,30,148,31,242,31,3,31,186,31,186,30,108,31,96,31,161,31,72,31,3,31,223,31,223,30,243,31,134,31,134,30,134,29,90,31,80,31,97,31,207,31,207,30,207,29,53,31,121,31,62,31,13,31,112,31,240,31,45,31,42,31,50,31,9,31,33,31,244,31,94,31,94,30,225,31,48,31,21,31,203,31,83,31,31,31,201,31,131,31,131,30,222,31,178,31,145,31,145,30,20,31,161,31,158,31,196,31,91,31,137,31,137,30,174,31,145,31,247,31,247,30,241,31,153,31,10,31,30,31,31,31,220,31,220,30,27,31,25,31,161,31,161,30,3,31,3,30,3,29,159,31,159,30,217,31,2,31,230,31,230,30,212,31,190,31,95,31,147,31,176,31,113,31,202,31,130,31,185,31,86,31,110,31,99,31,235,31,96,31,198,31,191,31,207,31,87,31,87,30,135,31,228,31,254,31,179,31,120,31,211,31,231,31,59,31,12,31,53,31,235,31,140,31,10,31,10,30,84,31,84,30,247,31,247,30,247,29,240,31,240,30,140,31,28,31,190,31,214,31,191,31,191,30,191,29,99,31,197,31,57,31,148,31,148,30,132,31,150,31,198,31,25,31,209,31,209,30,209,29,26,31,117,31,117,30,85,31,5,31,18,31,18,30,68,31,127,31,187,31,187,30,210,31,204,31,54,31,214,31,137,31,137,30,205,31,234,31,211,31,183,31,59,31,252,31,40,31,248,31,96,31,130,31,130,30,158,31,158,30,19,31,21,31,47,31,141,31,147,31,108,31,108,30,206,31,25,31,25,30,162,31,162,30,230,31,107,31,108,31,137,31,137,30,148,31,181,31,181,30,85,31,110,31,110,30,238,31,125,31,179,31,56,31,193,31,118,31,82,31,202,31,111,31,252,31,140,31,140,30,7,31,118,31,136,31,124,31,78,31,95,31,147,31,168,31,26,31,5,31,246,31,12,31,41,31,41,30,174,31,86,31,183,31,102,31,242,31,207,31,220,31,87,31,87,30,244,31,225,31,84,31,159,31,6,31,6,30,6,29,198,31,69,31,32,31,71,31,207,31,122,31,230,31,51,31,225,31,173,31,170,31,1,31,186,31,186,30,202,31,202,31,202,30,135,31,204,31,148,31,158,31,45,31,65,31,196,31,216,31,6,31,113,31,249,31,173,31,98,31,98,30,159,31,73,31,241,31,197,31,121,31,140,31,218,31,185,31,103,31,103,31,48,31,178,31,164,31,164,30,113,31,200,31,116,31,229,31,229,30,229,29,229,28,205,31,106,31,148,31,148,30,80,31,180,31,255,31,212,31,234,31,17,31,17,30,173,31,241,31,204,31,119,31,225,31,225,30,135,31,155,31,155,30,224,31,125,31,249,31,107,31,2,31,129,31,204,31,172,31,64,31,101,31,214,31,214,30,166,31,15,31,225,31,199,31,133,31,141,31,182,31,107,31,136,31,27,31,224,31,98,31,98,30,239,31,68,31,93,31,93,30,93,29,93,28,75,31,139,31,124,31,215,31,215,30,56,31,45,31,45,30,180,31,180,30,28,31,134,31,134,30,52,31,135,31,65,31,65,30,140,31,207,31,207,30,202,31,232,31,92,31,193,31,193,30,194,31,194,30,194,29,194,28,79,31,18,31,225,31,232,31,97,31,78,31,78,30,121,31,165,31,165,30,231,31,80,31,39,31,58,31,34,31,107,31,22,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
