-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_235 is
end project_tb_235;

architecture project_tb_arch_235 of project_tb_235 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 810;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (74,0,215,0,32,0,27,0,143,0,69,0,20,0,182,0,15,0,23,0,253,0,68,0,241,0,72,0,104,0,101,0,200,0,95,0,191,0,0,0,64,0,0,0,176,0,0,0,225,0,11,0,148,0,29,0,42,0,0,0,24,0,90,0,140,0,82,0,145,0,26,0,151,0,45,0,0,0,231,0,134,0,86,0,148,0,131,0,82,0,27,0,139,0,228,0,2,0,239,0,61,0,0,0,17,0,208,0,197,0,0,0,0,0,220,0,99,0,164,0,74,0,104,0,126,0,99,0,15,0,150,0,21,0,248,0,79,0,209,0,222,0,247,0,26,0,98,0,150,0,31,0,198,0,99,0,207,0,251,0,146,0,125,0,12,0,98,0,231,0,31,0,0,0,0,0,73,0,0,0,0,0,18,0,230,0,0,0,252,0,0,0,65,0,237,0,155,0,98,0,79,0,162,0,127,0,242,0,22,0,154,0,114,0,198,0,200,0,0,0,139,0,0,0,174,0,30,0,88,0,213,0,3,0,110,0,62,0,209,0,105,0,0,0,52,0,216,0,219,0,74,0,97,0,86,0,139,0,0,0,93,0,0,0,184,0,191,0,72,0,157,0,0,0,16,0,25,0,156,0,122,0,125,0,245,0,95,0,193,0,0,0,116,0,51,0,68,0,0,0,0,0,46,0,218,0,179,0,0,0,0,0,222,0,223,0,0,0,35,0,103,0,20,0,64,0,41,0,42,0,215,0,90,0,188,0,147,0,225,0,0,0,133,0,4,0,63,0,0,0,59,0,174,0,80,0,0,0,152,0,65,0,0,0,155,0,255,0,246,0,0,0,171,0,59,0,0,0,0,0,0,0,149,0,32,0,215,0,11,0,106,0,18,0,131,0,108,0,211,0,17,0,228,0,0,0,0,0,9,0,4,0,125,0,54,0,24,0,101,0,219,0,84,0,40,0,79,0,177,0,36,0,18,0,0,0,43,0,0,0,0,0,53,0,225,0,182,0,0,0,11,0,173,0,99,0,98,0,121,0,230,0,61,0,0,0,57,0,157,0,212,0,76,0,26,0,158,0,142,0,14,0,112,0,53,0,77,0,65,0,5,0,208,0,0,0,5,0,122,0,102,0,0,0,0,0,144,0,0,0,242,0,160,0,0,0,167,0,170,0,129,0,0,0,191,0,104,0,105,0,154,0,100,0,175,0,28,0,116,0,32,0,55,0,52,0,172,0,213,0,172,0,197,0,195,0,33,0,86,0,0,0,24,0,198,0,53,0,113,0,164,0,152,0,221,0,0,0,11,0,204,0,167,0,223,0,220,0,239,0,144,0,8,0,108,0,70,0,19,0,47,0,220,0,0,0,160,0,224,0,226,0,194,0,187,0,0,0,167,0,156,0,205,0,0,0,131,0,166,0,44,0,98,0,155,0,162,0,117,0,125,0,0,0,43,0,216,0,126,0,13,0,34,0,111,0,13,0,9,0,163,0,0,0,0,0,201,0,175,0,28,0,170,0,244,0,108,0,44,0,149,0,103,0,0,0,0,0,55,0,112,0,0,0,130,0,227,0,133,0,93,0,204,0,119,0,1,0,223,0,202,0,175,0,97,0,126,0,205,0,45,0,34,0,0,0,7,0,0,0,37,0,21,0,183,0,102,0,130,0,197,0,0,0,247,0,170,0,25,0,55,0,174,0,227,0,0,0,0,0,4,0,175,0,0,0,17,0,0,0,82,0,103,0,77,0,164,0,167,0,210,0,124,0,0,0,46,0,72,0,55,0,149,0,25,0,248,0,83,0,0,0,63,0,0,0,0,0,231,0,34,0,103,0,86,0,0,0,150,0,87,0,0,0,184,0,0,0,0,0,161,0,72,0,99,0,174,0,84,0,39,0,0,0,175,0,24,0,37,0,198,0,195,0,112,0,41,0,181,0,253,0,47,0,237,0,0,0,167,0,0,0,221,0,133,0,161,0,120,0,18,0,141,0,246,0,14,0,230,0,54,0,216,0,0,0,29,0,88,0,152,0,143,0,22,0,0,0,77,0,162,0,0,0,202,0,185,0,64,0,118,0,242,0,184,0,55,0,6,0,0,0,212,0,84,0,221,0,40,0,228,0,0,0,32,0,189,0,52,0,227,0,249,0,191,0,49,0,160,0,35,0,208,0,0,0,24,0,118,0,0,0,163,0,129,0,239,0,23,0,186,0,189,0,114,0,216,0,182,0,0,0,0,0,192,0,141,0,204,0,51,0,186,0,43,0,211,0,79,0,0,0,192,0,0,0,141,0,0,0,136,0,0,0,0,0,26,0,97,0,59,0,131,0,0,0,63,0,2,0,121,0,47,0,0,0,14,0,221,0,52,0,239,0,97,0,86,0,47,0,153,0,244,0,107,0,0,0,117,0,192,0,171,0,77,0,0,0,51,0,0,0,0,0,114,0,49,0,57,0,53,0,243,0,0,0,160,0,35,0,30,0,225,0,131,0,191,0,223,0,198,0,116,0,62,0,228,0,0,0,235,0,98,0,174,0,192,0,0,0,15,0,233,0,0,0,0,0,136,0,246,0,23,0,24,0,52,0,10,0,59,0,15,0,0,0,100,0,254,0,71,0,64,0,0,0,186,0,6,0,203,0,0,0,0,0,0,0,22,0,0,0,199,0,0,0,94,0,31,0,34,0,224,0,195,0,239,0,35,0,155,0,106,0,122,0,0,0,199,0,230,0,148,0,19,0,243,0,176,0,189,0,20,0,0,0,94,0,20,0,231,0,189,0,231,0,156,0,110,0,148,0,0,0,0,0,208,0,117,0,26,0,0,0,228,0,165,0,0,0,79,0,0,0,72,0,137,0,0,0,6,0,0,0,130,0,207,0,131,0,0,0,107,0,0,0,57,0,70,0,251,0,0,0,121,0,108,0,120,0,2,0,0,0,117,0,241,0,154,0,47,0,122,0,47,0,198,0,0,0,25,0,0,0,157,0,213,0,0,0,88,0,175,0,30,0,154,0,198,0,172,0,57,0,231,0,43,0,187,0,12,0,0,0,128,0,0,0,126,0,0,0,56,0,216,0,239,0,177,0,50,0,0,0,0,0,158,0,248,0,154,0,180,0,42,0,10,0,0,0,246,0,86,0,0,0,2,0,21,0,108,0,224,0,65,0,105,0,36,0,180,0,146,0,37,0,44,0,165,0,0,0,48,0,67,0,183,0,209,0,0,0,153,0,60,0,140,0,142,0,30,0,96,0,152,0,0,0,33,0,67,0,95,0,89,0,157,0,58,0,114,0,19,0,2,0,0,0,38,0,234,0,0,0,159,0,0,0,109,0,218,0,0,0,162,0,0,0,45,0,19,0,229,0,233,0,127,0,58,0,0,0,95,0,0,0,251,0,45,0,94,0,0,0,0,0,169,0,235,0,183,0,97,0,94,0,62,0,197,0,0,0,23,0,153,0,0,0,42,0,177,0,150,0,52,0,16,0,44,0,18,0,138,0,57,0,181,0,97,0,47,0,104,0,169,0,0,0,14,0,45,0,169,0,32,0,216,0,14,0,150,0,59,0,237,0,18,0,242,0,74,0,28,0,169,0,103,0,215,0,78,0,180,0,0,0,62,0,95,0,48,0,241,0,215,0,114,0,36,0);
signal scenario_full  : scenario_type := (74,31,215,31,32,31,27,31,143,31,69,31,20,31,182,31,15,31,23,31,253,31,68,31,241,31,72,31,104,31,101,31,200,31,95,31,191,31,191,30,64,31,64,30,176,31,176,30,225,31,11,31,148,31,29,31,42,31,42,30,24,31,90,31,140,31,82,31,145,31,26,31,151,31,45,31,45,30,231,31,134,31,86,31,148,31,131,31,82,31,27,31,139,31,228,31,2,31,239,31,61,31,61,30,17,31,208,31,197,31,197,30,197,29,220,31,99,31,164,31,74,31,104,31,126,31,99,31,15,31,150,31,21,31,248,31,79,31,209,31,222,31,247,31,26,31,98,31,150,31,31,31,198,31,99,31,207,31,251,31,146,31,125,31,12,31,98,31,231,31,31,31,31,30,31,29,73,31,73,30,73,29,18,31,230,31,230,30,252,31,252,30,65,31,237,31,155,31,98,31,79,31,162,31,127,31,242,31,22,31,154,31,114,31,198,31,200,31,200,30,139,31,139,30,174,31,30,31,88,31,213,31,3,31,110,31,62,31,209,31,105,31,105,30,52,31,216,31,219,31,74,31,97,31,86,31,139,31,139,30,93,31,93,30,184,31,191,31,72,31,157,31,157,30,16,31,25,31,156,31,122,31,125,31,245,31,95,31,193,31,193,30,116,31,51,31,68,31,68,30,68,29,46,31,218,31,179,31,179,30,179,29,222,31,223,31,223,30,35,31,103,31,20,31,64,31,41,31,42,31,215,31,90,31,188,31,147,31,225,31,225,30,133,31,4,31,63,31,63,30,59,31,174,31,80,31,80,30,152,31,65,31,65,30,155,31,255,31,246,31,246,30,171,31,59,31,59,30,59,29,59,28,149,31,32,31,215,31,11,31,106,31,18,31,131,31,108,31,211,31,17,31,228,31,228,30,228,29,9,31,4,31,125,31,54,31,24,31,101,31,219,31,84,31,40,31,79,31,177,31,36,31,18,31,18,30,43,31,43,30,43,29,53,31,225,31,182,31,182,30,11,31,173,31,99,31,98,31,121,31,230,31,61,31,61,30,57,31,157,31,212,31,76,31,26,31,158,31,142,31,14,31,112,31,53,31,77,31,65,31,5,31,208,31,208,30,5,31,122,31,102,31,102,30,102,29,144,31,144,30,242,31,160,31,160,30,167,31,170,31,129,31,129,30,191,31,104,31,105,31,154,31,100,31,175,31,28,31,116,31,32,31,55,31,52,31,172,31,213,31,172,31,197,31,195,31,33,31,86,31,86,30,24,31,198,31,53,31,113,31,164,31,152,31,221,31,221,30,11,31,204,31,167,31,223,31,220,31,239,31,144,31,8,31,108,31,70,31,19,31,47,31,220,31,220,30,160,31,224,31,226,31,194,31,187,31,187,30,167,31,156,31,205,31,205,30,131,31,166,31,44,31,98,31,155,31,162,31,117,31,125,31,125,30,43,31,216,31,126,31,13,31,34,31,111,31,13,31,9,31,163,31,163,30,163,29,201,31,175,31,28,31,170,31,244,31,108,31,44,31,149,31,103,31,103,30,103,29,55,31,112,31,112,30,130,31,227,31,133,31,93,31,204,31,119,31,1,31,223,31,202,31,175,31,97,31,126,31,205,31,45,31,34,31,34,30,7,31,7,30,37,31,21,31,183,31,102,31,130,31,197,31,197,30,247,31,170,31,25,31,55,31,174,31,227,31,227,30,227,29,4,31,175,31,175,30,17,31,17,30,82,31,103,31,77,31,164,31,167,31,210,31,124,31,124,30,46,31,72,31,55,31,149,31,25,31,248,31,83,31,83,30,63,31,63,30,63,29,231,31,34,31,103,31,86,31,86,30,150,31,87,31,87,30,184,31,184,30,184,29,161,31,72,31,99,31,174,31,84,31,39,31,39,30,175,31,24,31,37,31,198,31,195,31,112,31,41,31,181,31,253,31,47,31,237,31,237,30,167,31,167,30,221,31,133,31,161,31,120,31,18,31,141,31,246,31,14,31,230,31,54,31,216,31,216,30,29,31,88,31,152,31,143,31,22,31,22,30,77,31,162,31,162,30,202,31,185,31,64,31,118,31,242,31,184,31,55,31,6,31,6,30,212,31,84,31,221,31,40,31,228,31,228,30,32,31,189,31,52,31,227,31,249,31,191,31,49,31,160,31,35,31,208,31,208,30,24,31,118,31,118,30,163,31,129,31,239,31,23,31,186,31,189,31,114,31,216,31,182,31,182,30,182,29,192,31,141,31,204,31,51,31,186,31,43,31,211,31,79,31,79,30,192,31,192,30,141,31,141,30,136,31,136,30,136,29,26,31,97,31,59,31,131,31,131,30,63,31,2,31,121,31,47,31,47,30,14,31,221,31,52,31,239,31,97,31,86,31,47,31,153,31,244,31,107,31,107,30,117,31,192,31,171,31,77,31,77,30,51,31,51,30,51,29,114,31,49,31,57,31,53,31,243,31,243,30,160,31,35,31,30,31,225,31,131,31,191,31,223,31,198,31,116,31,62,31,228,31,228,30,235,31,98,31,174,31,192,31,192,30,15,31,233,31,233,30,233,29,136,31,246,31,23,31,24,31,52,31,10,31,59,31,15,31,15,30,100,31,254,31,71,31,64,31,64,30,186,31,6,31,203,31,203,30,203,29,203,28,22,31,22,30,199,31,199,30,94,31,31,31,34,31,224,31,195,31,239,31,35,31,155,31,106,31,122,31,122,30,199,31,230,31,148,31,19,31,243,31,176,31,189,31,20,31,20,30,94,31,20,31,231,31,189,31,231,31,156,31,110,31,148,31,148,30,148,29,208,31,117,31,26,31,26,30,228,31,165,31,165,30,79,31,79,30,72,31,137,31,137,30,6,31,6,30,130,31,207,31,131,31,131,30,107,31,107,30,57,31,70,31,251,31,251,30,121,31,108,31,120,31,2,31,2,30,117,31,241,31,154,31,47,31,122,31,47,31,198,31,198,30,25,31,25,30,157,31,213,31,213,30,88,31,175,31,30,31,154,31,198,31,172,31,57,31,231,31,43,31,187,31,12,31,12,30,128,31,128,30,126,31,126,30,56,31,216,31,239,31,177,31,50,31,50,30,50,29,158,31,248,31,154,31,180,31,42,31,10,31,10,30,246,31,86,31,86,30,2,31,21,31,108,31,224,31,65,31,105,31,36,31,180,31,146,31,37,31,44,31,165,31,165,30,48,31,67,31,183,31,209,31,209,30,153,31,60,31,140,31,142,31,30,31,96,31,152,31,152,30,33,31,67,31,95,31,89,31,157,31,58,31,114,31,19,31,2,31,2,30,38,31,234,31,234,30,159,31,159,30,109,31,218,31,218,30,162,31,162,30,45,31,19,31,229,31,233,31,127,31,58,31,58,30,95,31,95,30,251,31,45,31,94,31,94,30,94,29,169,31,235,31,183,31,97,31,94,31,62,31,197,31,197,30,23,31,153,31,153,30,42,31,177,31,150,31,52,31,16,31,44,31,18,31,138,31,57,31,181,31,97,31,47,31,104,31,169,31,169,30,14,31,45,31,169,31,32,31,216,31,14,31,150,31,59,31,237,31,18,31,242,31,74,31,28,31,169,31,103,31,215,31,78,31,180,31,180,30,62,31,95,31,48,31,241,31,215,31,114,31,36,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
