-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 221;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (110,0,189,0,39,0,116,0,27,0,230,0,203,0,3,0,208,0,224,0,250,0,3,0,55,0,218,0,189,0,119,0,0,0,108,0,53,0,142,0,0,0,161,0,143,0,192,0,0,0,128,0,70,0,51,0,0,0,168,0,0,0,230,0,0,0,97,0,231,0,222,0,253,0,184,0,0,0,0,0,249,0,142,0,247,0,126,0,97,0,155,0,0,0,66,0,154,0,116,0,5,0,124,0,71,0,141,0,0,0,93,0,0,0,0,0,13,0,0,0,13,0,245,0,179,0,210,0,0,0,14,0,0,0,0,0,29,0,219,0,24,0,21,0,201,0,177,0,173,0,185,0,221,0,146,0,254,0,14,0,154,0,127,0,45,0,255,0,0,0,85,0,135,0,19,0,202,0,0,0,253,0,198,0,11,0,28,0,249,0,216,0,0,0,0,0,250,0,209,0,235,0,132,0,0,0,0,0,0,0,185,0,110,0,66,0,27,0,168,0,0,0,85,0,22,0,238,0,162,0,239,0,223,0,67,0,0,0,231,0,106,0,185,0,0,0,252,0,3,0,95,0,0,0,112,0,0,0,0,0,121,0,141,0,160,0,0,0,0,0,30,0,106,0,130,0,41,0,86,0,0,0,153,0,212,0,0,0,182,0,78,0,133,0,109,0,0,0,161,0,162,0,161,0,112,0,0,0,107,0,129,0,232,0,1,0,78,0,154,0,174,0,101,0,240,0,0,0,102,0,0,0,73,0,69,0,122,0,97,0,205,0,180,0,82,0,241,0,0,0,64,0,204,0,167,0,0,0,107,0,53,0,0,0,3,0,133,0,253,0,182,0,7,0,0,0,109,0,143,0,235,0,0,0,0,0,0,0,0,0,37,0,152,0,0,0,0,0,251,0,85,0,0,0,163,0,0,0,177,0,111,0,206,0,0,0,111,0,209,0,5,0,0,0,138,0,151,0,51,0,118,0,0,0,0,0,233,0,73,0,156,0);
signal scenario_full  : scenario_type := (110,31,189,31,39,31,116,31,27,31,230,31,203,31,3,31,208,31,224,31,250,31,3,31,55,31,218,31,189,31,119,31,119,30,108,31,53,31,142,31,142,30,161,31,143,31,192,31,192,30,128,31,70,31,51,31,51,30,168,31,168,30,230,31,230,30,97,31,231,31,222,31,253,31,184,31,184,30,184,29,249,31,142,31,247,31,126,31,97,31,155,31,155,30,66,31,154,31,116,31,5,31,124,31,71,31,141,31,141,30,93,31,93,30,93,29,13,31,13,30,13,31,245,31,179,31,210,31,210,30,14,31,14,30,14,29,29,31,219,31,24,31,21,31,201,31,177,31,173,31,185,31,221,31,146,31,254,31,14,31,154,31,127,31,45,31,255,31,255,30,85,31,135,31,19,31,202,31,202,30,253,31,198,31,11,31,28,31,249,31,216,31,216,30,216,29,250,31,209,31,235,31,132,31,132,30,132,29,132,28,185,31,110,31,66,31,27,31,168,31,168,30,85,31,22,31,238,31,162,31,239,31,223,31,67,31,67,30,231,31,106,31,185,31,185,30,252,31,3,31,95,31,95,30,112,31,112,30,112,29,121,31,141,31,160,31,160,30,160,29,30,31,106,31,130,31,41,31,86,31,86,30,153,31,212,31,212,30,182,31,78,31,133,31,109,31,109,30,161,31,162,31,161,31,112,31,112,30,107,31,129,31,232,31,1,31,78,31,154,31,174,31,101,31,240,31,240,30,102,31,102,30,73,31,69,31,122,31,97,31,205,31,180,31,82,31,241,31,241,30,64,31,204,31,167,31,167,30,107,31,53,31,53,30,3,31,133,31,253,31,182,31,7,31,7,30,109,31,143,31,235,31,235,30,235,29,235,28,235,27,37,31,152,31,152,30,152,29,251,31,85,31,85,30,163,31,163,30,177,31,111,31,206,31,206,30,111,31,209,31,5,31,5,30,138,31,151,31,51,31,118,31,118,30,118,29,233,31,73,31,156,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
