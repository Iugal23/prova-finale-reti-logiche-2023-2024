-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 507;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,31,0,64,0,57,0,0,0,220,0,228,0,111,0,0,0,0,0,0,0,111,0,0,0,248,0,251,0,11,0,0,0,80,0,201,0,82,0,81,0,113,0,1,0,0,0,78,0,164,0,192,0,249,0,0,0,180,0,70,0,243,0,0,0,129,0,0,0,249,0,0,0,32,0,0,0,144,0,228,0,29,0,0,0,118,0,229,0,122,0,101,0,99,0,239,0,179,0,223,0,7,0,96,0,0,0,213,0,80,0,61,0,0,0,0,0,138,0,0,0,7,0,38,0,31,0,0,0,33,0,0,0,44,0,233,0,0,0,82,0,6,0,197,0,97,0,251,0,0,0,86,0,89,0,55,0,27,0,171,0,67,0,0,0,13,0,16,0,11,0,199,0,0,0,29,0,78,0,200,0,173,0,184,0,59,0,78,0,236,0,192,0,0,0,177,0,106,0,240,0,191,0,53,0,185,0,43,0,161,0,4,0,85,0,248,0,178,0,0,0,50,0,210,0,190,0,34,0,0,0,163,0,187,0,230,0,163,0,0,0,39,0,50,0,125,0,0,0,90,0,0,0,135,0,58,0,125,0,0,0,156,0,75,0,0,0,202,0,2,0,60,0,201,0,0,0,230,0,31,0,126,0,0,0,62,0,83,0,150,0,0,0,0,0,250,0,13,0,127,0,233,0,212,0,174,0,141,0,0,0,3,0,107,0,11,0,142,0,161,0,0,0,109,0,176,0,254,0,4,0,161,0,48,0,45,0,169,0,98,0,38,0,0,0,156,0,26,0,52,0,53,0,27,0,200,0,200,0,142,0,61,0,75,0,28,0,75,0,40,0,21,0,88,0,0,0,48,0,0,0,0,0,0,0,14,0,140,0,223,0,191,0,0,0,30,0,64,0,5,0,130,0,0,0,216,0,138,0,67,0,152,0,47,0,242,0,72,0,126,0,246,0,133,0,194,0,161,0,106,0,224,0,251,0,0,0,210,0,40,0,176,0,172,0,116,0,192,0,223,0,184,0,210,0,146,0,0,0,237,0,88,0,154,0,0,0,213,0,72,0,238,0,107,0,0,0,175,0,100,0,145,0,184,0,194,0,128,0,245,0,189,0,210,0,25,0,146,0,137,0,140,0,89,0,6,0,199,0,252,0,30,0,254,0,163,0,0,0,241,0,0,0,213,0,202,0,150,0,0,0,84,0,112,0,141,0,201,0,222,0,69,0,63,0,238,0,25,0,128,0,242,0,174,0,206,0,167,0,246,0,86,0,247,0,237,0,166,0,179,0,162,0,0,0,207,0,215,0,0,0,162,0,141,0,157,0,126,0,0,0,95,0,0,0,213,0,4,0,24,0,227,0,141,0,188,0,112,0,158,0,60,0,19,0,220,0,0,0,0,0,160,0,144,0,150,0,139,0,98,0,177,0,0,0,254,0,187,0,228,0,47,0,98,0,171,0,193,0,0,0,156,0,87,0,113,0,167,0,216,0,239,0,0,0,102,0,0,0,210,0,64,0,0,0,0,0,200,0,103,0,67,0,0,0,0,0,16,0,0,0,13,0,153,0,150,0,15,0,59,0,205,0,249,0,152,0,3,0,0,0,23,0,50,0,245,0,0,0,227,0,255,0,0,0,144,0,126,0,110,0,105,0,123,0,0,0,168,0,142,0,122,0,71,0,27,0,28,0,228,0,219,0,6,0,62,0,22,0,224,0,90,0,176,0,166,0,90,0,140,0,175,0,106,0,139,0,25,0,71,0,96,0,0,0,166,0,131,0,151,0,159,0,75,0,231,0,195,0,176,0,8,0,177,0,0,0,72,0,191,0,58,0,43,0,118,0,72,0,0,0,0,0,25,0,8,0,206,0,42,0,76,0,99,0,88,0,231,0,170,0,0,0,71,0,20,0,251,0,66,0,158,0,94,0,81,0,30,0,254,0,132,0,132,0,193,0,0,0,98,0,0,0,178,0,29,0,126,0,61,0,134,0,143,0,108,0,4,0,108,0,154,0,78,0,44,0,0,0,0,0,168,0,11,0,141,0,20,0,88,0,48,0,181,0,12,0,0,0,234,0,123,0,190,0,0,0,251,0,193,0,34,0,177,0,66,0,9,0,150,0,130,0,128,0,250,0,25,0,0,0,86,0,0,0,102,0,0,0,120,0,250,0,36,0,97,0,214,0,0,0,100,0,0,0,0,0,0,0,100,0,210,0,113,0,0,0,193,0,39,0,139,0,0,0,58,0,0,0,9,0,235,0,0,0,0,0,177,0,0,0,224,0);
signal scenario_full  : scenario_type := (0,0,31,31,64,31,57,31,57,30,220,31,228,31,111,31,111,30,111,29,111,28,111,31,111,30,248,31,251,31,11,31,11,30,80,31,201,31,82,31,81,31,113,31,1,31,1,30,78,31,164,31,192,31,249,31,249,30,180,31,70,31,243,31,243,30,129,31,129,30,249,31,249,30,32,31,32,30,144,31,228,31,29,31,29,30,118,31,229,31,122,31,101,31,99,31,239,31,179,31,223,31,7,31,96,31,96,30,213,31,80,31,61,31,61,30,61,29,138,31,138,30,7,31,38,31,31,31,31,30,33,31,33,30,44,31,233,31,233,30,82,31,6,31,197,31,97,31,251,31,251,30,86,31,89,31,55,31,27,31,171,31,67,31,67,30,13,31,16,31,11,31,199,31,199,30,29,31,78,31,200,31,173,31,184,31,59,31,78,31,236,31,192,31,192,30,177,31,106,31,240,31,191,31,53,31,185,31,43,31,161,31,4,31,85,31,248,31,178,31,178,30,50,31,210,31,190,31,34,31,34,30,163,31,187,31,230,31,163,31,163,30,39,31,50,31,125,31,125,30,90,31,90,30,135,31,58,31,125,31,125,30,156,31,75,31,75,30,202,31,2,31,60,31,201,31,201,30,230,31,31,31,126,31,126,30,62,31,83,31,150,31,150,30,150,29,250,31,13,31,127,31,233,31,212,31,174,31,141,31,141,30,3,31,107,31,11,31,142,31,161,31,161,30,109,31,176,31,254,31,4,31,161,31,48,31,45,31,169,31,98,31,38,31,38,30,156,31,26,31,52,31,53,31,27,31,200,31,200,31,142,31,61,31,75,31,28,31,75,31,40,31,21,31,88,31,88,30,48,31,48,30,48,29,48,28,14,31,140,31,223,31,191,31,191,30,30,31,64,31,5,31,130,31,130,30,216,31,138,31,67,31,152,31,47,31,242,31,72,31,126,31,246,31,133,31,194,31,161,31,106,31,224,31,251,31,251,30,210,31,40,31,176,31,172,31,116,31,192,31,223,31,184,31,210,31,146,31,146,30,237,31,88,31,154,31,154,30,213,31,72,31,238,31,107,31,107,30,175,31,100,31,145,31,184,31,194,31,128,31,245,31,189,31,210,31,25,31,146,31,137,31,140,31,89,31,6,31,199,31,252,31,30,31,254,31,163,31,163,30,241,31,241,30,213,31,202,31,150,31,150,30,84,31,112,31,141,31,201,31,222,31,69,31,63,31,238,31,25,31,128,31,242,31,174,31,206,31,167,31,246,31,86,31,247,31,237,31,166,31,179,31,162,31,162,30,207,31,215,31,215,30,162,31,141,31,157,31,126,31,126,30,95,31,95,30,213,31,4,31,24,31,227,31,141,31,188,31,112,31,158,31,60,31,19,31,220,31,220,30,220,29,160,31,144,31,150,31,139,31,98,31,177,31,177,30,254,31,187,31,228,31,47,31,98,31,171,31,193,31,193,30,156,31,87,31,113,31,167,31,216,31,239,31,239,30,102,31,102,30,210,31,64,31,64,30,64,29,200,31,103,31,67,31,67,30,67,29,16,31,16,30,13,31,153,31,150,31,15,31,59,31,205,31,249,31,152,31,3,31,3,30,23,31,50,31,245,31,245,30,227,31,255,31,255,30,144,31,126,31,110,31,105,31,123,31,123,30,168,31,142,31,122,31,71,31,27,31,28,31,228,31,219,31,6,31,62,31,22,31,224,31,90,31,176,31,166,31,90,31,140,31,175,31,106,31,139,31,25,31,71,31,96,31,96,30,166,31,131,31,151,31,159,31,75,31,231,31,195,31,176,31,8,31,177,31,177,30,72,31,191,31,58,31,43,31,118,31,72,31,72,30,72,29,25,31,8,31,206,31,42,31,76,31,99,31,88,31,231,31,170,31,170,30,71,31,20,31,251,31,66,31,158,31,94,31,81,31,30,31,254,31,132,31,132,31,193,31,193,30,98,31,98,30,178,31,29,31,126,31,61,31,134,31,143,31,108,31,4,31,108,31,154,31,78,31,44,31,44,30,44,29,168,31,11,31,141,31,20,31,88,31,48,31,181,31,12,31,12,30,234,31,123,31,190,31,190,30,251,31,193,31,34,31,177,31,66,31,9,31,150,31,130,31,128,31,250,31,25,31,25,30,86,31,86,30,102,31,102,30,120,31,250,31,36,31,97,31,214,31,214,30,100,31,100,30,100,29,100,28,100,31,210,31,113,31,113,30,193,31,39,31,139,31,139,30,58,31,58,30,9,31,235,31,235,30,235,29,177,31,177,30,224,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
