-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 684;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (137,0,0,0,228,0,96,0,195,0,118,0,0,0,0,0,171,0,235,0,211,0,176,0,169,0,66,0,149,0,165,0,194,0,187,0,113,0,36,0,170,0,0,0,212,0,218,0,15,0,188,0,241,0,241,0,173,0,15,0,20,0,165,0,19,0,46,0,0,0,223,0,12,0,178,0,103,0,0,0,214,0,16,0,0,0,88,0,138,0,0,0,86,0,79,0,39,0,13,0,82,0,231,0,191,0,145,0,134,0,12,0,150,0,172,0,249,0,182,0,0,0,244,0,0,0,245,0,248,0,118,0,11,0,242,0,222,0,0,0,0,0,76,0,251,0,237,0,253,0,0,0,60,0,238,0,0,0,244,0,199,0,0,0,138,0,78,0,243,0,29,0,252,0,88,0,222,0,136,0,81,0,253,0,220,0,226,0,169,0,95,0,217,0,0,0,37,0,60,0,159,0,0,0,0,0,94,0,98,0,123,0,0,0,32,0,113,0,0,0,140,0,143,0,217,0,4,0,121,0,251,0,128,0,242,0,25,0,132,0,254,0,94,0,143,0,9,0,0,0,252,0,178,0,48,0,119,0,0,0,50,0,160,0,183,0,137,0,250,0,79,0,165,0,36,0,61,0,0,0,159,0,150,0,0,0,0,0,0,0,0,0,161,0,113,0,149,0,109,0,90,0,20,0,0,0,98,0,137,0,8,0,120,0,161,0,0,0,11,0,59,0,58,0,0,0,0,0,133,0,168,0,250,0,96,0,49,0,219,0,126,0,0,0,2,0,92,0,242,0,162,0,0,0,0,0,87,0,107,0,159,0,0,0,151,0,0,0,219,0,0,0,210,0,19,0,91,0,244,0,76,0,38,0,0,0,236,0,0,0,89,0,193,0,69,0,210,0,0,0,154,0,201,0,150,0,189,0,0,0,0,0,181,0,134,0,203,0,81,0,5,0,0,0,231,0,251,0,0,0,0,0,0,0,3,0,177,0,0,0,37,0,0,0,199,0,132,0,34,0,8,0,165,0,0,0,81,0,126,0,95,0,91,0,0,0,127,0,106,0,111,0,158,0,36,0,0,0,216,0,0,0,168,0,123,0,166,0,0,0,136,0,157,0,1,0,102,0,53,0,207,0,89,0,177,0,198,0,17,0,0,0,0,0,0,0,0,0,164,0,228,0,0,0,36,0,118,0,237,0,77,0,202,0,0,0,119,0,0,0,78,0,110,0,206,0,0,0,103,0,123,0,61,0,0,0,0,0,114,0,186,0,0,0,114,0,243,0,207,0,61,0,130,0,236,0,110,0,0,0,154,0,80,0,127,0,184,0,28,0,85,0,83,0,108,0,226,0,227,0,243,0,0,0,119,0,195,0,148,0,143,0,148,0,198,0,254,0,215,0,161,0,0,0,90,0,123,0,0,0,34,0,240,0,202,0,58,0,0,0,0,0,63,0,0,0,126,0,0,0,0,0,167,0,32,0,0,0,0,0,242,0,73,0,225,0,105,0,50,0,113,0,144,0,184,0,78,0,61,0,117,0,171,0,33,0,84,0,177,0,19,0,229,0,154,0,62,0,216,0,0,0,64,0,0,0,0,0,0,0,196,0,109,0,234,0,0,0,15,0,134,0,28,0,172,0,55,0,144,0,6,0,46,0,245,0,37,0,50,0,166,0,202,0,163,0,98,0,128,0,0,0,91,0,241,0,0,0,166,0,62,0,80,0,49,0,107,0,38,0,27,0,156,0,0,0,0,0,252,0,99,0,245,0,81,0,16,0,94,0,28,0,18,0,224,0,0,0,175,0,56,0,219,0,230,0,0,0,0,0,172,0,55,0,0,0,0,0,189,0,71,0,207,0,83,0,224,0,174,0,172,0,5,0,0,0,0,0,122,0,106,0,111,0,213,0,27,0,137,0,134,0,0,0,151,0,34,0,0,0,124,0,196,0,208,0,204,0,224,0,0,0,208,0,90,0,0,0,143,0,203,0,153,0,233,0,117,0,0,0,140,0,71,0,73,0,132,0,77,0,196,0,114,0,62,0,16,0,232,0,86,0,222,0,212,0,177,0,0,0,2,0,57,0,0,0,233,0,53,0,169,0,0,0,150,0,34,0,234,0,249,0,82,0,244,0,154,0,101,0,0,0,250,0,196,0,34,0,237,0,155,0,71,0,0,0,39,0,84,0,136,0,0,0,224,0,157,0,200,0,189,0,0,0,175,0,215,0,0,0,103,0,170,0,0,0,220,0,44,0,41,0,244,0,50,0,40,0,127,0,215,0,161,0,141,0,150,0,0,0,203,0,139,0,148,0,101,0,24,0,226,0,242,0,241,0,81,0,0,0,72,0,121,0,242,0,110,0,147,0,138,0,227,0,0,0,229,0,98,0,172,0,59,0,0,0,112,0,3,0,7,0,0,0,171,0,109,0,218,0,241,0,135,0,106,0,173,0,0,0,0,0,0,0,0,0,196,0,213,0,0,0,130,0,170,0,12,0,251,0,145,0,239,0,208,0,0,0,189,0,228,0,181,0,74,0,0,0,123,0,169,0,169,0,164,0,172,0,0,0,231,0,0,0,154,0,124,0,0,0,1,0,43,0,210,0,170,0,71,0,152,0,0,0,201,0,68,0,153,0,13,0,31,0,50,0,57,0,168,0,137,0,74,0,35,0,19,0,0,0,75,0,72,0,219,0,0,0,199,0,252,0,124,0,57,0,153,0,68,0,229,0,60,0,193,0,0,0,0,0,55,0,49,0,92,0,94,0,75,0,207,0,71,0,41,0,126,0,66,0,0,0,208,0,154,0,137,0,0,0,160,0,44,0,230,0,83,0,239,0,0,0,0,0,0,0,181,0,78,0,224,0,57,0,76,0,0,0,212,0,233,0,0,0,209,0,217,0,98,0,0,0,218,0,200,0,49,0,48,0,222,0,149,0,164,0,249,0,89,0,190,0,155,0,248,0,103,0,91,0,189,0,232,0,194,0,117,0,250,0,0,0,133,0,13,0,203,0,25,0,152,0,9,0,143,0,42,0,158,0,212,0,0,0,115,0,119,0,212,0,32,0,0,0,159,0,104,0);
signal scenario_full  : scenario_type := (137,31,137,30,228,31,96,31,195,31,118,31,118,30,118,29,171,31,235,31,211,31,176,31,169,31,66,31,149,31,165,31,194,31,187,31,113,31,36,31,170,31,170,30,212,31,218,31,15,31,188,31,241,31,241,31,173,31,15,31,20,31,165,31,19,31,46,31,46,30,223,31,12,31,178,31,103,31,103,30,214,31,16,31,16,30,88,31,138,31,138,30,86,31,79,31,39,31,13,31,82,31,231,31,191,31,145,31,134,31,12,31,150,31,172,31,249,31,182,31,182,30,244,31,244,30,245,31,248,31,118,31,11,31,242,31,222,31,222,30,222,29,76,31,251,31,237,31,253,31,253,30,60,31,238,31,238,30,244,31,199,31,199,30,138,31,78,31,243,31,29,31,252,31,88,31,222,31,136,31,81,31,253,31,220,31,226,31,169,31,95,31,217,31,217,30,37,31,60,31,159,31,159,30,159,29,94,31,98,31,123,31,123,30,32,31,113,31,113,30,140,31,143,31,217,31,4,31,121,31,251,31,128,31,242,31,25,31,132,31,254,31,94,31,143,31,9,31,9,30,252,31,178,31,48,31,119,31,119,30,50,31,160,31,183,31,137,31,250,31,79,31,165,31,36,31,61,31,61,30,159,31,150,31,150,30,150,29,150,28,150,27,161,31,113,31,149,31,109,31,90,31,20,31,20,30,98,31,137,31,8,31,120,31,161,31,161,30,11,31,59,31,58,31,58,30,58,29,133,31,168,31,250,31,96,31,49,31,219,31,126,31,126,30,2,31,92,31,242,31,162,31,162,30,162,29,87,31,107,31,159,31,159,30,151,31,151,30,219,31,219,30,210,31,19,31,91,31,244,31,76,31,38,31,38,30,236,31,236,30,89,31,193,31,69,31,210,31,210,30,154,31,201,31,150,31,189,31,189,30,189,29,181,31,134,31,203,31,81,31,5,31,5,30,231,31,251,31,251,30,251,29,251,28,3,31,177,31,177,30,37,31,37,30,199,31,132,31,34,31,8,31,165,31,165,30,81,31,126,31,95,31,91,31,91,30,127,31,106,31,111,31,158,31,36,31,36,30,216,31,216,30,168,31,123,31,166,31,166,30,136,31,157,31,1,31,102,31,53,31,207,31,89,31,177,31,198,31,17,31,17,30,17,29,17,28,17,27,164,31,228,31,228,30,36,31,118,31,237,31,77,31,202,31,202,30,119,31,119,30,78,31,110,31,206,31,206,30,103,31,123,31,61,31,61,30,61,29,114,31,186,31,186,30,114,31,243,31,207,31,61,31,130,31,236,31,110,31,110,30,154,31,80,31,127,31,184,31,28,31,85,31,83,31,108,31,226,31,227,31,243,31,243,30,119,31,195,31,148,31,143,31,148,31,198,31,254,31,215,31,161,31,161,30,90,31,123,31,123,30,34,31,240,31,202,31,58,31,58,30,58,29,63,31,63,30,126,31,126,30,126,29,167,31,32,31,32,30,32,29,242,31,73,31,225,31,105,31,50,31,113,31,144,31,184,31,78,31,61,31,117,31,171,31,33,31,84,31,177,31,19,31,229,31,154,31,62,31,216,31,216,30,64,31,64,30,64,29,64,28,196,31,109,31,234,31,234,30,15,31,134,31,28,31,172,31,55,31,144,31,6,31,46,31,245,31,37,31,50,31,166,31,202,31,163,31,98,31,128,31,128,30,91,31,241,31,241,30,166,31,62,31,80,31,49,31,107,31,38,31,27,31,156,31,156,30,156,29,252,31,99,31,245,31,81,31,16,31,94,31,28,31,18,31,224,31,224,30,175,31,56,31,219,31,230,31,230,30,230,29,172,31,55,31,55,30,55,29,189,31,71,31,207,31,83,31,224,31,174,31,172,31,5,31,5,30,5,29,122,31,106,31,111,31,213,31,27,31,137,31,134,31,134,30,151,31,34,31,34,30,124,31,196,31,208,31,204,31,224,31,224,30,208,31,90,31,90,30,143,31,203,31,153,31,233,31,117,31,117,30,140,31,71,31,73,31,132,31,77,31,196,31,114,31,62,31,16,31,232,31,86,31,222,31,212,31,177,31,177,30,2,31,57,31,57,30,233,31,53,31,169,31,169,30,150,31,34,31,234,31,249,31,82,31,244,31,154,31,101,31,101,30,250,31,196,31,34,31,237,31,155,31,71,31,71,30,39,31,84,31,136,31,136,30,224,31,157,31,200,31,189,31,189,30,175,31,215,31,215,30,103,31,170,31,170,30,220,31,44,31,41,31,244,31,50,31,40,31,127,31,215,31,161,31,141,31,150,31,150,30,203,31,139,31,148,31,101,31,24,31,226,31,242,31,241,31,81,31,81,30,72,31,121,31,242,31,110,31,147,31,138,31,227,31,227,30,229,31,98,31,172,31,59,31,59,30,112,31,3,31,7,31,7,30,171,31,109,31,218,31,241,31,135,31,106,31,173,31,173,30,173,29,173,28,173,27,196,31,213,31,213,30,130,31,170,31,12,31,251,31,145,31,239,31,208,31,208,30,189,31,228,31,181,31,74,31,74,30,123,31,169,31,169,31,164,31,172,31,172,30,231,31,231,30,154,31,124,31,124,30,1,31,43,31,210,31,170,31,71,31,152,31,152,30,201,31,68,31,153,31,13,31,31,31,50,31,57,31,168,31,137,31,74,31,35,31,19,31,19,30,75,31,72,31,219,31,219,30,199,31,252,31,124,31,57,31,153,31,68,31,229,31,60,31,193,31,193,30,193,29,55,31,49,31,92,31,94,31,75,31,207,31,71,31,41,31,126,31,66,31,66,30,208,31,154,31,137,31,137,30,160,31,44,31,230,31,83,31,239,31,239,30,239,29,239,28,181,31,78,31,224,31,57,31,76,31,76,30,212,31,233,31,233,30,209,31,217,31,98,31,98,30,218,31,200,31,49,31,48,31,222,31,149,31,164,31,249,31,89,31,190,31,155,31,248,31,103,31,91,31,189,31,232,31,194,31,117,31,250,31,250,30,133,31,13,31,203,31,25,31,152,31,9,31,143,31,42,31,158,31,212,31,212,30,115,31,119,31,212,31,32,31,32,30,159,31,104,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
