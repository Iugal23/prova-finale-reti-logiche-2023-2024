-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_96 is
end project_tb_96;

architecture project_tb_arch_96 of project_tb_96 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 696;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (135,0,167,0,184,0,142,0,0,0,181,0,5,0,76,0,88,0,228,0,0,0,206,0,154,0,245,0,0,0,201,0,45,0,154,0,184,0,182,0,0,0,141,0,117,0,177,0,89,0,189,0,0,0,193,0,121,0,0,0,0,0,0,0,161,0,180,0,0,0,91,0,164,0,178,0,152,0,207,0,0,0,174,0,196,0,0,0,0,0,196,0,180,0,235,0,205,0,82,0,0,0,104,0,145,0,54,0,80,0,128,0,138,0,166,0,167,0,54,0,123,0,240,0,0,0,0,0,13,0,61,0,239,0,130,0,91,0,135,0,205,0,244,0,19,0,202,0,0,0,68,0,254,0,116,0,0,0,0,0,98,0,185,0,181,0,213,0,178,0,186,0,201,0,38,0,208,0,118,0,171,0,0,0,0,0,0,0,42,0,210,0,50,0,91,0,35,0,17,0,235,0,0,0,6,0,69,0,14,0,61,0,0,0,130,0,52,0,0,0,0,0,211,0,37,0,182,0,133,0,138,0,243,0,116,0,0,0,64,0,129,0,45,0,61,0,0,0,221,0,205,0,0,0,156,0,0,0,0,0,24,0,98,0,77,0,242,0,172,0,128,0,0,0,107,0,28,0,69,0,154,0,112,0,0,0,245,0,231,0,129,0,196,0,247,0,0,0,55,0,184,0,220,0,0,0,97,0,74,0,0,0,123,0,136,0,148,0,226,0,147,0,216,0,167,0,85,0,12,0,234,0,0,0,0,0,44,0,245,0,0,0,48,0,50,0,19,0,36,0,22,0,179,0,207,0,190,0,0,0,221,0,28,0,130,0,151,0,76,0,206,0,203,0,2,0,209,0,78,0,138,0,106,0,0,0,112,0,195,0,235,0,0,0,195,0,71,0,114,0,0,0,238,0,30,0,97,0,51,0,191,0,75,0,23,0,35,0,0,0,250,0,157,0,254,0,232,0,231,0,25,0,82,0,236,0,113,0,57,0,0,0,67,0,0,0,172,0,248,0,1,0,156,0,74,0,0,0,252,0,251,0,203,0,0,0,0,0,9,0,34,0,121,0,203,0,162,0,0,0,86,0,1,0,105,0,163,0,157,0,25,0,123,0,48,0,139,0,129,0,0,0,13,0,181,0,179,0,45,0,0,0,181,0,235,0,195,0,150,0,0,0,158,0,0,0,25,0,0,0,217,0,0,0,0,0,54,0,165,0,143,0,0,0,0,0,192,0,241,0,0,0,249,0,103,0,122,0,160,0,100,0,159,0,105,0,84,0,0,0,221,0,213,0,216,0,140,0,237,0,173,0,29,0,87,0,8,0,252,0,105,0,228,0,0,0,222,0,37,0,86,0,35,0,195,0,81,0,53,0,22,0,100,0,156,0,0,0,252,0,71,0,148,0,138,0,18,0,0,0,50,0,0,0,0,0,161,0,27,0,92,0,5,0,49,0,206,0,56,0,65,0,36,0,204,0,61,0,0,0,39,0,189,0,110,0,253,0,0,0,133,0,137,0,0,0,28,0,0,0,20,0,0,0,92,0,44,0,103,0,182,0,93,0,251,0,69,0,160,0,234,0,0,0,139,0,126,0,105,0,224,0,199,0,0,0,88,0,118,0,93,0,111,0,0,0,81,0,176,0,251,0,116,0,99,0,0,0,15,0,0,0,114,0,158,0,0,0,0,0,0,0,130,0,34,0,173,0,0,0,56,0,210,0,124,0,236,0,135,0,153,0,37,0,247,0,33,0,178,0,0,0,190,0,119,0,0,0,243,0,161,0,140,0,20,0,17,0,65,0,146,0,192,0,22,0,202,0,175,0,158,0,221,0,199,0,120,0,156,0,213,0,0,0,210,0,99,0,34,0,130,0,88,0,0,0,156,0,126,0,212,0,240,0,0,0,19,0,232,0,179,0,0,0,0,0,0,0,27,0,0,0,199,0,0,0,93,0,89,0,0,0,121,0,81,0,191,0,50,0,62,0,142,0,28,0,57,0,191,0,0,0,220,0,150,0,0,0,231,0,216,0,234,0,0,0,203,0,76,0,54,0,95,0,39,0,113,0,94,0,175,0,132,0,244,0,165,0,205,0,133,0,89,0,214,0,0,0,253,0,188,0,183,0,117,0,0,0,163,0,187,0,0,0,228,0,0,0,234,0,65,0,11,0,58,0,76,0,203,0,156,0,26,0,243,0,218,0,86,0,0,0,160,0,108,0,157,0,11,0,44,0,181,0,253,0,17,0,0,0,250,0,197,0,62,0,196,0,202,0,241,0,68,0,81,0,50,0,200,0,137,0,23,0,234,0,13,0,45,0,0,0,75,0,14,0,230,0,238,0,159,0,16,0,179,0,0,0,72,0,80,0,61,0,231,0,12,0,92,0,231,0,132,0,54,0,212,0,221,0,0,0,68,0,21,0,164,0,168,0,163,0,0,0,218,0,0,0,0,0,42,0,210,0,193,0,0,0,88,0,102,0,0,0,251,0,228,0,200,0,72,0,231,0,38,0,137,0,22,0,0,0,5,0,66,0,17,0,0,0,178,0,191,0,249,0,0,0,0,0,141,0,118,0,0,0,25,0,130,0,0,0,49,0,37,0,0,0,6,0,0,0,34,0,74,0,124,0,110,0,151,0,0,0,85,0,135,0,0,0,0,0,0,0,0,0,25,0,1,0,80,0,227,0,141,0,22,0,181,0,42,0,0,0,0,0,114,0,102,0,181,0,68,0,251,0,0,0,107,0,171,0,154,0,127,0,156,0,24,0,165,0,165,0,0,0,187,0,144,0,128,0,238,0,59,0,191,0,227,0,0,0,157,0,255,0,0,0,110,0,24,0,0,0,242,0,79,0,46,0,132,0,26,0,0,0,245,0,212,0,152,0,124,0,164,0,70,0,83,0,8,0,0,0,231,0,84,0,0,0,169,0,226,0,150,0,0,0,32,0,0,0,44,0,228,0,247,0,0,0,0,0,240,0,201,0,154,0,76,0,52,0,105,0,18,0,0,0,115,0,73,0,0,0,203,0,68,0,155,0,0,0,0,0,51,0,55,0,11,0,223,0,65,0,38,0,0,0,254,0,52,0,82,0,87,0,237,0,0,0,226,0,162,0,165,0,181,0,101,0,157,0);
signal scenario_full  : scenario_type := (135,31,167,31,184,31,142,31,142,30,181,31,5,31,76,31,88,31,228,31,228,30,206,31,154,31,245,31,245,30,201,31,45,31,154,31,184,31,182,31,182,30,141,31,117,31,177,31,89,31,189,31,189,30,193,31,121,31,121,30,121,29,121,28,161,31,180,31,180,30,91,31,164,31,178,31,152,31,207,31,207,30,174,31,196,31,196,30,196,29,196,31,180,31,235,31,205,31,82,31,82,30,104,31,145,31,54,31,80,31,128,31,138,31,166,31,167,31,54,31,123,31,240,31,240,30,240,29,13,31,61,31,239,31,130,31,91,31,135,31,205,31,244,31,19,31,202,31,202,30,68,31,254,31,116,31,116,30,116,29,98,31,185,31,181,31,213,31,178,31,186,31,201,31,38,31,208,31,118,31,171,31,171,30,171,29,171,28,42,31,210,31,50,31,91,31,35,31,17,31,235,31,235,30,6,31,69,31,14,31,61,31,61,30,130,31,52,31,52,30,52,29,211,31,37,31,182,31,133,31,138,31,243,31,116,31,116,30,64,31,129,31,45,31,61,31,61,30,221,31,205,31,205,30,156,31,156,30,156,29,24,31,98,31,77,31,242,31,172,31,128,31,128,30,107,31,28,31,69,31,154,31,112,31,112,30,245,31,231,31,129,31,196,31,247,31,247,30,55,31,184,31,220,31,220,30,97,31,74,31,74,30,123,31,136,31,148,31,226,31,147,31,216,31,167,31,85,31,12,31,234,31,234,30,234,29,44,31,245,31,245,30,48,31,50,31,19,31,36,31,22,31,179,31,207,31,190,31,190,30,221,31,28,31,130,31,151,31,76,31,206,31,203,31,2,31,209,31,78,31,138,31,106,31,106,30,112,31,195,31,235,31,235,30,195,31,71,31,114,31,114,30,238,31,30,31,97,31,51,31,191,31,75,31,23,31,35,31,35,30,250,31,157,31,254,31,232,31,231,31,25,31,82,31,236,31,113,31,57,31,57,30,67,31,67,30,172,31,248,31,1,31,156,31,74,31,74,30,252,31,251,31,203,31,203,30,203,29,9,31,34,31,121,31,203,31,162,31,162,30,86,31,1,31,105,31,163,31,157,31,25,31,123,31,48,31,139,31,129,31,129,30,13,31,181,31,179,31,45,31,45,30,181,31,235,31,195,31,150,31,150,30,158,31,158,30,25,31,25,30,217,31,217,30,217,29,54,31,165,31,143,31,143,30,143,29,192,31,241,31,241,30,249,31,103,31,122,31,160,31,100,31,159,31,105,31,84,31,84,30,221,31,213,31,216,31,140,31,237,31,173,31,29,31,87,31,8,31,252,31,105,31,228,31,228,30,222,31,37,31,86,31,35,31,195,31,81,31,53,31,22,31,100,31,156,31,156,30,252,31,71,31,148,31,138,31,18,31,18,30,50,31,50,30,50,29,161,31,27,31,92,31,5,31,49,31,206,31,56,31,65,31,36,31,204,31,61,31,61,30,39,31,189,31,110,31,253,31,253,30,133,31,137,31,137,30,28,31,28,30,20,31,20,30,92,31,44,31,103,31,182,31,93,31,251,31,69,31,160,31,234,31,234,30,139,31,126,31,105,31,224,31,199,31,199,30,88,31,118,31,93,31,111,31,111,30,81,31,176,31,251,31,116,31,99,31,99,30,15,31,15,30,114,31,158,31,158,30,158,29,158,28,130,31,34,31,173,31,173,30,56,31,210,31,124,31,236,31,135,31,153,31,37,31,247,31,33,31,178,31,178,30,190,31,119,31,119,30,243,31,161,31,140,31,20,31,17,31,65,31,146,31,192,31,22,31,202,31,175,31,158,31,221,31,199,31,120,31,156,31,213,31,213,30,210,31,99,31,34,31,130,31,88,31,88,30,156,31,126,31,212,31,240,31,240,30,19,31,232,31,179,31,179,30,179,29,179,28,27,31,27,30,199,31,199,30,93,31,89,31,89,30,121,31,81,31,191,31,50,31,62,31,142,31,28,31,57,31,191,31,191,30,220,31,150,31,150,30,231,31,216,31,234,31,234,30,203,31,76,31,54,31,95,31,39,31,113,31,94,31,175,31,132,31,244,31,165,31,205,31,133,31,89,31,214,31,214,30,253,31,188,31,183,31,117,31,117,30,163,31,187,31,187,30,228,31,228,30,234,31,65,31,11,31,58,31,76,31,203,31,156,31,26,31,243,31,218,31,86,31,86,30,160,31,108,31,157,31,11,31,44,31,181,31,253,31,17,31,17,30,250,31,197,31,62,31,196,31,202,31,241,31,68,31,81,31,50,31,200,31,137,31,23,31,234,31,13,31,45,31,45,30,75,31,14,31,230,31,238,31,159,31,16,31,179,31,179,30,72,31,80,31,61,31,231,31,12,31,92,31,231,31,132,31,54,31,212,31,221,31,221,30,68,31,21,31,164,31,168,31,163,31,163,30,218,31,218,30,218,29,42,31,210,31,193,31,193,30,88,31,102,31,102,30,251,31,228,31,200,31,72,31,231,31,38,31,137,31,22,31,22,30,5,31,66,31,17,31,17,30,178,31,191,31,249,31,249,30,249,29,141,31,118,31,118,30,25,31,130,31,130,30,49,31,37,31,37,30,6,31,6,30,34,31,74,31,124,31,110,31,151,31,151,30,85,31,135,31,135,30,135,29,135,28,135,27,25,31,1,31,80,31,227,31,141,31,22,31,181,31,42,31,42,30,42,29,114,31,102,31,181,31,68,31,251,31,251,30,107,31,171,31,154,31,127,31,156,31,24,31,165,31,165,31,165,30,187,31,144,31,128,31,238,31,59,31,191,31,227,31,227,30,157,31,255,31,255,30,110,31,24,31,24,30,242,31,79,31,46,31,132,31,26,31,26,30,245,31,212,31,152,31,124,31,164,31,70,31,83,31,8,31,8,30,231,31,84,31,84,30,169,31,226,31,150,31,150,30,32,31,32,30,44,31,228,31,247,31,247,30,247,29,240,31,201,31,154,31,76,31,52,31,105,31,18,31,18,30,115,31,73,31,73,30,203,31,68,31,155,31,155,30,155,29,51,31,55,31,11,31,223,31,65,31,38,31,38,30,254,31,52,31,82,31,87,31,237,31,237,30,226,31,162,31,165,31,181,31,101,31,157,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
