-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_308 is
end project_tb_308;

architecture project_tb_arch_308 of project_tb_308 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 384;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (244,0,154,0,0,0,234,0,96,0,23,0,27,0,145,0,65,0,143,0,34,0,224,0,77,0,210,0,206,0,0,0,123,0,158,0,0,0,174,0,0,0,37,0,149,0,0,0,157,0,206,0,230,0,160,0,71,0,0,0,89,0,0,0,2,0,145,0,56,0,0,0,0,0,253,0,192,0,4,0,0,0,0,0,124,0,36,0,113,0,188,0,179,0,0,0,162,0,78,0,115,0,198,0,89,0,0,0,0,0,169,0,31,0,4,0,39,0,0,0,102,0,7,0,0,0,26,0,125,0,146,0,151,0,19,0,195,0,246,0,205,0,56,0,194,0,250,0,54,0,178,0,211,0,5,0,153,0,84,0,39,0,8,0,0,0,0,0,12,0,149,0,8,0,61,0,0,0,195,0,202,0,54,0,146,0,95,0,19,0,173,0,28,0,163,0,151,0,139,0,139,0,194,0,253,0,65,0,106,0,0,0,0,0,10,0,227,0,244,0,16,0,0,0,0,0,237,0,152,0,91,0,215,0,30,0,1,0,222,0,244,0,24,0,0,0,12,0,44,0,153,0,0,0,0,0,232,0,178,0,169,0,0,0,0,0,130,0,25,0,127,0,34,0,19,0,0,0,107,0,138,0,220,0,0,0,137,0,0,0,55,0,45,0,233,0,0,0,220,0,0,0,155,0,27,0,22,0,4,0,212,0,225,0,195,0,183,0,0,0,145,0,138,0,0,0,227,0,0,0,0,0,75,0,92,0,99,0,0,0,60,0,75,0,223,0,216,0,27,0,138,0,251,0,108,0,231,0,244,0,0,0,31,0,222,0,0,0,146,0,147,0,0,0,160,0,234,0,71,0,123,0,107,0,160,0,7,0,65,0,194,0,80,0,2,0,69,0,250,0,168,0,0,0,83,0,219,0,58,0,90,0,216,0,196,0,89,0,85,0,243,0,108,0,0,0,72,0,124,0,196,0,171,0,0,0,46,0,210,0,182,0,124,0,234,0,73,0,43,0,241,0,40,0,0,0,239,0,68,0,216,0,0,0,39,0,199,0,215,0,197,0,44,0,58,0,0,0,0,0,0,0,182,0,121,0,0,0,121,0,0,0,183,0,77,0,213,0,77,0,107,0,50,0,84,0,0,0,166,0,238,0,252,0,100,0,183,0,0,0,105,0,0,0,0,0,187,0,0,0,80,0,0,0,62,0,161,0,249,0,72,0,225,0,0,0,214,0,251,0,0,0,54,0,247,0,56,0,202,0,125,0,0,0,173,0,227,0,75,0,165,0,0,0,161,0,253,0,2,0,119,0,193,0,0,0,157,0,8,0,174,0,0,0,11,0,218,0,214,0,91,0,3,0,55,0,109,0,9,0,223,0,0,0,136,0,236,0,0,0,0,0,114,0,246,0,101,0,212,0,0,0,199,0,147,0,227,0,79,0,0,0,0,0,147,0,176,0,68,0,133,0,30,0,206,0,27,0,0,0,0,0,220,0,123,0,0,0,93,0,184,0,170,0,185,0,88,0,21,0,152,0,197,0,10,0,216,0,199,0,207,0,74,0,31,0,204,0,71,0,172,0,0,0,0,0,83,0,0,0,29,0,0,0,0,0,157,0,134,0,0,0,171,0,131,0,234,0,216,0,0,0,167,0,11,0,0,0,131,0,116,0,0,0,229,0,95,0,0,0,60,0,186,0,0,0,160,0,238,0,163,0,51,0,53,0,0,0);
signal scenario_full  : scenario_type := (244,31,154,31,154,30,234,31,96,31,23,31,27,31,145,31,65,31,143,31,34,31,224,31,77,31,210,31,206,31,206,30,123,31,158,31,158,30,174,31,174,30,37,31,149,31,149,30,157,31,206,31,230,31,160,31,71,31,71,30,89,31,89,30,2,31,145,31,56,31,56,30,56,29,253,31,192,31,4,31,4,30,4,29,124,31,36,31,113,31,188,31,179,31,179,30,162,31,78,31,115,31,198,31,89,31,89,30,89,29,169,31,31,31,4,31,39,31,39,30,102,31,7,31,7,30,26,31,125,31,146,31,151,31,19,31,195,31,246,31,205,31,56,31,194,31,250,31,54,31,178,31,211,31,5,31,153,31,84,31,39,31,8,31,8,30,8,29,12,31,149,31,8,31,61,31,61,30,195,31,202,31,54,31,146,31,95,31,19,31,173,31,28,31,163,31,151,31,139,31,139,31,194,31,253,31,65,31,106,31,106,30,106,29,10,31,227,31,244,31,16,31,16,30,16,29,237,31,152,31,91,31,215,31,30,31,1,31,222,31,244,31,24,31,24,30,12,31,44,31,153,31,153,30,153,29,232,31,178,31,169,31,169,30,169,29,130,31,25,31,127,31,34,31,19,31,19,30,107,31,138,31,220,31,220,30,137,31,137,30,55,31,45,31,233,31,233,30,220,31,220,30,155,31,27,31,22,31,4,31,212,31,225,31,195,31,183,31,183,30,145,31,138,31,138,30,227,31,227,30,227,29,75,31,92,31,99,31,99,30,60,31,75,31,223,31,216,31,27,31,138,31,251,31,108,31,231,31,244,31,244,30,31,31,222,31,222,30,146,31,147,31,147,30,160,31,234,31,71,31,123,31,107,31,160,31,7,31,65,31,194,31,80,31,2,31,69,31,250,31,168,31,168,30,83,31,219,31,58,31,90,31,216,31,196,31,89,31,85,31,243,31,108,31,108,30,72,31,124,31,196,31,171,31,171,30,46,31,210,31,182,31,124,31,234,31,73,31,43,31,241,31,40,31,40,30,239,31,68,31,216,31,216,30,39,31,199,31,215,31,197,31,44,31,58,31,58,30,58,29,58,28,182,31,121,31,121,30,121,31,121,30,183,31,77,31,213,31,77,31,107,31,50,31,84,31,84,30,166,31,238,31,252,31,100,31,183,31,183,30,105,31,105,30,105,29,187,31,187,30,80,31,80,30,62,31,161,31,249,31,72,31,225,31,225,30,214,31,251,31,251,30,54,31,247,31,56,31,202,31,125,31,125,30,173,31,227,31,75,31,165,31,165,30,161,31,253,31,2,31,119,31,193,31,193,30,157,31,8,31,174,31,174,30,11,31,218,31,214,31,91,31,3,31,55,31,109,31,9,31,223,31,223,30,136,31,236,31,236,30,236,29,114,31,246,31,101,31,212,31,212,30,199,31,147,31,227,31,79,31,79,30,79,29,147,31,176,31,68,31,133,31,30,31,206,31,27,31,27,30,27,29,220,31,123,31,123,30,93,31,184,31,170,31,185,31,88,31,21,31,152,31,197,31,10,31,216,31,199,31,207,31,74,31,31,31,204,31,71,31,172,31,172,30,172,29,83,31,83,30,29,31,29,30,29,29,157,31,134,31,134,30,171,31,131,31,234,31,216,31,216,30,167,31,11,31,11,30,131,31,116,31,116,30,229,31,95,31,95,30,60,31,186,31,186,30,160,31,238,31,163,31,51,31,53,31,53,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
