-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_275 is
end project_tb_275;

architecture project_tb_arch_275 of project_tb_275 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 924;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,203,0,52,0,54,0,0,0,74,0,0,0,8,0,241,0,7,0,86,0,12,0,178,0,78,0,138,0,55,0,164,0,17,0,33,0,0,0,188,0,175,0,0,0,58,0,206,0,151,0,103,0,138,0,0,0,141,0,142,0,146,0,0,0,40,0,1,0,0,0,91,0,108,0,187,0,147,0,107,0,0,0,229,0,0,0,0,0,101,0,44,0,188,0,142,0,0,0,100,0,136,0,81,0,43,0,166,0,203,0,185,0,0,0,200,0,124,0,0,0,0,0,229,0,120,0,146,0,134,0,108,0,144,0,162,0,34,0,179,0,214,0,17,0,0,0,102,0,121,0,13,0,225,0,41,0,0,0,0,0,100,0,98,0,141,0,34,0,0,0,119,0,118,0,30,0,0,0,31,0,0,0,0,0,83,0,91,0,235,0,79,0,175,0,14,0,135,0,8,0,116,0,46,0,0,0,0,0,1,0,93,0,3,0,111,0,77,0,135,0,124,0,0,0,0,0,0,0,214,0,139,0,91,0,41,0,0,0,0,0,245,0,150,0,16,0,13,0,138,0,147,0,148,0,0,0,119,0,143,0,0,0,118,0,145,0,238,0,39,0,193,0,201,0,163,0,219,0,155,0,207,0,43,0,232,0,11,0,227,0,163,0,214,0,3,0,244,0,0,0,208,0,203,0,189,0,187,0,208,0,186,0,118,0,0,0,120,0,30,0,64,0,106,0,123,0,0,0,215,0,255,0,152,0,28,0,165,0,105,0,254,0,69,0,180,0,59,0,0,0,202,0,101,0,151,0,251,0,44,0,0,0,0,0,141,0,46,0,248,0,182,0,83,0,249,0,125,0,49,0,184,0,43,0,13,0,0,0,247,0,0,0,49,0,0,0,233,0,115,0,108,0,145,0,187,0,97,0,112,0,79,0,236,0,131,0,37,0,214,0,114,0,46,0,186,0,193,0,13,0,183,0,0,0,180,0,210,0,135,0,17,0,122,0,231,0,96,0,196,0,155,0,145,0,26,0,253,0,0,0,6,0,189,0,130,0,75,0,75,0,0,0,0,0,217,0,0,0,132,0,45,0,212,0,135,0,139,0,7,0,0,0,0,0,66,0,0,0,163,0,53,0,183,0,64,0,0,0,0,0,152,0,0,0,100,0,120,0,0,0,47,0,156,0,0,0,52,0,234,0,0,0,206,0,137,0,141,0,114,0,180,0,220,0,143,0,132,0,0,0,97,0,81,0,119,0,220,0,183,0,73,0,19,0,26,0,213,0,173,0,163,0,40,0,157,0,97,0,146,0,158,0,0,0,205,0,0,0,42,0,120,0,143,0,170,0,56,0,60,0,95,0,93,0,77,0,229,0,236,0,237,0,43,0,6,0,45,0,124,0,95,0,0,0,124,0,0,0,177,0,147,0,3,0,0,0,143,0,0,0,34,0,96,0,0,0,75,0,0,0,146,0,40,0,0,0,42,0,59,0,247,0,12,0,119,0,64,0,2,0,132,0,172,0,250,0,122,0,96,0,85,0,211,0,175,0,126,0,216,0,226,0,235,0,0,0,14,0,0,0,141,0,0,0,156,0,144,0,194,0,225,0,189,0,186,0,114,0,24,0,32,0,176,0,187,0,0,0,99,0,0,0,0,0,196,0,22,0,116,0,29,0,0,0,166,0,59,0,204,0,64,0,234,0,15,0,24,0,0,0,0,0,0,0,133,0,33,0,168,0,144,0,0,0,0,0,18,0,132,0,105,0,94,0,0,0,121,0,0,0,0,0,0,0,92,0,214,0,179,0,44,0,31,0,14,0,55,0,0,0,156,0,0,0,105,0,36,0,136,0,111,0,161,0,171,0,194,0,128,0,78,0,142,0,200,0,138,0,9,0,0,0,96,0,0,0,161,0,0,0,71,0,21,0,103,0,0,0,201,0,39,0,179,0,138,0,204,0,153,0,24,0,16,0,230,0,57,0,59,0,0,0,116,0,0,0,152,0,245,0,0,0,101,0,0,0,199,0,0,0,101,0,93,0,205,0,131,0,191,0,131,0,118,0,4,0,48,0,76,0,8,0,0,0,0,0,0,0,137,0,209,0,19,0,67,0,145,0,83,0,64,0,0,0,149,0,0,0,177,0,45,0,55,0,96,0,112,0,85,0,53,0,0,0,250,0,62,0,156,0,151,0,0,0,163,0,167,0,166,0,204,0,126,0,253,0,0,0,118,0,192,0,83,0,176,0,59,0,198,0,203,0,0,0,0,0,160,0,0,0,195,0,249,0,0,0,36,0,13,0,0,0,244,0,107,0,29,0,77,0,0,0,40,0,92,0,0,0,8,0,167,0,106,0,113,0,0,0,157,0,111,0,31,0,34,0,20,0,28,0,130,0,199,0,110,0,120,0,211,0,144,0,79,0,0,0,74,0,235,0,26,0,180,0,0,0,200,0,67,0,30,0,101,0,221,0,240,0,167,0,0,0,179,0,178,0,0,0,0,0,0,0,0,0,159,0,250,0,159,0,49,0,0,0,217,0,212,0,12,0,235,0,173,0,118,0,208,0,178,0,65,0,26,0,116,0,21,0,95,0,144,0,221,0,93,0,1,0,132,0,12,0,71,0,202,0,0,0,168,0,0,0,41,0,0,0,228,0,134,0,147,0,191,0,200,0,37,0,74,0,0,0,120,0,98,0,138,0,113,0,178,0,98,0,0,0,54,0,233,0,217,0,7,0,0,0,0,0,183,0,50,0,10,0,78,0,0,0,0,0,111,0,145,0,253,0,6,0,172,0,109,0,169,0,54,0,0,0,2,0,0,0,35,0,0,0,137,0,211,0,0,0,147,0,46,0,113,0,165,0,57,0,138,0,205,0,71,0,0,0,106,0,0,0,2,0,208,0,57,0,120,0,16,0,71,0,230,0,0,0,0,0,220,0,131,0,101,0,166,0,0,0,4,0,18,0,92,0,0,0,4,0,207,0,0,0,148,0,34,0,125,0,8,0,238,0,235,0,162,0,144,0,173,0,0,0,0,0,0,0,179,0,87,0,124,0,39,0,83,0,180,0,168,0,39,0,225,0,48,0,62,0,255,0,56,0,0,0,142,0,148,0,118,0,71,0,0,0,50,0,8,0,0,0,96,0,22,0,0,0,0,0,0,0,0,0,0,0,233,0,158,0,0,0,86,0,110,0,68,0,170,0,161,0,16,0,204,0,167,0,212,0,162,0,236,0,0,0,0,0,158,0,12,0,55,0,225,0,157,0,209,0,143,0,149,0,123,0,0,0,0,0,0,0,61,0,17,0,62,0,171,0,152,0,255,0,64,0,70,0,81,0,0,0,254,0,50,0,170,0,215,0,0,0,198,0,0,0,230,0,115,0,131,0,222,0,64,0,140,0,149,0,6,0,0,0,187,0,53,0,91,0,0,0,255,0,151,0,0,0,170,0,18,0,106,0,0,0,40,0,61,0,240,0,149,0,42,0,250,0,165,0,223,0,229,0,111,0,68,0,164,0,168,0,59,0,0,0,177,0,253,0,38,0,159,0,93,0,38,0,177,0,105,0,0,0,0,0,0,0,226,0,238,0,92,0,18,0,0,0,37,0,0,0,133,0,0,0,0,0,7,0,39,0,85,0,147,0,254,0,250,0,124,0,12,0,131,0,82,0,154,0,51,0,153,0,80,0,231,0,0,0,127,0,0,0,172,0,189,0,0,0,65,0,0,0,77,0,219,0,43,0,223,0,38,0,0,0,36,0,0,0,254,0,0,0,33,0,156,0,178,0,245,0,211,0,213,0,0,0,111,0,215,0,112,0,143,0,0,0,127,0,0,0,118,0,3,0,78,0,4,0,15,0,122,0,0,0,0,0,0,0,234,0,27,0,63,0,47,0,143,0,71,0,210,0,209,0,180,0,114,0,0,0,0,0,120,0,221,0,133,0,10,0,184,0,84,0,226,0,28,0,160,0,0,0,108,0,115,0,104,0,65,0,102,0,0,0,0,0,186,0,80,0,247,0,195,0,97,0,165,0,0,0,166,0,8,0,54,0,37,0,220,0,136,0,0,0,65,0,204,0,228,0,0,0,44,0,120,0,23,0,182,0,0,0,114,0,0,0,207,0,206,0,168,0,4,0,21,0,0,0,90,0,0,0);
signal scenario_full  : scenario_type := (0,0,203,31,52,31,54,31,54,30,74,31,74,30,8,31,241,31,7,31,86,31,12,31,178,31,78,31,138,31,55,31,164,31,17,31,33,31,33,30,188,31,175,31,175,30,58,31,206,31,151,31,103,31,138,31,138,30,141,31,142,31,146,31,146,30,40,31,1,31,1,30,91,31,108,31,187,31,147,31,107,31,107,30,229,31,229,30,229,29,101,31,44,31,188,31,142,31,142,30,100,31,136,31,81,31,43,31,166,31,203,31,185,31,185,30,200,31,124,31,124,30,124,29,229,31,120,31,146,31,134,31,108,31,144,31,162,31,34,31,179,31,214,31,17,31,17,30,102,31,121,31,13,31,225,31,41,31,41,30,41,29,100,31,98,31,141,31,34,31,34,30,119,31,118,31,30,31,30,30,31,31,31,30,31,29,83,31,91,31,235,31,79,31,175,31,14,31,135,31,8,31,116,31,46,31,46,30,46,29,1,31,93,31,3,31,111,31,77,31,135,31,124,31,124,30,124,29,124,28,214,31,139,31,91,31,41,31,41,30,41,29,245,31,150,31,16,31,13,31,138,31,147,31,148,31,148,30,119,31,143,31,143,30,118,31,145,31,238,31,39,31,193,31,201,31,163,31,219,31,155,31,207,31,43,31,232,31,11,31,227,31,163,31,214,31,3,31,244,31,244,30,208,31,203,31,189,31,187,31,208,31,186,31,118,31,118,30,120,31,30,31,64,31,106,31,123,31,123,30,215,31,255,31,152,31,28,31,165,31,105,31,254,31,69,31,180,31,59,31,59,30,202,31,101,31,151,31,251,31,44,31,44,30,44,29,141,31,46,31,248,31,182,31,83,31,249,31,125,31,49,31,184,31,43,31,13,31,13,30,247,31,247,30,49,31,49,30,233,31,115,31,108,31,145,31,187,31,97,31,112,31,79,31,236,31,131,31,37,31,214,31,114,31,46,31,186,31,193,31,13,31,183,31,183,30,180,31,210,31,135,31,17,31,122,31,231,31,96,31,196,31,155,31,145,31,26,31,253,31,253,30,6,31,189,31,130,31,75,31,75,31,75,30,75,29,217,31,217,30,132,31,45,31,212,31,135,31,139,31,7,31,7,30,7,29,66,31,66,30,163,31,53,31,183,31,64,31,64,30,64,29,152,31,152,30,100,31,120,31,120,30,47,31,156,31,156,30,52,31,234,31,234,30,206,31,137,31,141,31,114,31,180,31,220,31,143,31,132,31,132,30,97,31,81,31,119,31,220,31,183,31,73,31,19,31,26,31,213,31,173,31,163,31,40,31,157,31,97,31,146,31,158,31,158,30,205,31,205,30,42,31,120,31,143,31,170,31,56,31,60,31,95,31,93,31,77,31,229,31,236,31,237,31,43,31,6,31,45,31,124,31,95,31,95,30,124,31,124,30,177,31,147,31,3,31,3,30,143,31,143,30,34,31,96,31,96,30,75,31,75,30,146,31,40,31,40,30,42,31,59,31,247,31,12,31,119,31,64,31,2,31,132,31,172,31,250,31,122,31,96,31,85,31,211,31,175,31,126,31,216,31,226,31,235,31,235,30,14,31,14,30,141,31,141,30,156,31,144,31,194,31,225,31,189,31,186,31,114,31,24,31,32,31,176,31,187,31,187,30,99,31,99,30,99,29,196,31,22,31,116,31,29,31,29,30,166,31,59,31,204,31,64,31,234,31,15,31,24,31,24,30,24,29,24,28,133,31,33,31,168,31,144,31,144,30,144,29,18,31,132,31,105,31,94,31,94,30,121,31,121,30,121,29,121,28,92,31,214,31,179,31,44,31,31,31,14,31,55,31,55,30,156,31,156,30,105,31,36,31,136,31,111,31,161,31,171,31,194,31,128,31,78,31,142,31,200,31,138,31,9,31,9,30,96,31,96,30,161,31,161,30,71,31,21,31,103,31,103,30,201,31,39,31,179,31,138,31,204,31,153,31,24,31,16,31,230,31,57,31,59,31,59,30,116,31,116,30,152,31,245,31,245,30,101,31,101,30,199,31,199,30,101,31,93,31,205,31,131,31,191,31,131,31,118,31,4,31,48,31,76,31,8,31,8,30,8,29,8,28,137,31,209,31,19,31,67,31,145,31,83,31,64,31,64,30,149,31,149,30,177,31,45,31,55,31,96,31,112,31,85,31,53,31,53,30,250,31,62,31,156,31,151,31,151,30,163,31,167,31,166,31,204,31,126,31,253,31,253,30,118,31,192,31,83,31,176,31,59,31,198,31,203,31,203,30,203,29,160,31,160,30,195,31,249,31,249,30,36,31,13,31,13,30,244,31,107,31,29,31,77,31,77,30,40,31,92,31,92,30,8,31,167,31,106,31,113,31,113,30,157,31,111,31,31,31,34,31,20,31,28,31,130,31,199,31,110,31,120,31,211,31,144,31,79,31,79,30,74,31,235,31,26,31,180,31,180,30,200,31,67,31,30,31,101,31,221,31,240,31,167,31,167,30,179,31,178,31,178,30,178,29,178,28,178,27,159,31,250,31,159,31,49,31,49,30,217,31,212,31,12,31,235,31,173,31,118,31,208,31,178,31,65,31,26,31,116,31,21,31,95,31,144,31,221,31,93,31,1,31,132,31,12,31,71,31,202,31,202,30,168,31,168,30,41,31,41,30,228,31,134,31,147,31,191,31,200,31,37,31,74,31,74,30,120,31,98,31,138,31,113,31,178,31,98,31,98,30,54,31,233,31,217,31,7,31,7,30,7,29,183,31,50,31,10,31,78,31,78,30,78,29,111,31,145,31,253,31,6,31,172,31,109,31,169,31,54,31,54,30,2,31,2,30,35,31,35,30,137,31,211,31,211,30,147,31,46,31,113,31,165,31,57,31,138,31,205,31,71,31,71,30,106,31,106,30,2,31,208,31,57,31,120,31,16,31,71,31,230,31,230,30,230,29,220,31,131,31,101,31,166,31,166,30,4,31,18,31,92,31,92,30,4,31,207,31,207,30,148,31,34,31,125,31,8,31,238,31,235,31,162,31,144,31,173,31,173,30,173,29,173,28,179,31,87,31,124,31,39,31,83,31,180,31,168,31,39,31,225,31,48,31,62,31,255,31,56,31,56,30,142,31,148,31,118,31,71,31,71,30,50,31,8,31,8,30,96,31,22,31,22,30,22,29,22,28,22,27,22,26,233,31,158,31,158,30,86,31,110,31,68,31,170,31,161,31,16,31,204,31,167,31,212,31,162,31,236,31,236,30,236,29,158,31,12,31,55,31,225,31,157,31,209,31,143,31,149,31,123,31,123,30,123,29,123,28,61,31,17,31,62,31,171,31,152,31,255,31,64,31,70,31,81,31,81,30,254,31,50,31,170,31,215,31,215,30,198,31,198,30,230,31,115,31,131,31,222,31,64,31,140,31,149,31,6,31,6,30,187,31,53,31,91,31,91,30,255,31,151,31,151,30,170,31,18,31,106,31,106,30,40,31,61,31,240,31,149,31,42,31,250,31,165,31,223,31,229,31,111,31,68,31,164,31,168,31,59,31,59,30,177,31,253,31,38,31,159,31,93,31,38,31,177,31,105,31,105,30,105,29,105,28,226,31,238,31,92,31,18,31,18,30,37,31,37,30,133,31,133,30,133,29,7,31,39,31,85,31,147,31,254,31,250,31,124,31,12,31,131,31,82,31,154,31,51,31,153,31,80,31,231,31,231,30,127,31,127,30,172,31,189,31,189,30,65,31,65,30,77,31,219,31,43,31,223,31,38,31,38,30,36,31,36,30,254,31,254,30,33,31,156,31,178,31,245,31,211,31,213,31,213,30,111,31,215,31,112,31,143,31,143,30,127,31,127,30,118,31,3,31,78,31,4,31,15,31,122,31,122,30,122,29,122,28,234,31,27,31,63,31,47,31,143,31,71,31,210,31,209,31,180,31,114,31,114,30,114,29,120,31,221,31,133,31,10,31,184,31,84,31,226,31,28,31,160,31,160,30,108,31,115,31,104,31,65,31,102,31,102,30,102,29,186,31,80,31,247,31,195,31,97,31,165,31,165,30,166,31,8,31,54,31,37,31,220,31,136,31,136,30,65,31,204,31,228,31,228,30,44,31,120,31,23,31,182,31,182,30,114,31,114,30,207,31,206,31,168,31,4,31,21,31,21,30,90,31,90,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
