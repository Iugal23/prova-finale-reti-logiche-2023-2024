-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_768 is
end project_tb_768;

architecture project_tb_arch_768 of project_tb_768 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 814;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,65,0,57,0,79,0,0,0,0,0,0,0,192,0,121,0,89,0,74,0,100,0,64,0,117,0,235,0,134,0,166,0,0,0,235,0,172,0,136,0,162,0,98,0,214,0,43,0,196,0,214,0,120,0,179,0,0,0,236,0,188,0,60,0,24,0,231,0,202,0,0,0,25,0,51,0,235,0,132,0,89,0,100,0,41,0,115,0,152,0,250,0,240,0,153,0,143,0,0,0,12,0,57,0,60,0,0,0,0,0,211,0,11,0,64,0,8,0,0,0,33,0,215,0,239,0,115,0,8,0,79,0,120,0,0,0,0,0,149,0,94,0,69,0,55,0,0,0,0,0,230,0,168,0,0,0,4,0,186,0,168,0,203,0,0,0,84,0,9,0,0,0,167,0,0,0,193,0,161,0,135,0,145,0,238,0,0,0,65,0,0,0,16,0,216,0,0,0,170,0,0,0,156,0,120,0,246,0,133,0,0,0,224,0,154,0,155,0,31,0,54,0,138,0,9,0,59,0,223,0,102,0,199,0,125,0,183,0,128,0,67,0,143,0,88,0,202,0,164,0,0,0,145,0,0,0,0,0,120,0,193,0,96,0,72,0,220,0,79,0,0,0,235,0,206,0,75,0,138,0,249,0,105,0,67,0,18,0,53,0,0,0,87,0,114,0,2,0,103,0,0,0,177,0,189,0,170,0,35,0,202,0,34,0,12,0,0,0,71,0,0,0,92,0,0,0,115,0,221,0,99,0,21,0,40,0,32,0,76,0,61,0,231,0,124,0,69,0,114,0,58,0,134,0,15,0,164,0,136,0,143,0,87,0,147,0,238,0,185,0,74,0,108,0,167,0,226,0,107,0,0,0,34,0,97,0,117,0,45,0,140,0,154,0,21,0,156,0,78,0,17,0,0,0,82,0,0,0,112,0,179,0,13,0,162,0,32,0,28,0,54,0,100,0,250,0,0,0,80,0,0,0,134,0,27,0,0,0,43,0,87,0,0,0,199,0,239,0,136,0,1,0,0,0,44,0,3,0,0,0,0,0,170,0,167,0,249,0,94,0,0,0,189,0,175,0,97,0,69,0,52,0,13,0,166,0,210,0,131,0,20,0,0,0,100,0,90,0,138,0,0,0,246,0,166,0,30,0,80,0,247,0,225,0,0,0,0,0,206,0,180,0,0,0,0,0,40,0,180,0,10,0,111,0,71,0,72,0,0,0,18,0,79,0,136,0,223,0,146,0,223,0,20,0,190,0,106,0,56,0,0,0,159,0,230,0,0,0,144,0,239,0,19,0,37,0,178,0,147,0,174,0,254,0,84,0,134,0,5,0,223,0,32,0,144,0,174,0,18,0,41,0,0,0,39,0,35,0,97,0,223,0,219,0,0,0,0,0,197,0,23,0,213,0,155,0,60,0,147,0,215,0,159,0,0,0,19,0,128,0,171,0,202,0,30,0,118,0,0,0,94,0,0,0,0,0,170,0,207,0,140,0,0,0,185,0,50,0,0,0,0,0,0,0,0,0,220,0,135,0,134,0,19,0,159,0,173,0,97,0,84,0,216,0,53,0,213,0,245,0,141,0,56,0,0,0,0,0,207,0,252,0,0,0,2,0,229,0,113,0,196,0,52,0,202,0,193,0,0,0,99,0,193,0,67,0,162,0,0,0,100,0,200,0,228,0,101,0,107,0,109,0,0,0,61,0,0,0,116,0,7,0,14,0,212,0,77,0,73,0,0,0,5,0,184,0,184,0,0,0,4,0,94,0,66,0,0,0,199,0,139,0,180,0,75,0,194,0,0,0,248,0,106,0,171,0,43,0,141,0,0,0,0,0,194,0,57,0,78,0,104,0,73,0,241,0,58,0,55,0,218,0,55,0,13,0,37,0,52,0,0,0,230,0,243,0,82,0,11,0,0,0,0,0,171,0,12,0,201,0,38,0,3,0,197,0,176,0,0,0,10,0,0,0,251,0,124,0,64,0,0,0,57,0,70,0,0,0,206,0,162,0,243,0,0,0,72,0,0,0,97,0,20,0,141,0,234,0,88,0,127,0,234,0,248,0,83,0,82,0,40,0,78,0,0,0,24,0,119,0,0,0,2,0,0,0,0,0,237,0,154,0,39,0,0,0,95,0,22,0,47,0,238,0,193,0,75,0,47,0,184,0,98,0,30,0,0,0,136,0,36,0,151,0,15,0,130,0,0,0,0,0,20,0,51,0,110,0,135,0,92,0,0,0,90,0,109,0,0,0,231,0,247,0,80,0,108,0,139,0,12,0,14,0,0,0,33,0,248,0,248,0,57,0,233,0,146,0,0,0,232,0,132,0,199,0,97,0,152,0,10,0,251,0,58,0,167,0,17,0,30,0,201,0,44,0,206,0,194,0,138,0,207,0,216,0,0,0,24,0,103,0,106,0,107,0,78,0,235,0,171,0,18,0,98,0,47,0,2,0,183,0,68,0,39,0,103,0,0,0,128,0,253,0,29,0,208,0,105,0,0,0,0,0,0,0,0,0,173,0,0,0,92,0,210,0,131,0,93,0,189,0,186,0,67,0,144,0,81,0,73,0,0,0,0,0,25,0,88,0,0,0,65,0,89,0,72,0,240,0,0,0,34,0,177,0,224,0,92,0,0,0,123,0,159,0,239,0,178,0,95,0,0,0,152,0,204,0,96,0,28,0,0,0,0,0,223,0,72,0,53,0,0,0,0,0,31,0,244,0,0,0,121,0,63,0,47,0,26,0,0,0,236,0,241,0,180,0,96,0,66,0,0,0,113,0,236,0,190,0,0,0,224,0,105,0,114,0,14,0,9,0,234,0,236,0,86,0,0,0,217,0,217,0,179,0,84,0,65,0,239,0,94,0,237,0,177,0,97,0,235,0,200,0,60,0,240,0,18,0,240,0,181,0,143,0,111,0,103,0,162,0,164,0,172,0,0,0,22,0,245,0,248,0,0,0,100,0,53,0,0,0,96,0,129,0,111,0,205,0,15,0,64,0,233,0,67,0,115,0,0,0,130,0,16,0,155,0,127,0,193,0,4,0,41,0,61,0,231,0,0,0,46,0,4,0,241,0,116,0,183,0,0,0,0,0,191,0,254,0,189,0,51,0,214,0,240,0,127,0,244,0,102,0,152,0,142,0,0,0,58,0,211,0,0,0,218,0,0,0,0,0,0,0,0,0,202,0,15,0,251,0,0,0,94,0,28,0,146,0,137,0,94,0,146,0,0,0,107,0,255,0,214,0,120,0,234,0,117,0,181,0,125,0,94,0,0,0,101,0,114,0,137,0,0,0,72,0,0,0,168,0,240,0,142,0,0,0,22,0,6,0,98,0,0,0,67,0,104,0,42,0,93,0,0,0,212,0,0,0,231,0,4,0,133,0,148,0,40,0,172,0,126,0,197,0,241,0,0,0,80,0,0,0,145,0,157,0,114,0,155,0,43,0,0,0,0,0,133,0,177,0,237,0,171,0,0,0,243,0,73,0,209,0,14,0,124,0,56,0,142,0,65,0,19,0,165,0,11,0,0,0,119,0,220,0,111,0,195,0,113,0,0,0,0,0,76,0,45,0,195,0,254,0,69,0,144,0,47,0,225,0,159,0,16,0,241,0,224,0,58,0,193,0,95,0,92,0,181,0,153,0,124,0,181,0);
signal scenario_full  : scenario_type := (0,0,65,31,57,31,79,31,79,30,79,29,79,28,192,31,121,31,89,31,74,31,100,31,64,31,117,31,235,31,134,31,166,31,166,30,235,31,172,31,136,31,162,31,98,31,214,31,43,31,196,31,214,31,120,31,179,31,179,30,236,31,188,31,60,31,24,31,231,31,202,31,202,30,25,31,51,31,235,31,132,31,89,31,100,31,41,31,115,31,152,31,250,31,240,31,153,31,143,31,143,30,12,31,57,31,60,31,60,30,60,29,211,31,11,31,64,31,8,31,8,30,33,31,215,31,239,31,115,31,8,31,79,31,120,31,120,30,120,29,149,31,94,31,69,31,55,31,55,30,55,29,230,31,168,31,168,30,4,31,186,31,168,31,203,31,203,30,84,31,9,31,9,30,167,31,167,30,193,31,161,31,135,31,145,31,238,31,238,30,65,31,65,30,16,31,216,31,216,30,170,31,170,30,156,31,120,31,246,31,133,31,133,30,224,31,154,31,155,31,31,31,54,31,138,31,9,31,59,31,223,31,102,31,199,31,125,31,183,31,128,31,67,31,143,31,88,31,202,31,164,31,164,30,145,31,145,30,145,29,120,31,193,31,96,31,72,31,220,31,79,31,79,30,235,31,206,31,75,31,138,31,249,31,105,31,67,31,18,31,53,31,53,30,87,31,114,31,2,31,103,31,103,30,177,31,189,31,170,31,35,31,202,31,34,31,12,31,12,30,71,31,71,30,92,31,92,30,115,31,221,31,99,31,21,31,40,31,32,31,76,31,61,31,231,31,124,31,69,31,114,31,58,31,134,31,15,31,164,31,136,31,143,31,87,31,147,31,238,31,185,31,74,31,108,31,167,31,226,31,107,31,107,30,34,31,97,31,117,31,45,31,140,31,154,31,21,31,156,31,78,31,17,31,17,30,82,31,82,30,112,31,179,31,13,31,162,31,32,31,28,31,54,31,100,31,250,31,250,30,80,31,80,30,134,31,27,31,27,30,43,31,87,31,87,30,199,31,239,31,136,31,1,31,1,30,44,31,3,31,3,30,3,29,170,31,167,31,249,31,94,31,94,30,189,31,175,31,97,31,69,31,52,31,13,31,166,31,210,31,131,31,20,31,20,30,100,31,90,31,138,31,138,30,246,31,166,31,30,31,80,31,247,31,225,31,225,30,225,29,206,31,180,31,180,30,180,29,40,31,180,31,10,31,111,31,71,31,72,31,72,30,18,31,79,31,136,31,223,31,146,31,223,31,20,31,190,31,106,31,56,31,56,30,159,31,230,31,230,30,144,31,239,31,19,31,37,31,178,31,147,31,174,31,254,31,84,31,134,31,5,31,223,31,32,31,144,31,174,31,18,31,41,31,41,30,39,31,35,31,97,31,223,31,219,31,219,30,219,29,197,31,23,31,213,31,155,31,60,31,147,31,215,31,159,31,159,30,19,31,128,31,171,31,202,31,30,31,118,31,118,30,94,31,94,30,94,29,170,31,207,31,140,31,140,30,185,31,50,31,50,30,50,29,50,28,50,27,220,31,135,31,134,31,19,31,159,31,173,31,97,31,84,31,216,31,53,31,213,31,245,31,141,31,56,31,56,30,56,29,207,31,252,31,252,30,2,31,229,31,113,31,196,31,52,31,202,31,193,31,193,30,99,31,193,31,67,31,162,31,162,30,100,31,200,31,228,31,101,31,107,31,109,31,109,30,61,31,61,30,116,31,7,31,14,31,212,31,77,31,73,31,73,30,5,31,184,31,184,31,184,30,4,31,94,31,66,31,66,30,199,31,139,31,180,31,75,31,194,31,194,30,248,31,106,31,171,31,43,31,141,31,141,30,141,29,194,31,57,31,78,31,104,31,73,31,241,31,58,31,55,31,218,31,55,31,13,31,37,31,52,31,52,30,230,31,243,31,82,31,11,31,11,30,11,29,171,31,12,31,201,31,38,31,3,31,197,31,176,31,176,30,10,31,10,30,251,31,124,31,64,31,64,30,57,31,70,31,70,30,206,31,162,31,243,31,243,30,72,31,72,30,97,31,20,31,141,31,234,31,88,31,127,31,234,31,248,31,83,31,82,31,40,31,78,31,78,30,24,31,119,31,119,30,2,31,2,30,2,29,237,31,154,31,39,31,39,30,95,31,22,31,47,31,238,31,193,31,75,31,47,31,184,31,98,31,30,31,30,30,136,31,36,31,151,31,15,31,130,31,130,30,130,29,20,31,51,31,110,31,135,31,92,31,92,30,90,31,109,31,109,30,231,31,247,31,80,31,108,31,139,31,12,31,14,31,14,30,33,31,248,31,248,31,57,31,233,31,146,31,146,30,232,31,132,31,199,31,97,31,152,31,10,31,251,31,58,31,167,31,17,31,30,31,201,31,44,31,206,31,194,31,138,31,207,31,216,31,216,30,24,31,103,31,106,31,107,31,78,31,235,31,171,31,18,31,98,31,47,31,2,31,183,31,68,31,39,31,103,31,103,30,128,31,253,31,29,31,208,31,105,31,105,30,105,29,105,28,105,27,173,31,173,30,92,31,210,31,131,31,93,31,189,31,186,31,67,31,144,31,81,31,73,31,73,30,73,29,25,31,88,31,88,30,65,31,89,31,72,31,240,31,240,30,34,31,177,31,224,31,92,31,92,30,123,31,159,31,239,31,178,31,95,31,95,30,152,31,204,31,96,31,28,31,28,30,28,29,223,31,72,31,53,31,53,30,53,29,31,31,244,31,244,30,121,31,63,31,47,31,26,31,26,30,236,31,241,31,180,31,96,31,66,31,66,30,113,31,236,31,190,31,190,30,224,31,105,31,114,31,14,31,9,31,234,31,236,31,86,31,86,30,217,31,217,31,179,31,84,31,65,31,239,31,94,31,237,31,177,31,97,31,235,31,200,31,60,31,240,31,18,31,240,31,181,31,143,31,111,31,103,31,162,31,164,31,172,31,172,30,22,31,245,31,248,31,248,30,100,31,53,31,53,30,96,31,129,31,111,31,205,31,15,31,64,31,233,31,67,31,115,31,115,30,130,31,16,31,155,31,127,31,193,31,4,31,41,31,61,31,231,31,231,30,46,31,4,31,241,31,116,31,183,31,183,30,183,29,191,31,254,31,189,31,51,31,214,31,240,31,127,31,244,31,102,31,152,31,142,31,142,30,58,31,211,31,211,30,218,31,218,30,218,29,218,28,218,27,202,31,15,31,251,31,251,30,94,31,28,31,146,31,137,31,94,31,146,31,146,30,107,31,255,31,214,31,120,31,234,31,117,31,181,31,125,31,94,31,94,30,101,31,114,31,137,31,137,30,72,31,72,30,168,31,240,31,142,31,142,30,22,31,6,31,98,31,98,30,67,31,104,31,42,31,93,31,93,30,212,31,212,30,231,31,4,31,133,31,148,31,40,31,172,31,126,31,197,31,241,31,241,30,80,31,80,30,145,31,157,31,114,31,155,31,43,31,43,30,43,29,133,31,177,31,237,31,171,31,171,30,243,31,73,31,209,31,14,31,124,31,56,31,142,31,65,31,19,31,165,31,11,31,11,30,119,31,220,31,111,31,195,31,113,31,113,30,113,29,76,31,45,31,195,31,254,31,69,31,144,31,47,31,225,31,159,31,16,31,241,31,224,31,58,31,193,31,95,31,92,31,181,31,153,31,124,31,181,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
