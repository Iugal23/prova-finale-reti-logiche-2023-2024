-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 196;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (130,0,159,0,28,0,188,0,14,0,175,0,13,0,0,0,56,0,29,0,131,0,242,0,160,0,26,0,143,0,0,0,0,0,103,0,211,0,159,0,86,0,41,0,54,0,128,0,231,0,0,0,233,0,240,0,43,0,240,0,22,0,45,0,101,0,228,0,141,0,0,0,242,0,186,0,0,0,43,0,132,0,62,0,48,0,206,0,152,0,82,0,0,0,184,0,113,0,97,0,80,0,0,0,237,0,152,0,150,0,128,0,0,0,178,0,95,0,0,0,142,0,0,0,0,0,154,0,8,0,25,0,198,0,0,0,71,0,149,0,0,0,174,0,0,0,74,0,0,0,133,0,214,0,254,0,127,0,76,0,12,0,104,0,66,0,131,0,213,0,33,0,170,0,249,0,0,0,0,0,181,0,148,0,181,0,219,0,116,0,135,0,41,0,0,0,148,0,134,0,0,0,187,0,179,0,27,0,248,0,9,0,0,0,0,0,116,0,28,0,135,0,15,0,79,0,0,0,178,0,227,0,34,0,186,0,231,0,89,0,148,0,199,0,166,0,0,0,27,0,145,0,1,0,191,0,0,0,6,0,64,0,42,0,16,0,201,0,109,0,150,0,218,0,86,0,24,0,179,0,215,0,0,0,218,0,234,0,156,0,0,0,185,0,152,0,224,0,0,0,0,0,105,0,64,0,0,0,182,0,196,0,0,0,41,0,213,0,68,0,70,0,165,0,129,0,0,0,219,0,0,0,74,0,255,0,0,0,21,0,70,0,158,0,0,0,0,0,39,0,191,0,0,0,26,0,252,0,95,0,65,0,34,0,5,0,8,0,145,0,248,0,0,0,38,0,93,0,146,0,186,0,0,0,115,0,108,0,0,0,194,0);
signal scenario_full  : scenario_type := (130,31,159,31,28,31,188,31,14,31,175,31,13,31,13,30,56,31,29,31,131,31,242,31,160,31,26,31,143,31,143,30,143,29,103,31,211,31,159,31,86,31,41,31,54,31,128,31,231,31,231,30,233,31,240,31,43,31,240,31,22,31,45,31,101,31,228,31,141,31,141,30,242,31,186,31,186,30,43,31,132,31,62,31,48,31,206,31,152,31,82,31,82,30,184,31,113,31,97,31,80,31,80,30,237,31,152,31,150,31,128,31,128,30,178,31,95,31,95,30,142,31,142,30,142,29,154,31,8,31,25,31,198,31,198,30,71,31,149,31,149,30,174,31,174,30,74,31,74,30,133,31,214,31,254,31,127,31,76,31,12,31,104,31,66,31,131,31,213,31,33,31,170,31,249,31,249,30,249,29,181,31,148,31,181,31,219,31,116,31,135,31,41,31,41,30,148,31,134,31,134,30,187,31,179,31,27,31,248,31,9,31,9,30,9,29,116,31,28,31,135,31,15,31,79,31,79,30,178,31,227,31,34,31,186,31,231,31,89,31,148,31,199,31,166,31,166,30,27,31,145,31,1,31,191,31,191,30,6,31,64,31,42,31,16,31,201,31,109,31,150,31,218,31,86,31,24,31,179,31,215,31,215,30,218,31,234,31,156,31,156,30,185,31,152,31,224,31,224,30,224,29,105,31,64,31,64,30,182,31,196,31,196,30,41,31,213,31,68,31,70,31,165,31,129,31,129,30,219,31,219,30,74,31,255,31,255,30,21,31,70,31,158,31,158,30,158,29,39,31,191,31,191,30,26,31,252,31,95,31,65,31,34,31,5,31,8,31,145,31,248,31,248,30,38,31,93,31,146,31,186,31,186,30,115,31,108,31,108,30,194,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
