-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_324 is
end project_tb_324;

architecture project_tb_arch_324 of project_tb_324 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 311;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,88,0,0,0,0,0,196,0,87,0,0,0,0,0,32,0,194,0,0,0,0,0,83,0,0,0,229,0,148,0,39,0,196,0,79,0,129,0,138,0,168,0,155,0,149,0,172,0,177,0,211,0,201,0,157,0,240,0,28,0,248,0,111,0,103,0,44,0,147,0,236,0,1,0,0,0,180,0,0,0,156,0,0,0,44,0,0,0,38,0,4,0,111,0,187,0,0,0,75,0,116,0,205,0,0,0,181,0,245,0,87,0,219,0,217,0,0,0,175,0,146,0,44,0,165,0,40,0,111,0,0,0,0,0,207,0,213,0,145,0,71,0,241,0,220,0,0,0,2,0,0,0,92,0,37,0,0,0,78,0,88,0,216,0,0,0,0,0,0,0,69,0,108,0,100,0,150,0,0,0,61,0,0,0,143,0,0,0,88,0,0,0,194,0,186,0,45,0,212,0,141,0,0,0,13,0,0,0,0,0,117,0,134,0,238,0,0,0,183,0,43,0,0,0,0,0,108,0,100,0,140,0,231,0,29,0,42,0,0,0,1,0,59,0,46,0,235,0,0,0,56,0,117,0,0,0,187,0,119,0,133,0,192,0,199,0,141,0,0,0,210,0,117,0,51,0,79,0,132,0,143,0,96,0,57,0,0,0,51,0,133,0,156,0,184,0,0,0,95,0,73,0,98,0,243,0,249,0,170,0,116,0,60,0,55,0,211,0,208,0,108,0,68,0,255,0,108,0,169,0,213,0,15,0,45,0,75,0,178,0,19,0,147,0,0,0,64,0,168,0,212,0,97,0,219,0,0,0,103,0,185,0,204,0,156,0,147,0,166,0,41,0,183,0,0,0,109,0,50,0,180,0,235,0,0,0,0,0,2,0,0,0,185,0,201,0,0,0,63,0,232,0,246,0,122,0,42,0,148,0,16,0,161,0,103,0,0,0,255,0,213,0,144,0,36,0,76,0,38,0,203,0,126,0,21,0,105,0,96,0,241,0,48,0,0,0,157,0,226,0,195,0,150,0,245,0,0,0,0,0,0,0,0,0,219,0,249,0,99,0,0,0,215,0,38,0,71,0,91,0,117,0,152,0,175,0,175,0,22,0,250,0,110,0,140,0,0,0,203,0,0,0,58,0,207,0,167,0,171,0,177,0,189,0,227,0,198,0,208,0,119,0,219,0,0,0,245,0,104,0,232,0,0,0,51,0,0,0,213,0,185,0,0,0,0,0,242,0,227,0,191,0,183,0,142,0,82,0,63,0,111,0,92,0,0,0,5,0,245,0,0,0,125,0,33,0,154,0,0,0,247,0,0,0,90,0,0,0,53,0,76,0,5,0,156,0,233,0,39,0,91,0,4,0,23,0,42,0,218,0,78,0,161,0,108,0,31,0,17,0);
signal scenario_full  : scenario_type := (0,0,88,31,88,30,88,29,196,31,87,31,87,30,87,29,32,31,194,31,194,30,194,29,83,31,83,30,229,31,148,31,39,31,196,31,79,31,129,31,138,31,168,31,155,31,149,31,172,31,177,31,211,31,201,31,157,31,240,31,28,31,248,31,111,31,103,31,44,31,147,31,236,31,1,31,1,30,180,31,180,30,156,31,156,30,44,31,44,30,38,31,4,31,111,31,187,31,187,30,75,31,116,31,205,31,205,30,181,31,245,31,87,31,219,31,217,31,217,30,175,31,146,31,44,31,165,31,40,31,111,31,111,30,111,29,207,31,213,31,145,31,71,31,241,31,220,31,220,30,2,31,2,30,92,31,37,31,37,30,78,31,88,31,216,31,216,30,216,29,216,28,69,31,108,31,100,31,150,31,150,30,61,31,61,30,143,31,143,30,88,31,88,30,194,31,186,31,45,31,212,31,141,31,141,30,13,31,13,30,13,29,117,31,134,31,238,31,238,30,183,31,43,31,43,30,43,29,108,31,100,31,140,31,231,31,29,31,42,31,42,30,1,31,59,31,46,31,235,31,235,30,56,31,117,31,117,30,187,31,119,31,133,31,192,31,199,31,141,31,141,30,210,31,117,31,51,31,79,31,132,31,143,31,96,31,57,31,57,30,51,31,133,31,156,31,184,31,184,30,95,31,73,31,98,31,243,31,249,31,170,31,116,31,60,31,55,31,211,31,208,31,108,31,68,31,255,31,108,31,169,31,213,31,15,31,45,31,75,31,178,31,19,31,147,31,147,30,64,31,168,31,212,31,97,31,219,31,219,30,103,31,185,31,204,31,156,31,147,31,166,31,41,31,183,31,183,30,109,31,50,31,180,31,235,31,235,30,235,29,2,31,2,30,185,31,201,31,201,30,63,31,232,31,246,31,122,31,42,31,148,31,16,31,161,31,103,31,103,30,255,31,213,31,144,31,36,31,76,31,38,31,203,31,126,31,21,31,105,31,96,31,241,31,48,31,48,30,157,31,226,31,195,31,150,31,245,31,245,30,245,29,245,28,245,27,219,31,249,31,99,31,99,30,215,31,38,31,71,31,91,31,117,31,152,31,175,31,175,31,22,31,250,31,110,31,140,31,140,30,203,31,203,30,58,31,207,31,167,31,171,31,177,31,189,31,227,31,198,31,208,31,119,31,219,31,219,30,245,31,104,31,232,31,232,30,51,31,51,30,213,31,185,31,185,30,185,29,242,31,227,31,191,31,183,31,142,31,82,31,63,31,111,31,92,31,92,30,5,31,245,31,245,30,125,31,33,31,154,31,154,30,247,31,247,30,90,31,90,30,53,31,76,31,5,31,156,31,233,31,39,31,91,31,4,31,23,31,42,31,218,31,78,31,161,31,108,31,31,31,17,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
