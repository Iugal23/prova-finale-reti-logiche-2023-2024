-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 800;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (60,0,241,0,196,0,202,0,238,0,215,0,0,0,54,0,100,0,148,0,4,0,0,0,0,0,145,0,0,0,77,0,151,0,185,0,63,0,20,0,222,0,176,0,244,0,236,0,60,0,21,0,90,0,49,0,0,0,0,0,56,0,91,0,0,0,217,0,199,0,130,0,0,0,205,0,0,0,95,0,188,0,76,0,51,0,54,0,184,0,0,0,44,0,155,0,65,0,75,0,69,0,142,0,122,0,95,0,154,0,0,0,87,0,5,0,121,0,132,0,17,0,193,0,171,0,0,0,218,0,131,0,96,0,15,0,23,0,199,0,70,0,184,0,0,0,222,0,41,0,0,0,0,0,22,0,65,0,103,0,81,0,71,0,244,0,50,0,105,0,0,0,171,0,59,0,0,0,10,0,0,0,183,0,158,0,219,0,174,0,142,0,2,0,0,0,0,0,155,0,188,0,99,0,0,0,149,0,250,0,0,0,110,0,0,0,0,0,0,0,9,0,198,0,155,0,0,0,108,0,169,0,199,0,159,0,72,0,38,0,76,0,212,0,147,0,18,0,114,0,52,0,167,0,56,0,225,0,87,0,157,0,155,0,203,0,137,0,104,0,147,0,196,0,156,0,173,0,103,0,136,0,174,0,177,0,51,0,86,0,89,0,97,0,114,0,161,0,152,0,0,0,200,0,113,0,0,0,99,0,81,0,0,0,203,0,255,0,206,0,186,0,162,0,0,0,54,0,137,0,0,0,51,0,156,0,229,0,169,0,86,0,144,0,0,0,203,0,153,0,0,0,46,0,205,0,153,0,115,0,97,0,0,0,193,0,239,0,161,0,0,0,150,0,0,0,14,0,0,0,135,0,32,0,63,0,93,0,143,0,178,0,3,0,45,0,199,0,0,0,0,0,85,0,191,0,64,0,160,0,180,0,29,0,120,0,82,0,180,0,131,0,156,0,109,0,64,0,47,0,0,0,90,0,153,0,194,0,91,0,2,0,119,0,2,0,236,0,210,0,237,0,0,0,0,0,0,0,144,0,241,0,73,0,231,0,219,0,164,0,118,0,68,0,0,0,102,0,171,0,0,0,137,0,197,0,34,0,0,0,18,0,48,0,0,0,0,0,65,0,90,0,56,0,0,0,241,0,152,0,153,0,0,0,132,0,224,0,142,0,92,0,37,0,111,0,129,0,19,0,240,0,230,0,127,0,199,0,47,0,26,0,162,0,0,0,87,0,50,0,199,0,46,0,43,0,177,0,0,0,99,0,173,0,0,0,23,0,0,0,0,0,65,0,35,0,169,0,0,0,177,0,168,0,185,0,0,0,8,0,243,0,0,0,0,0,16,0,34,0,39,0,20,0,202,0,24,0,210,0,101,0,156,0,14,0,148,0,168,0,40,0,204,0,10,0,235,0,131,0,240,0,0,0,32,0,0,0,207,0,80,0,0,0,96,0,225,0,92,0,140,0,95,0,53,0,115,0,54,0,207,0,153,0,226,0,175,0,197,0,179,0,0,0,199,0,0,0,0,0,0,0,0,0,124,0,8,0,0,0,0,0,58,0,104,0,103,0,217,0,0,0,103,0,211,0,191,0,239,0,108,0,0,0,0,0,15,0,193,0,95,0,0,0,0,0,90,0,196,0,243,0,190,0,0,0,172,0,0,0,4,0,130,0,89,0,99,0,194,0,164,0,241,0,20,0,194,0,186,0,142,0,105,0,99,0,91,0,65,0,235,0,118,0,9,0,219,0,127,0,237,0,2,0,0,0,0,0,37,0,127,0,0,0,0,0,171,0,244,0,0,0,168,0,0,0,146,0,222,0,89,0,47,0,67,0,43,0,52,0,0,0,130,0,0,0,0,0,144,0,0,0,13,0,31,0,162,0,89,0,230,0,0,0,209,0,212,0,0,0,49,0,0,0,247,0,0,0,0,0,6,0,58,0,115,0,98,0,121,0,23,0,161,0,210,0,18,0,222,0,0,0,19,0,236,0,151,0,12,0,173,0,0,0,208,0,7,0,98,0,130,0,211,0,112,0,198,0,148,0,0,0,155,0,178,0,215,0,197,0,235,0,146,0,0,0,0,0,0,0,60,0,0,0,0,0,0,0,217,0,211,0,0,0,1,0,0,0,102,0,4,0,243,0,57,0,227,0,109,0,0,0,108,0,79,0,0,0,124,0,94,0,75,0,180,0,31,0,132,0,185,0,255,0,58,0,10,0,224,0,140,0,160,0,235,0,96,0,165,0,204,0,153,0,196,0,0,0,0,0,113,0,0,0,96,0,85,0,136,0,42,0,191,0,91,0,21,0,141,0,150,0,97,0,97,0,128,0,88,0,250,0,214,0,42,0,192,0,0,0,94,0,82,0,175,0,87,0,18,0,199,0,69,0,82,0,241,0,166,0,170,0,73,0,64,0,0,0,46,0,94,0,239,0,119,0,0,0,187,0,15,0,225,0,90,0,156,0,120,0,150,0,2,0,61,0,39,0,210,0,47,0,165,0,158,0,64,0,85,0,64,0,0,0,124,0,0,0,85,0,65,0,209,0,0,0,0,0,167,0,245,0,129,0,229,0,110,0,0,0,157,0,219,0,0,0,247,0,66,0,246,0,210,0,173,0,0,0,19,0,218,0,254,0,123,0,235,0,26,0,192,0,227,0,246,0,126,0,127,0,0,0,0,0,187,0,74,0,252,0,233,0,154,0,134,0,110,0,229,0,217,0,255,0,96,0,180,0,206,0,16,0,202,0,65,0,177,0,6,0,154,0,211,0,0,0,100,0,195,0,0,0,157,0,0,0,0,0,176,0,92,0,0,0,145,0,94,0,0,0,124,0,223,0,58,0,164,0,253,0,217,0,152,0,0,0,143,0,138,0,164,0,243,0,110,0,222,0,0,0,204,0,114,0,67,0,60,0,236,0,115,0,0,0,31,0,49,0,63,0,248,0,7,0,0,0,251,0,153,0,131,0,177,0,51,0,0,0,94,0,0,0,90,0,194,0,71,0,77,0,248,0,108,0,224,0,137,0,253,0,96,0,4,0,0,0,215,0,213,0,46,0,25,0,198,0,0,0,245,0,200,0,102,0,160,0,110,0,199,0,120,0,0,0,112,0,214,0,225,0,93,0,239,0,95,0,227,0,208,0,0,0,28,0,96,0,121,0,152,0,0,0,0,0,13,0,0,0,150,0,33,0,160,0,104,0,0,0,156,0,64,0,63,0,120,0,0,0,3,0,2,0,153,0,115,0,181,0,220,0,144,0,4,0,162,0,0,0,0,0,127,0,207,0,0,0,120,0,0,0,109,0,58,0,85,0,189,0,209,0,214,0,0,0,120,0,2,0,76,0,49,0,150,0,114,0,0,0,1,0,15,0,132,0,104,0,0,0,180,0,178,0,219,0,0,0,223,0,221,0,131,0,24,0,0,0,0,0,11,0,0,0,0,0,37,0,173,0,202,0,165,0,0,0,156,0,47,0,0,0,0,0,250,0,228,0,234,0,109,0,9,0,226,0,0,0,197,0,26,0,151,0,0,0,91,0,0,0,200,0,58,0,227,0,0,0,255,0,88,0,80,0,201,0,189,0,17,0,239,0);
signal scenario_full  : scenario_type := (60,31,241,31,196,31,202,31,238,31,215,31,215,30,54,31,100,31,148,31,4,31,4,30,4,29,145,31,145,30,77,31,151,31,185,31,63,31,20,31,222,31,176,31,244,31,236,31,60,31,21,31,90,31,49,31,49,30,49,29,56,31,91,31,91,30,217,31,199,31,130,31,130,30,205,31,205,30,95,31,188,31,76,31,51,31,54,31,184,31,184,30,44,31,155,31,65,31,75,31,69,31,142,31,122,31,95,31,154,31,154,30,87,31,5,31,121,31,132,31,17,31,193,31,171,31,171,30,218,31,131,31,96,31,15,31,23,31,199,31,70,31,184,31,184,30,222,31,41,31,41,30,41,29,22,31,65,31,103,31,81,31,71,31,244,31,50,31,105,31,105,30,171,31,59,31,59,30,10,31,10,30,183,31,158,31,219,31,174,31,142,31,2,31,2,30,2,29,155,31,188,31,99,31,99,30,149,31,250,31,250,30,110,31,110,30,110,29,110,28,9,31,198,31,155,31,155,30,108,31,169,31,199,31,159,31,72,31,38,31,76,31,212,31,147,31,18,31,114,31,52,31,167,31,56,31,225,31,87,31,157,31,155,31,203,31,137,31,104,31,147,31,196,31,156,31,173,31,103,31,136,31,174,31,177,31,51,31,86,31,89,31,97,31,114,31,161,31,152,31,152,30,200,31,113,31,113,30,99,31,81,31,81,30,203,31,255,31,206,31,186,31,162,31,162,30,54,31,137,31,137,30,51,31,156,31,229,31,169,31,86,31,144,31,144,30,203,31,153,31,153,30,46,31,205,31,153,31,115,31,97,31,97,30,193,31,239,31,161,31,161,30,150,31,150,30,14,31,14,30,135,31,32,31,63,31,93,31,143,31,178,31,3,31,45,31,199,31,199,30,199,29,85,31,191,31,64,31,160,31,180,31,29,31,120,31,82,31,180,31,131,31,156,31,109,31,64,31,47,31,47,30,90,31,153,31,194,31,91,31,2,31,119,31,2,31,236,31,210,31,237,31,237,30,237,29,237,28,144,31,241,31,73,31,231,31,219,31,164,31,118,31,68,31,68,30,102,31,171,31,171,30,137,31,197,31,34,31,34,30,18,31,48,31,48,30,48,29,65,31,90,31,56,31,56,30,241,31,152,31,153,31,153,30,132,31,224,31,142,31,92,31,37,31,111,31,129,31,19,31,240,31,230,31,127,31,199,31,47,31,26,31,162,31,162,30,87,31,50,31,199,31,46,31,43,31,177,31,177,30,99,31,173,31,173,30,23,31,23,30,23,29,65,31,35,31,169,31,169,30,177,31,168,31,185,31,185,30,8,31,243,31,243,30,243,29,16,31,34,31,39,31,20,31,202,31,24,31,210,31,101,31,156,31,14,31,148,31,168,31,40,31,204,31,10,31,235,31,131,31,240,31,240,30,32,31,32,30,207,31,80,31,80,30,96,31,225,31,92,31,140,31,95,31,53,31,115,31,54,31,207,31,153,31,226,31,175,31,197,31,179,31,179,30,199,31,199,30,199,29,199,28,199,27,124,31,8,31,8,30,8,29,58,31,104,31,103,31,217,31,217,30,103,31,211,31,191,31,239,31,108,31,108,30,108,29,15,31,193,31,95,31,95,30,95,29,90,31,196,31,243,31,190,31,190,30,172,31,172,30,4,31,130,31,89,31,99,31,194,31,164,31,241,31,20,31,194,31,186,31,142,31,105,31,99,31,91,31,65,31,235,31,118,31,9,31,219,31,127,31,237,31,2,31,2,30,2,29,37,31,127,31,127,30,127,29,171,31,244,31,244,30,168,31,168,30,146,31,222,31,89,31,47,31,67,31,43,31,52,31,52,30,130,31,130,30,130,29,144,31,144,30,13,31,31,31,162,31,89,31,230,31,230,30,209,31,212,31,212,30,49,31,49,30,247,31,247,30,247,29,6,31,58,31,115,31,98,31,121,31,23,31,161,31,210,31,18,31,222,31,222,30,19,31,236,31,151,31,12,31,173,31,173,30,208,31,7,31,98,31,130,31,211,31,112,31,198,31,148,31,148,30,155,31,178,31,215,31,197,31,235,31,146,31,146,30,146,29,146,28,60,31,60,30,60,29,60,28,217,31,211,31,211,30,1,31,1,30,102,31,4,31,243,31,57,31,227,31,109,31,109,30,108,31,79,31,79,30,124,31,94,31,75,31,180,31,31,31,132,31,185,31,255,31,58,31,10,31,224,31,140,31,160,31,235,31,96,31,165,31,204,31,153,31,196,31,196,30,196,29,113,31,113,30,96,31,85,31,136,31,42,31,191,31,91,31,21,31,141,31,150,31,97,31,97,31,128,31,88,31,250,31,214,31,42,31,192,31,192,30,94,31,82,31,175,31,87,31,18,31,199,31,69,31,82,31,241,31,166,31,170,31,73,31,64,31,64,30,46,31,94,31,239,31,119,31,119,30,187,31,15,31,225,31,90,31,156,31,120,31,150,31,2,31,61,31,39,31,210,31,47,31,165,31,158,31,64,31,85,31,64,31,64,30,124,31,124,30,85,31,65,31,209,31,209,30,209,29,167,31,245,31,129,31,229,31,110,31,110,30,157,31,219,31,219,30,247,31,66,31,246,31,210,31,173,31,173,30,19,31,218,31,254,31,123,31,235,31,26,31,192,31,227,31,246,31,126,31,127,31,127,30,127,29,187,31,74,31,252,31,233,31,154,31,134,31,110,31,229,31,217,31,255,31,96,31,180,31,206,31,16,31,202,31,65,31,177,31,6,31,154,31,211,31,211,30,100,31,195,31,195,30,157,31,157,30,157,29,176,31,92,31,92,30,145,31,94,31,94,30,124,31,223,31,58,31,164,31,253,31,217,31,152,31,152,30,143,31,138,31,164,31,243,31,110,31,222,31,222,30,204,31,114,31,67,31,60,31,236,31,115,31,115,30,31,31,49,31,63,31,248,31,7,31,7,30,251,31,153,31,131,31,177,31,51,31,51,30,94,31,94,30,90,31,194,31,71,31,77,31,248,31,108,31,224,31,137,31,253,31,96,31,4,31,4,30,215,31,213,31,46,31,25,31,198,31,198,30,245,31,200,31,102,31,160,31,110,31,199,31,120,31,120,30,112,31,214,31,225,31,93,31,239,31,95,31,227,31,208,31,208,30,28,31,96,31,121,31,152,31,152,30,152,29,13,31,13,30,150,31,33,31,160,31,104,31,104,30,156,31,64,31,63,31,120,31,120,30,3,31,2,31,153,31,115,31,181,31,220,31,144,31,4,31,162,31,162,30,162,29,127,31,207,31,207,30,120,31,120,30,109,31,58,31,85,31,189,31,209,31,214,31,214,30,120,31,2,31,76,31,49,31,150,31,114,31,114,30,1,31,15,31,132,31,104,31,104,30,180,31,178,31,219,31,219,30,223,31,221,31,131,31,24,31,24,30,24,29,11,31,11,30,11,29,37,31,173,31,202,31,165,31,165,30,156,31,47,31,47,30,47,29,250,31,228,31,234,31,109,31,9,31,226,31,226,30,197,31,26,31,151,31,151,30,91,31,91,30,200,31,58,31,227,31,227,30,255,31,88,31,80,31,201,31,189,31,17,31,239,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
