-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 575;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (91,0,106,0,31,0,173,0,0,0,0,0,165,0,29,0,166,0,121,0,0,0,60,0,204,0,180,0,166,0,50,0,202,0,233,0,109,0,197,0,177,0,0,0,70,0,58,0,0,0,225,0,226,0,0,0,110,0,209,0,252,0,75,0,29,0,168,0,177,0,234,0,165,0,227,0,19,0,156,0,191,0,24,0,244,0,177,0,22,0,51,0,0,0,38,0,99,0,172,0,0,0,134,0,0,0,40,0,69,0,13,0,189,0,184,0,189,0,17,0,0,0,197,0,20,0,0,0,0,0,245,0,177,0,106,0,189,0,127,0,115,0,153,0,104,0,1,0,0,0,0,0,102,0,77,0,66,0,143,0,59,0,213,0,116,0,0,0,42,0,207,0,0,0,73,0,0,0,133,0,0,0,94,0,17,0,232,0,191,0,228,0,10,0,161,0,8,0,0,0,102,0,36,0,142,0,0,0,250,0,236,0,25,0,225,0,133,0,201,0,222,0,246,0,123,0,0,0,243,0,105,0,0,0,33,0,237,0,0,0,6,0,95,0,39,0,87,0,126,0,212,0,64,0,0,0,0,0,243,0,119,0,209,0,89,0,0,0,229,0,77,0,212,0,147,0,80,0,101,0,116,0,185,0,14,0,252,0,235,0,223,0,65,0,155,0,83,0,0,0,157,0,232,0,16,0,0,0,124,0,45,0,14,0,83,0,179,0,130,0,0,0,26,0,111,0,22,0,254,0,149,0,110,0,182,0,22,0,0,0,208,0,197,0,81,0,198,0,231,0,214,0,130,0,237,0,165,0,229,0,203,0,221,0,72,0,246,0,203,0,0,0,208,0,204,0,0,0,0,0,5,0,177,0,114,0,194,0,0,0,67,0,225,0,0,0,98,0,94,0,56,0,83,0,133,0,0,0,11,0,190,0,92,0,5,0,0,0,86,0,36,0,89,0,67,0,75,0,8,0,159,0,30,0,0,0,94,0,217,0,240,0,191,0,0,0,64,0,33,0,6,0,74,0,0,0,0,0,136,0,119,0,220,0,0,0,6,0,143,0,92,0,206,0,32,0,95,0,0,0,4,0,122,0,255,0,83,0,119,0,148,0,35,0,91,0,0,0,78,0,174,0,0,0,0,0,82,0,239,0,26,0,4,0,220,0,29,0,31,0,148,0,31,0,106,0,66,0,208,0,67,0,31,0,34,0,227,0,109,0,210,0,0,0,0,0,154,0,0,0,112,0,191,0,0,0,94,0,37,0,193,0,147,0,0,0,139,0,164,0,177,0,0,0,250,0,121,0,0,0,23,0,40,0,172,0,193,0,223,0,196,0,254,0,71,0,250,0,161,0,4,0,0,0,96,0,135,0,252,0,47,0,101,0,165,0,23,0,245,0,0,0,0,0,92,0,167,0,200,0,0,0,15,0,42,0,161,0,40,0,104,0,222,0,0,0,92,0,99,0,57,0,83,0,0,0,193,0,154,0,0,0,196,0,179,0,0,0,245,0,0,0,204,0,135,0,64,0,141,0,207,0,0,0,206,0,102,0,57,0,253,0,28,0,39,0,20,0,216,0,74,0,255,0,0,0,199,0,176,0,20,0,150,0,157,0,156,0,77,0,0,0,207,0,108,0,251,0,50,0,221,0,58,0,171,0,0,0,233,0,178,0,57,0,60,0,84,0,39,0,11,0,67,0,192,0,197,0,175,0,134,0,140,0,49,0,94,0,120,0,70,0,122,0,0,0,75,0,44,0,247,0,148,0,189,0,115,0,46,0,0,0,115,0,152,0,65,0,44,0,188,0,66,0,88,0,162,0,106,0,0,0,254,0,0,0,205,0,31,0,0,0,248,0,129,0,204,0,211,0,0,0,39,0,140,0,203,0,131,0,79,0,14,0,10,0,63,0,132,0,220,0,32,0,165,0,228,0,80,0,0,0,82,0,190,0,0,0,220,0,0,0,136,0,77,0,51,0,234,0,0,0,30,0,80,0,0,0,85,0,221,0,64,0,15,0,166,0,62,0,222,0,145,0,129,0,244,0,88,0,194,0,0,0,118,0,0,0,0,0,0,0,35,0,0,0,231,0,178,0,203,0,83,0,11,0,100,0,31,0,40,0,235,0,144,0,0,0,75,0,0,0,55,0,27,0,235,0,7,0,64,0,0,0,117,0,152,0,127,0,0,0,176,0,246,0,52,0,225,0,176,0,0,0,0,0,79,0,0,0,89,0,0,0,182,0,185,0,0,0,106,0,122,0,190,0,150,0,13,0,0,0,79,0,104,0,40,0,153,0,135,0,193,0,87,0,117,0,0,0,162,0,0,0,188,0,242,0,165,0,0,0,110,0,78,0,48,0,72,0,205,0,0,0,47,0,172,0,192,0,0,0,0,0,167,0,80,0,54,0,229,0,205,0,202,0,78,0,190,0,211,0,129,0,0,0,22,0,92,0,174,0,190,0,116,0,3,0,35,0,176,0,9,0,32,0,0,0,69,0,115,0,100,0,238,0,0,0,0,0,46,0,14,0,0,0,252,0,208,0,202,0,77,0,0,0,89,0,54,0,210,0,76,0,171,0,223,0,102,0);
signal scenario_full  : scenario_type := (91,31,106,31,31,31,173,31,173,30,173,29,165,31,29,31,166,31,121,31,121,30,60,31,204,31,180,31,166,31,50,31,202,31,233,31,109,31,197,31,177,31,177,30,70,31,58,31,58,30,225,31,226,31,226,30,110,31,209,31,252,31,75,31,29,31,168,31,177,31,234,31,165,31,227,31,19,31,156,31,191,31,24,31,244,31,177,31,22,31,51,31,51,30,38,31,99,31,172,31,172,30,134,31,134,30,40,31,69,31,13,31,189,31,184,31,189,31,17,31,17,30,197,31,20,31,20,30,20,29,245,31,177,31,106,31,189,31,127,31,115,31,153,31,104,31,1,31,1,30,1,29,102,31,77,31,66,31,143,31,59,31,213,31,116,31,116,30,42,31,207,31,207,30,73,31,73,30,133,31,133,30,94,31,17,31,232,31,191,31,228,31,10,31,161,31,8,31,8,30,102,31,36,31,142,31,142,30,250,31,236,31,25,31,225,31,133,31,201,31,222,31,246,31,123,31,123,30,243,31,105,31,105,30,33,31,237,31,237,30,6,31,95,31,39,31,87,31,126,31,212,31,64,31,64,30,64,29,243,31,119,31,209,31,89,31,89,30,229,31,77,31,212,31,147,31,80,31,101,31,116,31,185,31,14,31,252,31,235,31,223,31,65,31,155,31,83,31,83,30,157,31,232,31,16,31,16,30,124,31,45,31,14,31,83,31,179,31,130,31,130,30,26,31,111,31,22,31,254,31,149,31,110,31,182,31,22,31,22,30,208,31,197,31,81,31,198,31,231,31,214,31,130,31,237,31,165,31,229,31,203,31,221,31,72,31,246,31,203,31,203,30,208,31,204,31,204,30,204,29,5,31,177,31,114,31,194,31,194,30,67,31,225,31,225,30,98,31,94,31,56,31,83,31,133,31,133,30,11,31,190,31,92,31,5,31,5,30,86,31,36,31,89,31,67,31,75,31,8,31,159,31,30,31,30,30,94,31,217,31,240,31,191,31,191,30,64,31,33,31,6,31,74,31,74,30,74,29,136,31,119,31,220,31,220,30,6,31,143,31,92,31,206,31,32,31,95,31,95,30,4,31,122,31,255,31,83,31,119,31,148,31,35,31,91,31,91,30,78,31,174,31,174,30,174,29,82,31,239,31,26,31,4,31,220,31,29,31,31,31,148,31,31,31,106,31,66,31,208,31,67,31,31,31,34,31,227,31,109,31,210,31,210,30,210,29,154,31,154,30,112,31,191,31,191,30,94,31,37,31,193,31,147,31,147,30,139,31,164,31,177,31,177,30,250,31,121,31,121,30,23,31,40,31,172,31,193,31,223,31,196,31,254,31,71,31,250,31,161,31,4,31,4,30,96,31,135,31,252,31,47,31,101,31,165,31,23,31,245,31,245,30,245,29,92,31,167,31,200,31,200,30,15,31,42,31,161,31,40,31,104,31,222,31,222,30,92,31,99,31,57,31,83,31,83,30,193,31,154,31,154,30,196,31,179,31,179,30,245,31,245,30,204,31,135,31,64,31,141,31,207,31,207,30,206,31,102,31,57,31,253,31,28,31,39,31,20,31,216,31,74,31,255,31,255,30,199,31,176,31,20,31,150,31,157,31,156,31,77,31,77,30,207,31,108,31,251,31,50,31,221,31,58,31,171,31,171,30,233,31,178,31,57,31,60,31,84,31,39,31,11,31,67,31,192,31,197,31,175,31,134,31,140,31,49,31,94,31,120,31,70,31,122,31,122,30,75,31,44,31,247,31,148,31,189,31,115,31,46,31,46,30,115,31,152,31,65,31,44,31,188,31,66,31,88,31,162,31,106,31,106,30,254,31,254,30,205,31,31,31,31,30,248,31,129,31,204,31,211,31,211,30,39,31,140,31,203,31,131,31,79,31,14,31,10,31,63,31,132,31,220,31,32,31,165,31,228,31,80,31,80,30,82,31,190,31,190,30,220,31,220,30,136,31,77,31,51,31,234,31,234,30,30,31,80,31,80,30,85,31,221,31,64,31,15,31,166,31,62,31,222,31,145,31,129,31,244,31,88,31,194,31,194,30,118,31,118,30,118,29,118,28,35,31,35,30,231,31,178,31,203,31,83,31,11,31,100,31,31,31,40,31,235,31,144,31,144,30,75,31,75,30,55,31,27,31,235,31,7,31,64,31,64,30,117,31,152,31,127,31,127,30,176,31,246,31,52,31,225,31,176,31,176,30,176,29,79,31,79,30,89,31,89,30,182,31,185,31,185,30,106,31,122,31,190,31,150,31,13,31,13,30,79,31,104,31,40,31,153,31,135,31,193,31,87,31,117,31,117,30,162,31,162,30,188,31,242,31,165,31,165,30,110,31,78,31,48,31,72,31,205,31,205,30,47,31,172,31,192,31,192,30,192,29,167,31,80,31,54,31,229,31,205,31,202,31,78,31,190,31,211,31,129,31,129,30,22,31,92,31,174,31,190,31,116,31,3,31,35,31,176,31,9,31,32,31,32,30,69,31,115,31,100,31,238,31,238,30,238,29,46,31,14,31,14,30,252,31,208,31,202,31,77,31,77,30,89,31,54,31,210,31,76,31,171,31,223,31,102,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
