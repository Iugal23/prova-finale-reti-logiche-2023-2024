-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 387;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (133,0,45,0,18,0,0,0,241,0,22,0,17,0,146,0,6,0,183,0,202,0,168,0,58,0,69,0,0,0,0,0,66,0,0,0,0,0,209,0,13,0,0,0,43,0,117,0,36,0,38,0,163,0,92,0,69,0,0,0,0,0,99,0,10,0,0,0,167,0,196,0,136,0,6,0,228,0,50,0,0,0,0,0,251,0,0,0,74,0,229,0,59,0,79,0,180,0,153,0,109,0,255,0,91,0,0,0,6,0,142,0,0,0,204,0,0,0,0,0,28,0,0,0,253,0,0,0,171,0,107,0,0,0,16,0,218,0,80,0,7,0,146,0,0,0,246,0,234,0,108,0,105,0,100,0,54,0,24,0,89,0,189,0,137,0,247,0,67,0,101,0,0,0,243,0,18,0,66,0,0,0,0,0,178,0,177,0,0,0,47,0,147,0,0,0,175,0,0,0,96,0,0,0,174,0,0,0,200,0,114,0,79,0,20,0,252,0,134,0,89,0,72,0,0,0,84,0,83,0,131,0,0,0,136,0,0,0,245,0,66,0,160,0,139,0,165,0,52,0,179,0,0,0,103,0,206,0,255,0,248,0,244,0,0,0,0,0,0,0,212,0,0,0,121,0,28,0,215,0,159,0,176,0,97,0,216,0,226,0,116,0,203,0,27,0,238,0,87,0,0,0,174,0,233,0,236,0,6,0,0,0,0,0,66,0,19,0,137,0,153,0,0,0,33,0,68,0,25,0,101,0,215,0,204,0,0,0,115,0,0,0,0,0,205,0,80,0,229,0,0,0,175,0,0,0,184,0,95,0,0,0,0,0,65,0,0,0,0,0,35,0,188,0,252,0,75,0,84,0,205,0,33,0,140,0,246,0,35,0,32,0,179,0,107,0,203,0,137,0,108,0,7,0,0,0,64,0,162,0,229,0,77,0,253,0,0,0,0,0,182,0,177,0,135,0,36,0,119,0,0,0,0,0,86,0,0,0,216,0,192,0,123,0,146,0,249,0,0,0,92,0,137,0,77,0,69,0,154,0,12,0,0,0,235,0,130,0,41,0,173,0,125,0,56,0,179,0,18,0,0,0,126,0,246,0,79,0,122,0,79,0,104,0,34,0,0,0,150,0,2,0,69,0,94,0,151,0,0,0,170,0,207,0,113,0,159,0,222,0,137,0,6,0,12,0,115,0,126,0,32,0,74,0,187,0,156,0,205,0,133,0,125,0,185,0,92,0,199,0,0,0,8,0,12,0,0,0,12,0,56,0,201,0,0,0,122,0,0,0,139,0,0,0,0,0,173,0,0,0,117,0,0,0,193,0,86,0,78,0,195,0,186,0,66,0,142,0,4,0,107,0,0,0,0,0,0,0,38,0,0,0,49,0,173,0,41,0,0,0,106,0,8,0,15,0,241,0,220,0,61,0,152,0,28,0,45,0,86,0,53,0,205,0,8,0,190,0,227,0,121,0,0,0,0,0,255,0,53,0,0,0,11,0,208,0,109,0,0,0,0,0,80,0,110,0,104,0,92,0,117,0,0,0,0,0,201,0,0,0,209,0,9,0,244,0,0,0,161,0,221,0,0,0,144,0,0,0,212,0,0,0,178,0,179,0,192,0,82,0,68,0,154,0,0,0,148,0,214,0,38,0,140,0,193,0,221,0,0,0,195,0,141,0,250,0,224,0,197,0,43,0,100,0,0,0,200,0,136,0,18,0,0,0,145,0,0,0,48,0,19,0,167,0);
signal scenario_full  : scenario_type := (133,31,45,31,18,31,18,30,241,31,22,31,17,31,146,31,6,31,183,31,202,31,168,31,58,31,69,31,69,30,69,29,66,31,66,30,66,29,209,31,13,31,13,30,43,31,117,31,36,31,38,31,163,31,92,31,69,31,69,30,69,29,99,31,10,31,10,30,167,31,196,31,136,31,6,31,228,31,50,31,50,30,50,29,251,31,251,30,74,31,229,31,59,31,79,31,180,31,153,31,109,31,255,31,91,31,91,30,6,31,142,31,142,30,204,31,204,30,204,29,28,31,28,30,253,31,253,30,171,31,107,31,107,30,16,31,218,31,80,31,7,31,146,31,146,30,246,31,234,31,108,31,105,31,100,31,54,31,24,31,89,31,189,31,137,31,247,31,67,31,101,31,101,30,243,31,18,31,66,31,66,30,66,29,178,31,177,31,177,30,47,31,147,31,147,30,175,31,175,30,96,31,96,30,174,31,174,30,200,31,114,31,79,31,20,31,252,31,134,31,89,31,72,31,72,30,84,31,83,31,131,31,131,30,136,31,136,30,245,31,66,31,160,31,139,31,165,31,52,31,179,31,179,30,103,31,206,31,255,31,248,31,244,31,244,30,244,29,244,28,212,31,212,30,121,31,28,31,215,31,159,31,176,31,97,31,216,31,226,31,116,31,203,31,27,31,238,31,87,31,87,30,174,31,233,31,236,31,6,31,6,30,6,29,66,31,19,31,137,31,153,31,153,30,33,31,68,31,25,31,101,31,215,31,204,31,204,30,115,31,115,30,115,29,205,31,80,31,229,31,229,30,175,31,175,30,184,31,95,31,95,30,95,29,65,31,65,30,65,29,35,31,188,31,252,31,75,31,84,31,205,31,33,31,140,31,246,31,35,31,32,31,179,31,107,31,203,31,137,31,108,31,7,31,7,30,64,31,162,31,229,31,77,31,253,31,253,30,253,29,182,31,177,31,135,31,36,31,119,31,119,30,119,29,86,31,86,30,216,31,192,31,123,31,146,31,249,31,249,30,92,31,137,31,77,31,69,31,154,31,12,31,12,30,235,31,130,31,41,31,173,31,125,31,56,31,179,31,18,31,18,30,126,31,246,31,79,31,122,31,79,31,104,31,34,31,34,30,150,31,2,31,69,31,94,31,151,31,151,30,170,31,207,31,113,31,159,31,222,31,137,31,6,31,12,31,115,31,126,31,32,31,74,31,187,31,156,31,205,31,133,31,125,31,185,31,92,31,199,31,199,30,8,31,12,31,12,30,12,31,56,31,201,31,201,30,122,31,122,30,139,31,139,30,139,29,173,31,173,30,117,31,117,30,193,31,86,31,78,31,195,31,186,31,66,31,142,31,4,31,107,31,107,30,107,29,107,28,38,31,38,30,49,31,173,31,41,31,41,30,106,31,8,31,15,31,241,31,220,31,61,31,152,31,28,31,45,31,86,31,53,31,205,31,8,31,190,31,227,31,121,31,121,30,121,29,255,31,53,31,53,30,11,31,208,31,109,31,109,30,109,29,80,31,110,31,104,31,92,31,117,31,117,30,117,29,201,31,201,30,209,31,9,31,244,31,244,30,161,31,221,31,221,30,144,31,144,30,212,31,212,30,178,31,179,31,192,31,82,31,68,31,154,31,154,30,148,31,214,31,38,31,140,31,193,31,221,31,221,30,195,31,141,31,250,31,224,31,197,31,43,31,100,31,100,30,200,31,136,31,18,31,18,30,145,31,145,30,48,31,19,31,167,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
