-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 769;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (1,0,209,0,100,0,159,0,81,0,0,0,2,0,251,0,39,0,22,0,91,0,0,0,140,0,246,0,99,0,0,0,0,0,167,0,0,0,0,0,224,0,130,0,217,0,7,0,0,0,232,0,221,0,196,0,187,0,58,0,143,0,114,0,19,0,174,0,0,0,0,0,90,0,20,0,74,0,119,0,0,0,162,0,0,0,99,0,0,0,149,0,233,0,89,0,0,0,126,0,0,0,191,0,180,0,236,0,11,0,82,0,105,0,121,0,163,0,44,0,0,0,128,0,0,0,101,0,143,0,107,0,0,0,0,0,0,0,248,0,76,0,253,0,166,0,124,0,0,0,162,0,68,0,247,0,34,0,0,0,168,0,243,0,137,0,224,0,0,0,224,0,0,0,0,0,138,0,38,0,167,0,0,0,0,0,0,0,38,0,242,0,210,0,0,0,179,0,0,0,193,0,136,0,201,0,126,0,193,0,193,0,80,0,54,0,185,0,236,0,71,0,107,0,139,0,0,0,169,0,134,0,250,0,171,0,75,0,0,0,18,0,107,0,0,0,0,0,0,0,124,0,0,0,33,0,0,0,165,0,82,0,0,0,253,0,50,0,152,0,217,0,163,0,80,0,211,0,0,0,39,0,182,0,4,0,82,0,183,0,219,0,114,0,0,0,227,0,0,0,56,0,15,0,224,0,101,0,92,0,142,0,91,0,0,0,0,0,131,0,99,0,202,0,121,0,3,0,0,0,0,0,200,0,0,0,55,0,0,0,114,0,99,0,235,0,29,0,219,0,203,0,116,0,166,0,0,0,201,0,0,0,155,0,44,0,151,0,0,0,134,0,37,0,179,0,14,0,147,0,2,0,0,0,158,0,185,0,70,0,202,0,129,0,189,0,181,0,0,0,0,0,249,0,117,0,146,0,29,0,0,0,56,0,2,0,0,0,172,0,111,0,77,0,27,0,44,0,219,0,79,0,65,0,239,0,64,0,175,0,207,0,70,0,0,0,191,0,149,0,0,0,112,0,209,0,200,0,0,0,234,0,0,0,24,0,7,0,18,0,125,0,0,0,0,0,9,0,162,0,0,0,0,0,203,0,61,0,0,0,95,0,136,0,0,0,0,0,81,0,191,0,206,0,0,0,19,0,31,0,81,0,99,0,113,0,13,0,139,0,238,0,111,0,211,0,0,0,93,0,226,0,241,0,0,0,185,0,156,0,190,0,136,0,47,0,224,0,0,0,66,0,118,0,0,0,150,0,157,0,0,0,238,0,116,0,0,0,245,0,20,0,124,0,11,0,151,0,0,0,0,0,237,0,0,0,0,0,0,0,0,0,141,0,63,0,222,0,129,0,182,0,75,0,15,0,0,0,154,0,91,0,120,0,10,0,0,0,243,0,137,0,190,0,109,0,225,0,14,0,184,0,81,0,75,0,126,0,0,0,104,0,107,0,232,0,128,0,118,0,90,0,0,0,77,0,23,0,0,0,68,0,147,0,47,0,0,0,0,0,4,0,96,0,70,0,150,0,0,0,212,0,52,0,154,0,145,0,192,0,185,0,60,0,71,0,14,0,0,0,145,0,3,0,0,0,0,0,151,0,5,0,253,0,187,0,161,0,0,0,41,0,131,0,28,0,0,0,25,0,0,0,8,0,84,0,0,0,248,0,51,0,8,0,73,0,78,0,0,0,0,0,0,0,197,0,208,0,0,0,0,0,250,0,93,0,125,0,0,0,253,0,172,0,189,0,17,0,173,0,96,0,237,0,171,0,0,0,229,0,156,0,0,0,125,0,250,0,31,0,65,0,118,0,85,0,204,0,202,0,117,0,235,0,219,0,66,0,0,0,206,0,69,0,101,0,75,0,29,0,124,0,0,0,0,0,99,0,58,0,196,0,166,0,0,0,201,0,17,0,206,0,11,0,0,0,226,0,70,0,24,0,16,0,167,0,82,0,98,0,242,0,42,0,0,0,201,0,26,0,199,0,148,0,0,0,147,0,158,0,149,0,172,0,55,0,220,0,0,0,194,0,0,0,168,0,214,0,180,0,0,0,188,0,27,0,60,0,200,0,200,0,91,0,109,0,165,0,186,0,151,0,253,0,20,0,110,0,108,0,78,0,137,0,160,0,95,0,197,0,157,0,0,0,235,0,169,0,245,0,0,0,9,0,190,0,146,0,0,0,0,0,162,0,115,0,0,0,244,0,162,0,105,0,200,0,254,0,202,0,74,0,134,0,0,0,240,0,78,0,0,0,0,0,109,0,242,0,160,0,0,0,166,0,223,0,0,0,227,0,247,0,187,0,243,0,101,0,0,0,0,0,53,0,156,0,0,0,97,0,189,0,116,0,201,0,146,0,0,0,0,0,56,0,160,0,233,0,0,0,143,0,134,0,69,0,0,0,19,0,0,0,0,0,60,0,226,0,117,0,231,0,96,0,173,0,22,0,242,0,0,0,184,0,90,0,96,0,207,0,88,0,0,0,252,0,0,0,228,0,202,0,163,0,191,0,16,0,0,0,204,0,0,0,176,0,235,0,235,0,186,0,185,0,151,0,126,0,254,0,18,0,8,0,69,0,0,0,0,0,97,0,58,0,215,0,227,0,224,0,188,0,0,0,0,0,20,0,66,0,14,0,160,0,111,0,212,0,131,0,201,0,82,0,186,0,26,0,53,0,67,0,154,0,125,0,0,0,129,0,240,0,253,0,62,0,0,0,108,0,0,0,154,0,242,0,163,0,39,0,186,0,90,0,0,0,185,0,252,0,0,0,12,0,146,0,127,0,45,0,137,0,0,0,140,0,234,0,183,0,106,0,14,0,3,0,0,0,204,0,0,0,144,0,35,0,31,0,0,0,169,0,50,0,145,0,99,0,0,0,175,0,0,0,122,0,54,0,227,0,236,0,0,0,185,0,194,0,164,0,250,0,17,0,221,0,0,0,236,0,0,0,0,0,121,0,121,0,54,0,34,0,0,0,252,0,218,0,198,0,109,0,162,0,0,0,182,0,196,0,117,0,224,0,140,0,0,0,236,0,195,0,234,0,119,0,7,0,0,0,195,0,0,0,11,0,0,0,224,0,0,0,168,0,85,0,20,0,39,0,224,0,208,0,77,0,123,0,0,0,185,0,206,0,173,0,110,0,143,0,217,0,170,0,124,0,226,0,0,0,192,0,242,0,222,0,105,0,90,0,159,0,0,0,124,0,253,0,0,0,91,0,95,0,81,0,184,0,194,0,187,0,101,0,74,0,104,0,63,0,55,0,162,0,0,0,188,0,140,0,0,0,238,0,93,0,188,0,70,0,246,0,90,0,167,0,230,0,132,0,242,0,251,0,180,0,161,0,169,0,0,0,91,0,0,0,216,0,20,0,57,0,213,0,0,0,230,0,217,0,225,0,0,0,136,0,65,0,120,0,37,0,102,0,218,0,0,0,186,0,0,0,230,0,157,0,111,0);
signal scenario_full  : scenario_type := (1,31,209,31,100,31,159,31,81,31,81,30,2,31,251,31,39,31,22,31,91,31,91,30,140,31,246,31,99,31,99,30,99,29,167,31,167,30,167,29,224,31,130,31,217,31,7,31,7,30,232,31,221,31,196,31,187,31,58,31,143,31,114,31,19,31,174,31,174,30,174,29,90,31,20,31,74,31,119,31,119,30,162,31,162,30,99,31,99,30,149,31,233,31,89,31,89,30,126,31,126,30,191,31,180,31,236,31,11,31,82,31,105,31,121,31,163,31,44,31,44,30,128,31,128,30,101,31,143,31,107,31,107,30,107,29,107,28,248,31,76,31,253,31,166,31,124,31,124,30,162,31,68,31,247,31,34,31,34,30,168,31,243,31,137,31,224,31,224,30,224,31,224,30,224,29,138,31,38,31,167,31,167,30,167,29,167,28,38,31,242,31,210,31,210,30,179,31,179,30,193,31,136,31,201,31,126,31,193,31,193,31,80,31,54,31,185,31,236,31,71,31,107,31,139,31,139,30,169,31,134,31,250,31,171,31,75,31,75,30,18,31,107,31,107,30,107,29,107,28,124,31,124,30,33,31,33,30,165,31,82,31,82,30,253,31,50,31,152,31,217,31,163,31,80,31,211,31,211,30,39,31,182,31,4,31,82,31,183,31,219,31,114,31,114,30,227,31,227,30,56,31,15,31,224,31,101,31,92,31,142,31,91,31,91,30,91,29,131,31,99,31,202,31,121,31,3,31,3,30,3,29,200,31,200,30,55,31,55,30,114,31,99,31,235,31,29,31,219,31,203,31,116,31,166,31,166,30,201,31,201,30,155,31,44,31,151,31,151,30,134,31,37,31,179,31,14,31,147,31,2,31,2,30,158,31,185,31,70,31,202,31,129,31,189,31,181,31,181,30,181,29,249,31,117,31,146,31,29,31,29,30,56,31,2,31,2,30,172,31,111,31,77,31,27,31,44,31,219,31,79,31,65,31,239,31,64,31,175,31,207,31,70,31,70,30,191,31,149,31,149,30,112,31,209,31,200,31,200,30,234,31,234,30,24,31,7,31,18,31,125,31,125,30,125,29,9,31,162,31,162,30,162,29,203,31,61,31,61,30,95,31,136,31,136,30,136,29,81,31,191,31,206,31,206,30,19,31,31,31,81,31,99,31,113,31,13,31,139,31,238,31,111,31,211,31,211,30,93,31,226,31,241,31,241,30,185,31,156,31,190,31,136,31,47,31,224,31,224,30,66,31,118,31,118,30,150,31,157,31,157,30,238,31,116,31,116,30,245,31,20,31,124,31,11,31,151,31,151,30,151,29,237,31,237,30,237,29,237,28,237,27,141,31,63,31,222,31,129,31,182,31,75,31,15,31,15,30,154,31,91,31,120,31,10,31,10,30,243,31,137,31,190,31,109,31,225,31,14,31,184,31,81,31,75,31,126,31,126,30,104,31,107,31,232,31,128,31,118,31,90,31,90,30,77,31,23,31,23,30,68,31,147,31,47,31,47,30,47,29,4,31,96,31,70,31,150,31,150,30,212,31,52,31,154,31,145,31,192,31,185,31,60,31,71,31,14,31,14,30,145,31,3,31,3,30,3,29,151,31,5,31,253,31,187,31,161,31,161,30,41,31,131,31,28,31,28,30,25,31,25,30,8,31,84,31,84,30,248,31,51,31,8,31,73,31,78,31,78,30,78,29,78,28,197,31,208,31,208,30,208,29,250,31,93,31,125,31,125,30,253,31,172,31,189,31,17,31,173,31,96,31,237,31,171,31,171,30,229,31,156,31,156,30,125,31,250,31,31,31,65,31,118,31,85,31,204,31,202,31,117,31,235,31,219,31,66,31,66,30,206,31,69,31,101,31,75,31,29,31,124,31,124,30,124,29,99,31,58,31,196,31,166,31,166,30,201,31,17,31,206,31,11,31,11,30,226,31,70,31,24,31,16,31,167,31,82,31,98,31,242,31,42,31,42,30,201,31,26,31,199,31,148,31,148,30,147,31,158,31,149,31,172,31,55,31,220,31,220,30,194,31,194,30,168,31,214,31,180,31,180,30,188,31,27,31,60,31,200,31,200,31,91,31,109,31,165,31,186,31,151,31,253,31,20,31,110,31,108,31,78,31,137,31,160,31,95,31,197,31,157,31,157,30,235,31,169,31,245,31,245,30,9,31,190,31,146,31,146,30,146,29,162,31,115,31,115,30,244,31,162,31,105,31,200,31,254,31,202,31,74,31,134,31,134,30,240,31,78,31,78,30,78,29,109,31,242,31,160,31,160,30,166,31,223,31,223,30,227,31,247,31,187,31,243,31,101,31,101,30,101,29,53,31,156,31,156,30,97,31,189,31,116,31,201,31,146,31,146,30,146,29,56,31,160,31,233,31,233,30,143,31,134,31,69,31,69,30,19,31,19,30,19,29,60,31,226,31,117,31,231,31,96,31,173,31,22,31,242,31,242,30,184,31,90,31,96,31,207,31,88,31,88,30,252,31,252,30,228,31,202,31,163,31,191,31,16,31,16,30,204,31,204,30,176,31,235,31,235,31,186,31,185,31,151,31,126,31,254,31,18,31,8,31,69,31,69,30,69,29,97,31,58,31,215,31,227,31,224,31,188,31,188,30,188,29,20,31,66,31,14,31,160,31,111,31,212,31,131,31,201,31,82,31,186,31,26,31,53,31,67,31,154,31,125,31,125,30,129,31,240,31,253,31,62,31,62,30,108,31,108,30,154,31,242,31,163,31,39,31,186,31,90,31,90,30,185,31,252,31,252,30,12,31,146,31,127,31,45,31,137,31,137,30,140,31,234,31,183,31,106,31,14,31,3,31,3,30,204,31,204,30,144,31,35,31,31,31,31,30,169,31,50,31,145,31,99,31,99,30,175,31,175,30,122,31,54,31,227,31,236,31,236,30,185,31,194,31,164,31,250,31,17,31,221,31,221,30,236,31,236,30,236,29,121,31,121,31,54,31,34,31,34,30,252,31,218,31,198,31,109,31,162,31,162,30,182,31,196,31,117,31,224,31,140,31,140,30,236,31,195,31,234,31,119,31,7,31,7,30,195,31,195,30,11,31,11,30,224,31,224,30,168,31,85,31,20,31,39,31,224,31,208,31,77,31,123,31,123,30,185,31,206,31,173,31,110,31,143,31,217,31,170,31,124,31,226,31,226,30,192,31,242,31,222,31,105,31,90,31,159,31,159,30,124,31,253,31,253,30,91,31,95,31,81,31,184,31,194,31,187,31,101,31,74,31,104,31,63,31,55,31,162,31,162,30,188,31,140,31,140,30,238,31,93,31,188,31,70,31,246,31,90,31,167,31,230,31,132,31,242,31,251,31,180,31,161,31,169,31,169,30,91,31,91,30,216,31,20,31,57,31,213,31,213,30,230,31,217,31,225,31,225,30,136,31,65,31,120,31,37,31,102,31,218,31,218,30,186,31,186,30,230,31,157,31,111,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
