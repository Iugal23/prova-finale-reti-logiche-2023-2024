-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 815;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (1,0,81,0,146,0,55,0,107,0,49,0,206,0,29,0,0,0,179,0,79,0,249,0,20,0,159,0,253,0,0,0,0,0,163,0,109,0,138,0,0,0,56,0,153,0,97,0,147,0,105,0,39,0,52,0,74,0,215,0,153,0,234,0,147,0,156,0,96,0,0,0,172,0,123,0,2,0,125,0,248,0,20,0,129,0,0,0,242,0,204,0,54,0,38,0,245,0,77,0,0,0,3,0,195,0,118,0,206,0,73,0,0,0,39,0,174,0,217,0,0,0,92,0,0,0,0,0,251,0,235,0,126,0,92,0,231,0,234,0,40,0,100,0,193,0,117,0,140,0,143,0,145,0,1,0,57,0,237,0,211,0,93,0,152,0,156,0,0,0,152,0,215,0,0,0,0,0,86,0,0,0,74,0,135,0,203,0,194,0,0,0,0,0,244,0,178,0,163,0,184,0,29,0,98,0,109,0,0,0,188,0,38,0,182,0,9,0,129,0,180,0,104,0,0,0,87,0,124,0,0,0,28,0,3,0,56,0,239,0,80,0,104,0,70,0,0,0,167,0,174,0,0,0,0,0,202,0,0,0,215,0,0,0,0,0,128,0,42,0,0,0,51,0,0,0,68,0,240,0,137,0,142,0,129,0,125,0,18,0,66,0,103,0,193,0,20,0,182,0,245,0,0,0,4,0,244,0,202,0,228,0,188,0,216,0,177,0,208,0,36,0,125,0,0,0,95,0,186,0,58,0,10,0,181,0,0,0,50,0,153,0,35,0,47,0,0,0,235,0,248,0,244,0,54,0,122,0,118,0,0,0,7,0,131,0,17,0,243,0,115,0,63,0,128,0,242,0,213,0,1,0,248,0,63,0,110,0,89,0,102,0,91,0,214,0,167,0,0,0,59,0,109,0,111,0,0,0,55,0,155,0,175,0,0,0,232,0,176,0,0,0,56,0,14,0,56,0,225,0,28,0,0,0,244,0,89,0,93,0,218,0,209,0,113,0,109,0,100,0,96,0,237,0,194,0,194,0,174,0,18,0,27,0,63,0,85,0,86,0,128,0,41,0,0,0,0,0,231,0,73,0,0,0,54,0,140,0,193,0,21,0,41,0,182,0,0,0,0,0,0,0,30,0,203,0,0,0,57,0,64,0,0,0,71,0,244,0,123,0,51,0,235,0,131,0,133,0,118,0,165,0,133,0,134,0,141,0,221,0,0,0,240,0,28,0,5,0,211,0,16,0,156,0,202,0,113,0,107,0,58,0,26,0,138,0,201,0,65,0,0,0,209,0,230,0,236,0,90,0,207,0,36,0,82,0,27,0,139,0,231,0,35,0,0,0,21,0,0,0,22,0,133,0,148,0,105,0,133,0,135,0,77,0,180,0,118,0,154,0,145,0,4,0,64,0,208,0,241,0,0,0,252,0,85,0,129,0,116,0,242,0,166,0,0,0,245,0,88,0,176,0,0,0,174,0,224,0,96,0,32,0,170,0,6,0,126,0,199,0,186,0,65,0,0,0,89,0,177,0,154,0,234,0,128,0,66,0,66,0,0,0,48,0,11,0,66,0,17,0,68,0,105,0,124,0,154,0,65,0,33,0,117,0,0,0,110,0,60,0,0,0,0,0,36,0,0,0,205,0,180,0,178,0,29,0,63,0,69,0,122,0,211,0,0,0,0,0,126,0,125,0,209,0,118,0,130,0,19,0,247,0,205,0,0,0,135,0,0,0,66,0,227,0,0,0,203,0,154,0,0,0,0,0,149,0,9,0,122,0,151,0,0,0,117,0,130,0,147,0,190,0,14,0,0,0,10,0,97,0,136,0,0,0,220,0,0,0,223,0,0,0,220,0,220,0,139,0,47,0,89,0,198,0,157,0,0,0,220,0,176,0,175,0,253,0,129,0,219,0,0,0,73,0,0,0,47,0,96,0,95,0,66,0,0,0,135,0,0,0,47,0,166,0,24,0,0,0,81,0,72,0,171,0,199,0,93,0,0,0,92,0,134,0,0,0,142,0,66,0,90,0,192,0,162,0,224,0,244,0,204,0,131,0,177,0,199,0,214,0,108,0,210,0,58,0,196,0,194,0,145,0,0,0,126,0,120,0,35,0,176,0,52,0,173,0,141,0,178,0,87,0,140,0,108,0,154,0,122,0,0,0,189,0,0,0,0,0,0,0,0,0,245,0,198,0,73,0,115,0,253,0,115,0,189,0,128,0,74,0,225,0,11,0,120,0,66,0,208,0,0,0,60,0,184,0,71,0,154,0,36,0,0,0,213,0,237,0,196,0,0,0,170,0,169,0,15,0,185,0,0,0,133,0,0,0,224,0,162,0,0,0,8,0,0,0,243,0,119,0,182,0,0,0,123,0,0,0,46,0,230,0,141,0,22,0,250,0,173,0,212,0,227,0,0,0,185,0,70,0,95,0,29,0,108,0,213,0,35,0,105,0,93,0,207,0,0,0,95,0,250,0,205,0,190,0,212,0,1,0,71,0,0,0,182,0,181,0,166,0,21,0,26,0,142,0,92,0,145,0,0,0,4,0,0,0,0,0,104,0,0,0,65,0,65,0,178,0,224,0,229,0,5,0,10,0,129,0,0,0,0,0,74,0,104,0,232,0,179,0,2,0,119,0,0,0,194,0,1,0,69,0,99,0,162,0,183,0,0,0,114,0,222,0,214,0,225,0,18,0,202,0,157,0,190,0,148,0,22,0,12,0,74,0,131,0,0,0,182,0,0,0,190,0,23,0,218,0,55,0,108,0,222,0,243,0,0,0,226,0,0,0,80,0,0,0,0,0,0,0,0,0,62,0,105,0,39,0,225,0,186,0,83,0,81,0,0,0,0,0,87,0,3,0,0,0,143,0,105,0,107,0,67,0,148,0,68,0,31,0,138,0,163,0,217,0,67,0,49,0,190,0,6,0,139,0,57,0,209,0,172,0,141,0,183,0,142,0,97,0,5,0,0,0,136,0,101,0,163,0,0,0,66,0,0,0,121,0,254,0,0,0,57,0,3,0,121,0,0,0,23,0,0,0,254,0,14,0,67,0,89,0,57,0,118,0,230,0,192,0,34,0,128,0,172,0,227,0,204,0,170,0,204,0,0,0,202,0,112,0,122,0,0,0,195,0,10,0,0,0,188,0,89,0,16,0,114,0,151,0,56,0,4,0,117,0,25,0,0,0,117,0,155,0,245,0,173,0,100,0,0,0,95,0,68,0,234,0,253,0,0,0,0,0,9,0,115,0,217,0,0,0,0,0,86,0,0,0,122,0,0,0,96,0,172,0,182,0,0,0,39,0,116,0,0,0,86,0,89,0,79,0,2,0,0,0,7,0,100,0,97,0,195,0,6,0,2,0,202,0,240,0,0,0,126,0,149,0,41,0,0,0,40,0,215,0,183,0,165,0,0,0,1,0,108,0,101,0,0,0,118,0,0,0,0,0,77,0,92,0,0,0,231,0,178,0,41,0,20,0,69,0,0,0,48,0,63,0,48,0,252,0,0,0,70,0,0,0,149,0,0,0,110,0,71,0,0,0,156,0,30,0,0,0,5,0,0,0,74,0,18,0,133,0,240,0,109,0,98,0,255,0,0,0,80,0,210,0,242,0,193,0,109,0,0,0,0,0,0,0,47,0,79,0,0,0,51,0,148,0);
signal scenario_full  : scenario_type := (1,31,81,31,146,31,55,31,107,31,49,31,206,31,29,31,29,30,179,31,79,31,249,31,20,31,159,31,253,31,253,30,253,29,163,31,109,31,138,31,138,30,56,31,153,31,97,31,147,31,105,31,39,31,52,31,74,31,215,31,153,31,234,31,147,31,156,31,96,31,96,30,172,31,123,31,2,31,125,31,248,31,20,31,129,31,129,30,242,31,204,31,54,31,38,31,245,31,77,31,77,30,3,31,195,31,118,31,206,31,73,31,73,30,39,31,174,31,217,31,217,30,92,31,92,30,92,29,251,31,235,31,126,31,92,31,231,31,234,31,40,31,100,31,193,31,117,31,140,31,143,31,145,31,1,31,57,31,237,31,211,31,93,31,152,31,156,31,156,30,152,31,215,31,215,30,215,29,86,31,86,30,74,31,135,31,203,31,194,31,194,30,194,29,244,31,178,31,163,31,184,31,29,31,98,31,109,31,109,30,188,31,38,31,182,31,9,31,129,31,180,31,104,31,104,30,87,31,124,31,124,30,28,31,3,31,56,31,239,31,80,31,104,31,70,31,70,30,167,31,174,31,174,30,174,29,202,31,202,30,215,31,215,30,215,29,128,31,42,31,42,30,51,31,51,30,68,31,240,31,137,31,142,31,129,31,125,31,18,31,66,31,103,31,193,31,20,31,182,31,245,31,245,30,4,31,244,31,202,31,228,31,188,31,216,31,177,31,208,31,36,31,125,31,125,30,95,31,186,31,58,31,10,31,181,31,181,30,50,31,153,31,35,31,47,31,47,30,235,31,248,31,244,31,54,31,122,31,118,31,118,30,7,31,131,31,17,31,243,31,115,31,63,31,128,31,242,31,213,31,1,31,248,31,63,31,110,31,89,31,102,31,91,31,214,31,167,31,167,30,59,31,109,31,111,31,111,30,55,31,155,31,175,31,175,30,232,31,176,31,176,30,56,31,14,31,56,31,225,31,28,31,28,30,244,31,89,31,93,31,218,31,209,31,113,31,109,31,100,31,96,31,237,31,194,31,194,31,174,31,18,31,27,31,63,31,85,31,86,31,128,31,41,31,41,30,41,29,231,31,73,31,73,30,54,31,140,31,193,31,21,31,41,31,182,31,182,30,182,29,182,28,30,31,203,31,203,30,57,31,64,31,64,30,71,31,244,31,123,31,51,31,235,31,131,31,133,31,118,31,165,31,133,31,134,31,141,31,221,31,221,30,240,31,28,31,5,31,211,31,16,31,156,31,202,31,113,31,107,31,58,31,26,31,138,31,201,31,65,31,65,30,209,31,230,31,236,31,90,31,207,31,36,31,82,31,27,31,139,31,231,31,35,31,35,30,21,31,21,30,22,31,133,31,148,31,105,31,133,31,135,31,77,31,180,31,118,31,154,31,145,31,4,31,64,31,208,31,241,31,241,30,252,31,85,31,129,31,116,31,242,31,166,31,166,30,245,31,88,31,176,31,176,30,174,31,224,31,96,31,32,31,170,31,6,31,126,31,199,31,186,31,65,31,65,30,89,31,177,31,154,31,234,31,128,31,66,31,66,31,66,30,48,31,11,31,66,31,17,31,68,31,105,31,124,31,154,31,65,31,33,31,117,31,117,30,110,31,60,31,60,30,60,29,36,31,36,30,205,31,180,31,178,31,29,31,63,31,69,31,122,31,211,31,211,30,211,29,126,31,125,31,209,31,118,31,130,31,19,31,247,31,205,31,205,30,135,31,135,30,66,31,227,31,227,30,203,31,154,31,154,30,154,29,149,31,9,31,122,31,151,31,151,30,117,31,130,31,147,31,190,31,14,31,14,30,10,31,97,31,136,31,136,30,220,31,220,30,223,31,223,30,220,31,220,31,139,31,47,31,89,31,198,31,157,31,157,30,220,31,176,31,175,31,253,31,129,31,219,31,219,30,73,31,73,30,47,31,96,31,95,31,66,31,66,30,135,31,135,30,47,31,166,31,24,31,24,30,81,31,72,31,171,31,199,31,93,31,93,30,92,31,134,31,134,30,142,31,66,31,90,31,192,31,162,31,224,31,244,31,204,31,131,31,177,31,199,31,214,31,108,31,210,31,58,31,196,31,194,31,145,31,145,30,126,31,120,31,35,31,176,31,52,31,173,31,141,31,178,31,87,31,140,31,108,31,154,31,122,31,122,30,189,31,189,30,189,29,189,28,189,27,245,31,198,31,73,31,115,31,253,31,115,31,189,31,128,31,74,31,225,31,11,31,120,31,66,31,208,31,208,30,60,31,184,31,71,31,154,31,36,31,36,30,213,31,237,31,196,31,196,30,170,31,169,31,15,31,185,31,185,30,133,31,133,30,224,31,162,31,162,30,8,31,8,30,243,31,119,31,182,31,182,30,123,31,123,30,46,31,230,31,141,31,22,31,250,31,173,31,212,31,227,31,227,30,185,31,70,31,95,31,29,31,108,31,213,31,35,31,105,31,93,31,207,31,207,30,95,31,250,31,205,31,190,31,212,31,1,31,71,31,71,30,182,31,181,31,166,31,21,31,26,31,142,31,92,31,145,31,145,30,4,31,4,30,4,29,104,31,104,30,65,31,65,31,178,31,224,31,229,31,5,31,10,31,129,31,129,30,129,29,74,31,104,31,232,31,179,31,2,31,119,31,119,30,194,31,1,31,69,31,99,31,162,31,183,31,183,30,114,31,222,31,214,31,225,31,18,31,202,31,157,31,190,31,148,31,22,31,12,31,74,31,131,31,131,30,182,31,182,30,190,31,23,31,218,31,55,31,108,31,222,31,243,31,243,30,226,31,226,30,80,31,80,30,80,29,80,28,80,27,62,31,105,31,39,31,225,31,186,31,83,31,81,31,81,30,81,29,87,31,3,31,3,30,143,31,105,31,107,31,67,31,148,31,68,31,31,31,138,31,163,31,217,31,67,31,49,31,190,31,6,31,139,31,57,31,209,31,172,31,141,31,183,31,142,31,97,31,5,31,5,30,136,31,101,31,163,31,163,30,66,31,66,30,121,31,254,31,254,30,57,31,3,31,121,31,121,30,23,31,23,30,254,31,14,31,67,31,89,31,57,31,118,31,230,31,192,31,34,31,128,31,172,31,227,31,204,31,170,31,204,31,204,30,202,31,112,31,122,31,122,30,195,31,10,31,10,30,188,31,89,31,16,31,114,31,151,31,56,31,4,31,117,31,25,31,25,30,117,31,155,31,245,31,173,31,100,31,100,30,95,31,68,31,234,31,253,31,253,30,253,29,9,31,115,31,217,31,217,30,217,29,86,31,86,30,122,31,122,30,96,31,172,31,182,31,182,30,39,31,116,31,116,30,86,31,89,31,79,31,2,31,2,30,7,31,100,31,97,31,195,31,6,31,2,31,202,31,240,31,240,30,126,31,149,31,41,31,41,30,40,31,215,31,183,31,165,31,165,30,1,31,108,31,101,31,101,30,118,31,118,30,118,29,77,31,92,31,92,30,231,31,178,31,41,31,20,31,69,31,69,30,48,31,63,31,48,31,252,31,252,30,70,31,70,30,149,31,149,30,110,31,71,31,71,30,156,31,30,31,30,30,5,31,5,30,74,31,18,31,133,31,240,31,109,31,98,31,255,31,255,30,80,31,210,31,242,31,193,31,109,31,109,30,109,29,109,28,47,31,79,31,79,30,51,31,148,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
