-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 869;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (29,0,129,0,108,0,15,0,119,0,249,0,248,0,252,0,109,0,214,0,100,0,158,0,82,0,209,0,186,0,0,0,253,0,25,0,0,0,156,0,182,0,151,0,0,0,83,0,186,0,45,0,187,0,9,0,0,0,156,0,74,0,0,0,35,0,1,0,58,0,135,0,192,0,0,0,237,0,43,0,0,0,93,0,80,0,214,0,76,0,202,0,182,0,201,0,244,0,0,0,10,0,0,0,197,0,0,0,45,0,0,0,80,0,70,0,0,0,16,0,23,0,172,0,82,0,159,0,37,0,107,0,247,0,173,0,207,0,129,0,19,0,75,0,58,0,20,0,196,0,101,0,0,0,178,0,98,0,0,0,93,0,0,0,72,0,203,0,0,0,198,0,0,0,0,0,19,0,0,0,68,0,193,0,60,0,242,0,185,0,3,0,210,0,0,0,13,0,0,0,188,0,226,0,172,0,224,0,135,0,15,0,202,0,126,0,91,0,91,0,0,0,0,0,238,0,51,0,0,0,130,0,55,0,237,0,232,0,40,0,76,0,186,0,109,0,0,0,35,0,206,0,38,0,190,0,240,0,5,0,0,0,0,0,248,0,119,0,0,0,114,0,0,0,0,0,151,0,0,0,156,0,98,0,63,0,247,0,26,0,116,0,27,0,0,0,201,0,245,0,0,0,173,0,0,0,133,0,0,0,84,0,69,0,85,0,237,0,45,0,168,0,124,0,48,0,0,0,132,0,14,0,0,0,5,0,95,0,0,0,34,0,127,0,0,0,133,0,231,0,28,0,68,0,4,0,203,0,26,0,121,0,0,0,244,0,185,0,93,0,19,0,180,0,225,0,172,0,137,0,26,0,0,0,0,0,211,0,0,0,0,0,38,0,2,0,17,0,214,0,35,0,131,0,24,0,97,0,42,0,37,0,160,0,182,0,147,0,151,0,197,0,68,0,35,0,38,0,0,0,0,0,84,0,194,0,0,0,0,0,120,0,0,0,169,0,78,0,0,0,100,0,155,0,47,0,125,0,186,0,190,0,117,0,85,0,214,0,186,0,87,0,169,0,95,0,115,0,194,0,0,0,114,0,167,0,0,0,169,0,182,0,19,0,113,0,167,0,0,0,58,0,211,0,132,0,32,0,0,0,18,0,127,0,178,0,235,0,178,0,167,0,190,0,211,0,205,0,0,0,0,0,0,0,144,0,83,0,0,0,240,0,208,0,0,0,191,0,0,0,79,0,79,0,200,0,0,0,0,0,0,0,148,0,67,0,0,0,114,0,160,0,5,0,160,0,133,0,87,0,230,0,209,0,48,0,110,0,223,0,28,0,21,0,13,0,22,0,130,0,0,0,68,0,185,0,78,0,8,0,94,0,142,0,151,0,16,0,59,0,100,0,17,0,50,0,66,0,0,0,222,0,188,0,0,0,0,0,23,0,134,0,0,0,0,0,31,0,103,0,225,0,123,0,71,0,128,0,142,0,118,0,108,0,96,0,0,0,0,0,0,0,198,0,13,0,190,0,0,0,49,0,4,0,21,0,185,0,237,0,107,0,242,0,248,0,188,0,158,0,0,0,75,0,144,0,134,0,157,0,104,0,0,0,154,0,155,0,27,0,210,0,0,0,8,0,0,0,0,0,34,0,225,0,230,0,86,0,0,0,0,0,66,0,237,0,108,0,214,0,75,0,154,0,0,0,209,0,0,0,244,0,250,0,232,0,185,0,0,0,168,0,0,0,75,0,0,0,214,0,166,0,139,0,97,0,0,0,127,0,150,0,23,0,71,0,185,0,46,0,220,0,107,0,14,0,220,0,96,0,186,0,0,0,87,0,242,0,192,0,158,0,83,0,107,0,0,0,0,0,199,0,217,0,40,0,43,0,66,0,61,0,255,0,79,0,78,0,55,0,101,0,8,0,241,0,148,0,33,0,7,0,13,0,229,0,247,0,97,0,0,0,16,0,21,0,42,0,25,0,96,0,32,0,218,0,59,0,45,0,208,0,159,0,0,0,24,0,66,0,16,0,38,0,193,0,0,0,45,0,0,0,51,0,11,0,3,0,156,0,255,0,159,0,71,0,121,0,0,0,149,0,249,0,200,0,99,0,127,0,0,0,0,0,13,0,167,0,39,0,0,0,0,0,0,0,218,0,0,0,172,0,0,0,227,0,38,0,151,0,0,0,24,0,165,0,81,0,230,0,143,0,119,0,109,0,194,0,173,0,126,0,16,0,77,0,70,0,56,0,96,0,155,0,236,0,0,0,156,0,114,0,174,0,0,0,162,0,0,0,1,0,0,0,232,0,122,0,232,0,252,0,205,0,0,0,226,0,0,0,180,0,145,0,81,0,38,0,118,0,0,0,73,0,0,0,140,0,128,0,239,0,157,0,225,0,218,0,81,0,137,0,0,0,189,0,80,0,48,0,23,0,0,0,179,0,65,0,233,0,137,0,116,0,225,0,0,0,71,0,0,0,166,0,49,0,20,0,80,0,0,0,240,0,12,0,43,0,129,0,132,0,126,0,226,0,0,0,0,0,231,0,0,0,218,0,59,0,19,0,205,0,31,0,80,0,85,0,206,0,63,0,139,0,0,0,114,0,55,0,216,0,223,0,0,0,240,0,107,0,244,0,214,0,249,0,0,0,0,0,90,0,139,0,133,0,232,0,200,0,165,0,152,0,127,0,202,0,0,0,54,0,101,0,20,0,0,0,174,0,192,0,211,0,169,0,0,0,195,0,149,0,0,0,169,0,0,0,0,0,0,0,84,0,21,0,97,0,0,0,176,0,18,0,85,0,27,0,100,0,207,0,165,0,0,0,146,0,190,0,198,0,175,0,44,0,24,0,175,0,0,0,62,0,8,0,232,0,0,0,0,0,154,0,207,0,39,0,210,0,0,0,15,0,191,0,31,0,255,0,0,0,0,0,196,0,0,0,208,0,242,0,0,0,252,0,165,0,67,0,0,0,158,0,145,0,0,0,7,0,106,0,31,0,58,0,220,0,0,0,35,0,0,0,0,0,36,0,0,0,124,0,60,0,122,0,212,0,85,0,148,0,195,0,38,0,0,0,197,0,159,0,173,0,17,0,0,0,99,0,145,0,37,0,170,0,15,0,0,0,0,0,202,0,0,0,213,0,165,0,24,0,121,0,0,0,103,0,202,0,223,0,63,0,245,0,213,0,166,0,199,0,63,0,19,0,10,0,0,0,230,0,0,0,0,0,212,0,151,0,0,0,97,0,0,0,141,0,120,0,0,0,117,0,0,0,0,0,245,0,198,0,57,0,146,0,201,0,15,0,66,0,50,0,53,0,0,0,28,0,207,0,252,0,148,0,0,0,0,0,85,0,0,0,234,0,221,0,200,0,0,0,0,0,32,0,0,0,0,0,21,0,0,0,253,0,163,0,202,0,137,0,27,0,8,0,44,0,214,0,214,0,60,0,181,0,16,0,205,0,0,0,121,0,133,0,160,0,0,0,19,0,234,0,52,0,201,0,214,0,40,0,0,0,185,0,75,0,0,0,145,0,57,0,0,0,212,0,104,0,59,0,97,0,216,0,10,0,47,0,0,0,187,0,146,0,236,0,255,0,202,0,159,0,0,0,151,0,6,0,0,0,0,0,36,0,20,0,125,0,60,0,0,0,205,0,11,0,149,0,64,0,0,0,145,0,40,0,134,0,0,0,93,0,234,0,35,0,0,0,83,0,164,0,162,0,0,0,108,0,115,0,0,0,168,0,0,0,0,0,0,0,236,0,91,0,0,0,232,0,190,0,40,0,209,0,174,0,105,0,0,0,126,0,70,0,29,0,36,0,97,0,231,0,0,0,134,0,2,0,0,0,103,0,0,0,179,0,112,0,245,0,197,0,250,0,45,0,138,0,113,0,153,0,0,0,166,0);
signal scenario_full  : scenario_type := (29,31,129,31,108,31,15,31,119,31,249,31,248,31,252,31,109,31,214,31,100,31,158,31,82,31,209,31,186,31,186,30,253,31,25,31,25,30,156,31,182,31,151,31,151,30,83,31,186,31,45,31,187,31,9,31,9,30,156,31,74,31,74,30,35,31,1,31,58,31,135,31,192,31,192,30,237,31,43,31,43,30,93,31,80,31,214,31,76,31,202,31,182,31,201,31,244,31,244,30,10,31,10,30,197,31,197,30,45,31,45,30,80,31,70,31,70,30,16,31,23,31,172,31,82,31,159,31,37,31,107,31,247,31,173,31,207,31,129,31,19,31,75,31,58,31,20,31,196,31,101,31,101,30,178,31,98,31,98,30,93,31,93,30,72,31,203,31,203,30,198,31,198,30,198,29,19,31,19,30,68,31,193,31,60,31,242,31,185,31,3,31,210,31,210,30,13,31,13,30,188,31,226,31,172,31,224,31,135,31,15,31,202,31,126,31,91,31,91,31,91,30,91,29,238,31,51,31,51,30,130,31,55,31,237,31,232,31,40,31,76,31,186,31,109,31,109,30,35,31,206,31,38,31,190,31,240,31,5,31,5,30,5,29,248,31,119,31,119,30,114,31,114,30,114,29,151,31,151,30,156,31,98,31,63,31,247,31,26,31,116,31,27,31,27,30,201,31,245,31,245,30,173,31,173,30,133,31,133,30,84,31,69,31,85,31,237,31,45,31,168,31,124,31,48,31,48,30,132,31,14,31,14,30,5,31,95,31,95,30,34,31,127,31,127,30,133,31,231,31,28,31,68,31,4,31,203,31,26,31,121,31,121,30,244,31,185,31,93,31,19,31,180,31,225,31,172,31,137,31,26,31,26,30,26,29,211,31,211,30,211,29,38,31,2,31,17,31,214,31,35,31,131,31,24,31,97,31,42,31,37,31,160,31,182,31,147,31,151,31,197,31,68,31,35,31,38,31,38,30,38,29,84,31,194,31,194,30,194,29,120,31,120,30,169,31,78,31,78,30,100,31,155,31,47,31,125,31,186,31,190,31,117,31,85,31,214,31,186,31,87,31,169,31,95,31,115,31,194,31,194,30,114,31,167,31,167,30,169,31,182,31,19,31,113,31,167,31,167,30,58,31,211,31,132,31,32,31,32,30,18,31,127,31,178,31,235,31,178,31,167,31,190,31,211,31,205,31,205,30,205,29,205,28,144,31,83,31,83,30,240,31,208,31,208,30,191,31,191,30,79,31,79,31,200,31,200,30,200,29,200,28,148,31,67,31,67,30,114,31,160,31,5,31,160,31,133,31,87,31,230,31,209,31,48,31,110,31,223,31,28,31,21,31,13,31,22,31,130,31,130,30,68,31,185,31,78,31,8,31,94,31,142,31,151,31,16,31,59,31,100,31,17,31,50,31,66,31,66,30,222,31,188,31,188,30,188,29,23,31,134,31,134,30,134,29,31,31,103,31,225,31,123,31,71,31,128,31,142,31,118,31,108,31,96,31,96,30,96,29,96,28,198,31,13,31,190,31,190,30,49,31,4,31,21,31,185,31,237,31,107,31,242,31,248,31,188,31,158,31,158,30,75,31,144,31,134,31,157,31,104,31,104,30,154,31,155,31,27,31,210,31,210,30,8,31,8,30,8,29,34,31,225,31,230,31,86,31,86,30,86,29,66,31,237,31,108,31,214,31,75,31,154,31,154,30,209,31,209,30,244,31,250,31,232,31,185,31,185,30,168,31,168,30,75,31,75,30,214,31,166,31,139,31,97,31,97,30,127,31,150,31,23,31,71,31,185,31,46,31,220,31,107,31,14,31,220,31,96,31,186,31,186,30,87,31,242,31,192,31,158,31,83,31,107,31,107,30,107,29,199,31,217,31,40,31,43,31,66,31,61,31,255,31,79,31,78,31,55,31,101,31,8,31,241,31,148,31,33,31,7,31,13,31,229,31,247,31,97,31,97,30,16,31,21,31,42,31,25,31,96,31,32,31,218,31,59,31,45,31,208,31,159,31,159,30,24,31,66,31,16,31,38,31,193,31,193,30,45,31,45,30,51,31,11,31,3,31,156,31,255,31,159,31,71,31,121,31,121,30,149,31,249,31,200,31,99,31,127,31,127,30,127,29,13,31,167,31,39,31,39,30,39,29,39,28,218,31,218,30,172,31,172,30,227,31,38,31,151,31,151,30,24,31,165,31,81,31,230,31,143,31,119,31,109,31,194,31,173,31,126,31,16,31,77,31,70,31,56,31,96,31,155,31,236,31,236,30,156,31,114,31,174,31,174,30,162,31,162,30,1,31,1,30,232,31,122,31,232,31,252,31,205,31,205,30,226,31,226,30,180,31,145,31,81,31,38,31,118,31,118,30,73,31,73,30,140,31,128,31,239,31,157,31,225,31,218,31,81,31,137,31,137,30,189,31,80,31,48,31,23,31,23,30,179,31,65,31,233,31,137,31,116,31,225,31,225,30,71,31,71,30,166,31,49,31,20,31,80,31,80,30,240,31,12,31,43,31,129,31,132,31,126,31,226,31,226,30,226,29,231,31,231,30,218,31,59,31,19,31,205,31,31,31,80,31,85,31,206,31,63,31,139,31,139,30,114,31,55,31,216,31,223,31,223,30,240,31,107,31,244,31,214,31,249,31,249,30,249,29,90,31,139,31,133,31,232,31,200,31,165,31,152,31,127,31,202,31,202,30,54,31,101,31,20,31,20,30,174,31,192,31,211,31,169,31,169,30,195,31,149,31,149,30,169,31,169,30,169,29,169,28,84,31,21,31,97,31,97,30,176,31,18,31,85,31,27,31,100,31,207,31,165,31,165,30,146,31,190,31,198,31,175,31,44,31,24,31,175,31,175,30,62,31,8,31,232,31,232,30,232,29,154,31,207,31,39,31,210,31,210,30,15,31,191,31,31,31,255,31,255,30,255,29,196,31,196,30,208,31,242,31,242,30,252,31,165,31,67,31,67,30,158,31,145,31,145,30,7,31,106,31,31,31,58,31,220,31,220,30,35,31,35,30,35,29,36,31,36,30,124,31,60,31,122,31,212,31,85,31,148,31,195,31,38,31,38,30,197,31,159,31,173,31,17,31,17,30,99,31,145,31,37,31,170,31,15,31,15,30,15,29,202,31,202,30,213,31,165,31,24,31,121,31,121,30,103,31,202,31,223,31,63,31,245,31,213,31,166,31,199,31,63,31,19,31,10,31,10,30,230,31,230,30,230,29,212,31,151,31,151,30,97,31,97,30,141,31,120,31,120,30,117,31,117,30,117,29,245,31,198,31,57,31,146,31,201,31,15,31,66,31,50,31,53,31,53,30,28,31,207,31,252,31,148,31,148,30,148,29,85,31,85,30,234,31,221,31,200,31,200,30,200,29,32,31,32,30,32,29,21,31,21,30,253,31,163,31,202,31,137,31,27,31,8,31,44,31,214,31,214,31,60,31,181,31,16,31,205,31,205,30,121,31,133,31,160,31,160,30,19,31,234,31,52,31,201,31,214,31,40,31,40,30,185,31,75,31,75,30,145,31,57,31,57,30,212,31,104,31,59,31,97,31,216,31,10,31,47,31,47,30,187,31,146,31,236,31,255,31,202,31,159,31,159,30,151,31,6,31,6,30,6,29,36,31,20,31,125,31,60,31,60,30,205,31,11,31,149,31,64,31,64,30,145,31,40,31,134,31,134,30,93,31,234,31,35,31,35,30,83,31,164,31,162,31,162,30,108,31,115,31,115,30,168,31,168,30,168,29,168,28,236,31,91,31,91,30,232,31,190,31,40,31,209,31,174,31,105,31,105,30,126,31,70,31,29,31,36,31,97,31,231,31,231,30,134,31,2,31,2,30,103,31,103,30,179,31,112,31,245,31,197,31,250,31,45,31,138,31,113,31,153,31,153,30,166,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
