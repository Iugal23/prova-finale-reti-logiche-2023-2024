-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_674 is
end project_tb_674;

architecture project_tb_arch_674 of project_tb_674 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 240;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,26,0,136,0,42,0,40,0,58,0,73,0,233,0,99,0,3,0,0,0,32,0,216,0,127,0,117,0,231,0,54,0,132,0,25,0,194,0,192,0,141,0,181,0,94,0,227,0,76,0,0,0,169,0,69,0,87,0,0,0,181,0,2,0,89,0,64,0,0,0,218,0,119,0,78,0,45,0,0,0,22,0,111,0,103,0,69,0,0,0,49,0,0,0,230,0,126,0,10,0,191,0,231,0,166,0,177,0,117,0,0,0,32,0,0,0,220,0,252,0,0,0,197,0,42,0,191,0,0,0,239,0,182,0,35,0,144,0,232,0,214,0,136,0,0,0,171,0,0,0,201,0,76,0,122,0,176,0,128,0,34,0,44,0,209,0,0,0,140,0,90,0,27,0,162,0,0,0,19,0,84,0,51,0,80,0,0,0,166,0,59,0,90,0,38,0,0,0,0,0,175,0,0,0,137,0,120,0,172,0,153,0,2,0,240,0,131,0,90,0,136,0,187,0,19,0,182,0,246,0,65,0,193,0,105,0,166,0,187,0,0,0,254,0,0,0,115,0,233,0,218,0,250,0,159,0,151,0,79,0,0,0,167,0,251,0,87,0,0,0,233,0,146,0,51,0,241,0,226,0,128,0,61,0,115,0,241,0,233,0,0,0,79,0,0,0,0,0,91,0,181,0,239,0,125,0,194,0,164,0,0,0,232,0,194,0,0,0,221,0,28,0,139,0,231,0,136,0,0,0,0,0,0,0,150,0,176,0,92,0,0,0,189,0,22,0,0,0,243,0,152,0,70,0,219,0,1,0,73,0,215,0,0,0,0,0,112,0,0,0,48,0,91,0,0,0,225,0,205,0,69,0,101,0,49,0,90,0,77,0,61,0,154,0,115,0,233,0,19,0,241,0,222,0,0,0,0,0,200,0,102,0,72,0,181,0,93,0,40,0,81,0,0,0,249,0,41,0,0,0,173,0,53,0,9,0,222,0,115,0,42,0,27,0,18,0,154,0,219,0,0,0,167,0,177,0,107,0,44,0,0,0,8,0,34,0,0,0,107,0,183,0,0,0,17,0,20,0);
signal scenario_full  : scenario_type := (0,0,26,31,136,31,42,31,40,31,58,31,73,31,233,31,99,31,3,31,3,30,32,31,216,31,127,31,117,31,231,31,54,31,132,31,25,31,194,31,192,31,141,31,181,31,94,31,227,31,76,31,76,30,169,31,69,31,87,31,87,30,181,31,2,31,89,31,64,31,64,30,218,31,119,31,78,31,45,31,45,30,22,31,111,31,103,31,69,31,69,30,49,31,49,30,230,31,126,31,10,31,191,31,231,31,166,31,177,31,117,31,117,30,32,31,32,30,220,31,252,31,252,30,197,31,42,31,191,31,191,30,239,31,182,31,35,31,144,31,232,31,214,31,136,31,136,30,171,31,171,30,201,31,76,31,122,31,176,31,128,31,34,31,44,31,209,31,209,30,140,31,90,31,27,31,162,31,162,30,19,31,84,31,51,31,80,31,80,30,166,31,59,31,90,31,38,31,38,30,38,29,175,31,175,30,137,31,120,31,172,31,153,31,2,31,240,31,131,31,90,31,136,31,187,31,19,31,182,31,246,31,65,31,193,31,105,31,166,31,187,31,187,30,254,31,254,30,115,31,233,31,218,31,250,31,159,31,151,31,79,31,79,30,167,31,251,31,87,31,87,30,233,31,146,31,51,31,241,31,226,31,128,31,61,31,115,31,241,31,233,31,233,30,79,31,79,30,79,29,91,31,181,31,239,31,125,31,194,31,164,31,164,30,232,31,194,31,194,30,221,31,28,31,139,31,231,31,136,31,136,30,136,29,136,28,150,31,176,31,92,31,92,30,189,31,22,31,22,30,243,31,152,31,70,31,219,31,1,31,73,31,215,31,215,30,215,29,112,31,112,30,48,31,91,31,91,30,225,31,205,31,69,31,101,31,49,31,90,31,77,31,61,31,154,31,115,31,233,31,19,31,241,31,222,31,222,30,222,29,200,31,102,31,72,31,181,31,93,31,40,31,81,31,81,30,249,31,41,31,41,30,173,31,53,31,9,31,222,31,115,31,42,31,27,31,18,31,154,31,219,31,219,30,167,31,177,31,107,31,44,31,44,30,8,31,34,31,34,30,107,31,183,31,183,30,17,31,20,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
