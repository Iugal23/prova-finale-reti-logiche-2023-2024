-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_179 is
end project_tb_179;

architecture project_tb_arch_179 of project_tb_179 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1011;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (22,0,234,0,0,0,0,0,0,0,44,0,43,0,50,0,7,0,79,0,20,0,108,0,0,0,248,0,161,0,146,0,0,0,0,0,40,0,170,0,16,0,59,0,25,0,82,0,237,0,172,0,6,0,93,0,218,0,0,0,5,0,0,0,18,0,87,0,254,0,4,0,174,0,134,0,164,0,0,0,252,0,70,0,190,0,195,0,18,0,63,0,77,0,170,0,0,0,51,0,140,0,163,0,114,0,0,0,67,0,0,0,78,0,162,0,206,0,46,0,148,0,11,0,174,0,78,0,228,0,150,0,117,0,65,0,151,0,63,0,90,0,119,0,86,0,149,0,40,0,255,0,0,0,201,0,0,0,206,0,105,0,78,0,35,0,83,0,186,0,24,0,5,0,217,0,51,0,52,0,57,0,0,0,208,0,94,0,55,0,0,0,201,0,185,0,0,0,241,0,250,0,182,0,142,0,57,0,0,0,159,0,149,0,232,0,0,0,191,0,144,0,67,0,0,0,0,0,131,0,0,0,79,0,0,0,126,0,160,0,57,0,209,0,169,0,28,0,161,0,38,0,167,0,179,0,163,0,67,0,55,0,149,0,73,0,23,0,143,0,0,0,255,0,235,0,98,0,241,0,26,0,189,0,72,0,0,0,0,0,0,0,0,0,128,0,121,0,108,0,49,0,0,0,191,0,246,0,103,0,0,0,118,0,0,0,151,0,137,0,9,0,0,0,176,0,162,0,210,0,0,0,138,0,0,0,160,0,0,0,245,0,169,0,35,0,23,0,211,0,0,0,118,0,234,0,192,0,0,0,0,0,0,0,169,0,122,0,154,0,0,0,166,0,0,0,33,0,190,0,131,0,164,0,0,0,83,0,137,0,203,0,108,0,209,0,222,0,207,0,106,0,0,0,206,0,41,0,245,0,56,0,0,0,1,0,200,0,227,0,165,0,209,0,209,0,55,0,0,0,4,0,55,0,172,0,35,0,81,0,0,0,0,0,91,0,24,0,208,0,0,0,193,0,85,0,0,0,156,0,41,0,167,0,18,0,0,0,45,0,0,0,41,0,85,0,0,0,190,0,213,0,223,0,152,0,99,0,223,0,3,0,9,0,110,0,238,0,236,0,190,0,26,0,163,0,228,0,32,0,2,0,71,0,48,0,103,0,171,0,0,0,241,0,234,0,48,0,116,0,147,0,0,0,0,0,211,0,156,0,144,0,236,0,56,0,175,0,106,0,0,0,32,0,134,0,147,0,198,0,0,0,108,0,208,0,17,0,0,0,207,0,189,0,99,0,147,0,94,0,68,0,132,0,0,0,238,0,0,0,55,0,198,0,77,0,237,0,0,0,0,0,225,0,181,0,223,0,239,0,214,0,235,0,154,0,39,0,222,0,255,0,0,0,132,0,20,0,92,0,0,0,11,0,0,0,110,0,91,0,189,0,162,0,14,0,0,0,0,0,94,0,159,0,221,0,179,0,113,0,0,0,0,0,0,0,25,0,182,0,104,0,34,0,71,0,209,0,138,0,0,0,14,0,107,0,220,0,165,0,0,0,42,0,158,0,17,0,14,0,123,0,165,0,169,0,78,0,0,0,207,0,188,0,171,0,9,0,3,0,21,0,159,0,0,0,155,0,155,0,221,0,150,0,0,0,44,0,0,0,213,0,181,0,111,0,0,0,0,0,194,0,0,0,24,0,0,0,38,0,194,0,0,0,134,0,202,0,232,0,0,0,234,0,138,0,120,0,16,0,218,0,148,0,106,0,92,0,0,0,163,0,0,0,201,0,47,0,0,0,187,0,79,0,18,0,57,0,0,0,235,0,156,0,27,0,241,0,207,0,105,0,52,0,0,0,174,0,123,0,16,0,23,0,151,0,0,0,0,0,253,0,11,0,0,0,231,0,0,0,0,0,95,0,0,0,108,0,58,0,0,0,166,0,47,0,87,0,41,0,194,0,0,0,0,0,75,0,139,0,242,0,0,0,37,0,167,0,8,0,231,0,79,0,242,0,144,0,0,0,43,0,0,0,44,0,153,0,48,0,127,0,200,0,0,0,94,0,0,0,0,0,113,0,206,0,230,0,172,0,0,0,0,0,0,0,145,0,0,0,219,0,64,0,103,0,0,0,196,0,124,0,55,0,247,0,55,0,142,0,0,0,188,0,0,0,246,0,96,0,10,0,56,0,0,0,125,0,3,0,149,0,209,0,231,0,167,0,226,0,168,0,234,0,92,0,159,0,22,0,38,0,193,0,0,0,220,0,235,0,213,0,68,0,165,0,165,0,242,0,3,0,253,0,137,0,28,0,0,0,0,0,0,0,202,0,171,0,249,0,121,0,214,0,242,0,0,0,0,0,126,0,212,0,135,0,153,0,145,0,45,0,0,0,62,0,8,0,199,0,239,0,239,0,115,0,37,0,226,0,179,0,224,0,171,0,96,0,28,0,0,0,245,0,209,0,245,0,182,0,196,0,111,0,0,0,30,0,0,0,95,0,239,0,0,0,202,0,50,0,151,0,3,0,73,0,155,0,0,0,8,0,12,0,53,0,185,0,56,0,54,0,5,0,171,0,53,0,196,0,121,0,50,0,0,0,83,0,148,0,232,0,199,0,162,0,253,0,32,0,67,0,195,0,104,0,221,0,0,0,219,0,221,0,222,0,186,0,67,0,102,0,204,0,75,0,198,0,230,0,0,0,70,0,135,0,0,0,91,0,230,0,110,0,148,0,0,0,0,0,242,0,0,0,144,0,0,0,0,0,231,0,132,0,214,0,102,0,116,0,205,0,23,0,253,0,169,0,156,0,233,0,0,0,216,0,56,0,213,0,242,0,0,0,209,0,167,0,237,0,151,0,0,0,186,0,119,0,33,0,0,0,99,0,0,0,220,0,121,0,139,0,55,0,81,0,240,0,255,0,64,0,242,0,253,0,211,0,11,0,204,0,231,0,81,0,64,0,52,0,0,0,120,0,199,0,158,0,120,0,0,0,242,0,53,0,123,0,61,0,181,0,55,0,74,0,71,0,79,0,95,0,56,0,4,0,26,0,123,0,100,0,218,0,174,0,178,0,88,0,243,0,0,0,0,0,186,0,184,0,247,0,108,0,11,0,105,0,249,0,0,0,129,0,23,0,155,0,83,0,0,0,0,0,34,0,162,0,248,0,220,0,230,0,244,0,158,0,178,0,74,0,142,0,140,0,93,0,189,0,203,0,146,0,238,0,31,0,187,0,249,0,118,0,76,0,202,0,165,0,0,0,0,0,243,0,255,0,135,0,128,0,0,0,2,0,134,0,195,0,126,0,65,0,62,0,137,0,209,0,39,0,0,0,28,0,0,0,99,0,222,0,254,0,0,0,66,0,69,0,125,0,8,0,154,0,178,0,220,0,253,0,189,0,206,0,253,0,0,0,29,0,194,0,93,0,54,0,0,0,15,0,211,0,243,0,71,0,126,0,0,0,137,0,185,0,241,0,0,0,26,0,155,0,100,0,0,0,118,0,0,0,81,0,154,0,0,0,137,0,207,0,192,0,236,0,218,0,0,0,241,0,103,0,46,0,211,0,0,0,222,0,195,0,33,0,172,0,0,0,182,0,181,0,62,0,139,0,62,0,169,0,0,0,119,0,209,0,0,0,228,0,23,0,0,0,30,0,56,0,251,0,0,0,157,0,48,0,25,0,120,0,51,0,82,0,0,0,161,0,250,0,49,0,180,0,196,0,225,0,0,0,83,0,108,0,160,0,221,0,15,0,165,0,61,0,59,0,61,0,178,0,0,0,0,0,0,0,101,0,81,0,0,0,39,0,247,0,216,0,229,0,133,0,211,0,105,0,0,0,80,0,23,0,0,0,179,0,0,0,26,0,138,0,143,0,81,0,178,0,119,0,182,0,116,0,0,0,0,0,250,0,0,0,0,0,88,0,0,0,187,0,90,0,16,0,81,0,184,0,190,0,171,0,0,0,250,0,253,0,35,0,115,0,108,0,122,0,86,0,170,0,216,0,13,0,150,0,188,0,17,0,49,0,11,0,27,0,139,0,25,0,0,0,153,0,105,0,0,0,0,0,15,0,170,0,205,0,0,0,0,0,173,0,214,0,0,0,0,0,0,0,215,0,151,0,0,0,243,0,121,0,0,0,190,0,181,0,237,0,34,0,14,0,146,0,78,0,0,0,232,0,152,0,199,0,212,0,238,0,151,0,15,0,198,0,105,0,92,0,229,0,168,0,78,0,139,0,207,0,119,0,122,0,160,0,215,0,177,0,0,0,81,0,71,0,0,0,203,0,109,0,52,0,73,0,44,0,0,0,137,0,199,0,57,0,94,0,123,0,252,0,137,0,73,0,131,0,129,0,207,0,122,0,143,0,65,0,169,0,132,0,67,0,0,0,210,0,240,0,172,0,233,0,192,0,70,0,85,0,251,0,38,0,72,0,0,0,102,0,0,0,0,0,115,0,175,0,135,0,133,0,14,0,62,0,0,0,0,0,50,0,217,0,0,0,0,0,122,0,75,0,224,0,0,0,103,0,24,0,184,0);
signal scenario_full  : scenario_type := (22,31,234,31,234,30,234,29,234,28,44,31,43,31,50,31,7,31,79,31,20,31,108,31,108,30,248,31,161,31,146,31,146,30,146,29,40,31,170,31,16,31,59,31,25,31,82,31,237,31,172,31,6,31,93,31,218,31,218,30,5,31,5,30,18,31,87,31,254,31,4,31,174,31,134,31,164,31,164,30,252,31,70,31,190,31,195,31,18,31,63,31,77,31,170,31,170,30,51,31,140,31,163,31,114,31,114,30,67,31,67,30,78,31,162,31,206,31,46,31,148,31,11,31,174,31,78,31,228,31,150,31,117,31,65,31,151,31,63,31,90,31,119,31,86,31,149,31,40,31,255,31,255,30,201,31,201,30,206,31,105,31,78,31,35,31,83,31,186,31,24,31,5,31,217,31,51,31,52,31,57,31,57,30,208,31,94,31,55,31,55,30,201,31,185,31,185,30,241,31,250,31,182,31,142,31,57,31,57,30,159,31,149,31,232,31,232,30,191,31,144,31,67,31,67,30,67,29,131,31,131,30,79,31,79,30,126,31,160,31,57,31,209,31,169,31,28,31,161,31,38,31,167,31,179,31,163,31,67,31,55,31,149,31,73,31,23,31,143,31,143,30,255,31,235,31,98,31,241,31,26,31,189,31,72,31,72,30,72,29,72,28,72,27,128,31,121,31,108,31,49,31,49,30,191,31,246,31,103,31,103,30,118,31,118,30,151,31,137,31,9,31,9,30,176,31,162,31,210,31,210,30,138,31,138,30,160,31,160,30,245,31,169,31,35,31,23,31,211,31,211,30,118,31,234,31,192,31,192,30,192,29,192,28,169,31,122,31,154,31,154,30,166,31,166,30,33,31,190,31,131,31,164,31,164,30,83,31,137,31,203,31,108,31,209,31,222,31,207,31,106,31,106,30,206,31,41,31,245,31,56,31,56,30,1,31,200,31,227,31,165,31,209,31,209,31,55,31,55,30,4,31,55,31,172,31,35,31,81,31,81,30,81,29,91,31,24,31,208,31,208,30,193,31,85,31,85,30,156,31,41,31,167,31,18,31,18,30,45,31,45,30,41,31,85,31,85,30,190,31,213,31,223,31,152,31,99,31,223,31,3,31,9,31,110,31,238,31,236,31,190,31,26,31,163,31,228,31,32,31,2,31,71,31,48,31,103,31,171,31,171,30,241,31,234,31,48,31,116,31,147,31,147,30,147,29,211,31,156,31,144,31,236,31,56,31,175,31,106,31,106,30,32,31,134,31,147,31,198,31,198,30,108,31,208,31,17,31,17,30,207,31,189,31,99,31,147,31,94,31,68,31,132,31,132,30,238,31,238,30,55,31,198,31,77,31,237,31,237,30,237,29,225,31,181,31,223,31,239,31,214,31,235,31,154,31,39,31,222,31,255,31,255,30,132,31,20,31,92,31,92,30,11,31,11,30,110,31,91,31,189,31,162,31,14,31,14,30,14,29,94,31,159,31,221,31,179,31,113,31,113,30,113,29,113,28,25,31,182,31,104,31,34,31,71,31,209,31,138,31,138,30,14,31,107,31,220,31,165,31,165,30,42,31,158,31,17,31,14,31,123,31,165,31,169,31,78,31,78,30,207,31,188,31,171,31,9,31,3,31,21,31,159,31,159,30,155,31,155,31,221,31,150,31,150,30,44,31,44,30,213,31,181,31,111,31,111,30,111,29,194,31,194,30,24,31,24,30,38,31,194,31,194,30,134,31,202,31,232,31,232,30,234,31,138,31,120,31,16,31,218,31,148,31,106,31,92,31,92,30,163,31,163,30,201,31,47,31,47,30,187,31,79,31,18,31,57,31,57,30,235,31,156,31,27,31,241,31,207,31,105,31,52,31,52,30,174,31,123,31,16,31,23,31,151,31,151,30,151,29,253,31,11,31,11,30,231,31,231,30,231,29,95,31,95,30,108,31,58,31,58,30,166,31,47,31,87,31,41,31,194,31,194,30,194,29,75,31,139,31,242,31,242,30,37,31,167,31,8,31,231,31,79,31,242,31,144,31,144,30,43,31,43,30,44,31,153,31,48,31,127,31,200,31,200,30,94,31,94,30,94,29,113,31,206,31,230,31,172,31,172,30,172,29,172,28,145,31,145,30,219,31,64,31,103,31,103,30,196,31,124,31,55,31,247,31,55,31,142,31,142,30,188,31,188,30,246,31,96,31,10,31,56,31,56,30,125,31,3,31,149,31,209,31,231,31,167,31,226,31,168,31,234,31,92,31,159,31,22,31,38,31,193,31,193,30,220,31,235,31,213,31,68,31,165,31,165,31,242,31,3,31,253,31,137,31,28,31,28,30,28,29,28,28,202,31,171,31,249,31,121,31,214,31,242,31,242,30,242,29,126,31,212,31,135,31,153,31,145,31,45,31,45,30,62,31,8,31,199,31,239,31,239,31,115,31,37,31,226,31,179,31,224,31,171,31,96,31,28,31,28,30,245,31,209,31,245,31,182,31,196,31,111,31,111,30,30,31,30,30,95,31,239,31,239,30,202,31,50,31,151,31,3,31,73,31,155,31,155,30,8,31,12,31,53,31,185,31,56,31,54,31,5,31,171,31,53,31,196,31,121,31,50,31,50,30,83,31,148,31,232,31,199,31,162,31,253,31,32,31,67,31,195,31,104,31,221,31,221,30,219,31,221,31,222,31,186,31,67,31,102,31,204,31,75,31,198,31,230,31,230,30,70,31,135,31,135,30,91,31,230,31,110,31,148,31,148,30,148,29,242,31,242,30,144,31,144,30,144,29,231,31,132,31,214,31,102,31,116,31,205,31,23,31,253,31,169,31,156,31,233,31,233,30,216,31,56,31,213,31,242,31,242,30,209,31,167,31,237,31,151,31,151,30,186,31,119,31,33,31,33,30,99,31,99,30,220,31,121,31,139,31,55,31,81,31,240,31,255,31,64,31,242,31,253,31,211,31,11,31,204,31,231,31,81,31,64,31,52,31,52,30,120,31,199,31,158,31,120,31,120,30,242,31,53,31,123,31,61,31,181,31,55,31,74,31,71,31,79,31,95,31,56,31,4,31,26,31,123,31,100,31,218,31,174,31,178,31,88,31,243,31,243,30,243,29,186,31,184,31,247,31,108,31,11,31,105,31,249,31,249,30,129,31,23,31,155,31,83,31,83,30,83,29,34,31,162,31,248,31,220,31,230,31,244,31,158,31,178,31,74,31,142,31,140,31,93,31,189,31,203,31,146,31,238,31,31,31,187,31,249,31,118,31,76,31,202,31,165,31,165,30,165,29,243,31,255,31,135,31,128,31,128,30,2,31,134,31,195,31,126,31,65,31,62,31,137,31,209,31,39,31,39,30,28,31,28,30,99,31,222,31,254,31,254,30,66,31,69,31,125,31,8,31,154,31,178,31,220,31,253,31,189,31,206,31,253,31,253,30,29,31,194,31,93,31,54,31,54,30,15,31,211,31,243,31,71,31,126,31,126,30,137,31,185,31,241,31,241,30,26,31,155,31,100,31,100,30,118,31,118,30,81,31,154,31,154,30,137,31,207,31,192,31,236,31,218,31,218,30,241,31,103,31,46,31,211,31,211,30,222,31,195,31,33,31,172,31,172,30,182,31,181,31,62,31,139,31,62,31,169,31,169,30,119,31,209,31,209,30,228,31,23,31,23,30,30,31,56,31,251,31,251,30,157,31,48,31,25,31,120,31,51,31,82,31,82,30,161,31,250,31,49,31,180,31,196,31,225,31,225,30,83,31,108,31,160,31,221,31,15,31,165,31,61,31,59,31,61,31,178,31,178,30,178,29,178,28,101,31,81,31,81,30,39,31,247,31,216,31,229,31,133,31,211,31,105,31,105,30,80,31,23,31,23,30,179,31,179,30,26,31,138,31,143,31,81,31,178,31,119,31,182,31,116,31,116,30,116,29,250,31,250,30,250,29,88,31,88,30,187,31,90,31,16,31,81,31,184,31,190,31,171,31,171,30,250,31,253,31,35,31,115,31,108,31,122,31,86,31,170,31,216,31,13,31,150,31,188,31,17,31,49,31,11,31,27,31,139,31,25,31,25,30,153,31,105,31,105,30,105,29,15,31,170,31,205,31,205,30,205,29,173,31,214,31,214,30,214,29,214,28,215,31,151,31,151,30,243,31,121,31,121,30,190,31,181,31,237,31,34,31,14,31,146,31,78,31,78,30,232,31,152,31,199,31,212,31,238,31,151,31,15,31,198,31,105,31,92,31,229,31,168,31,78,31,139,31,207,31,119,31,122,31,160,31,215,31,177,31,177,30,81,31,71,31,71,30,203,31,109,31,52,31,73,31,44,31,44,30,137,31,199,31,57,31,94,31,123,31,252,31,137,31,73,31,131,31,129,31,207,31,122,31,143,31,65,31,169,31,132,31,67,31,67,30,210,31,240,31,172,31,233,31,192,31,70,31,85,31,251,31,38,31,72,31,72,30,102,31,102,30,102,29,115,31,175,31,135,31,133,31,14,31,62,31,62,30,62,29,50,31,217,31,217,30,217,29,122,31,75,31,224,31,224,30,103,31,24,31,184,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
