-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 949;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (172,0,231,0,167,0,238,0,231,0,184,0,228,0,197,0,0,0,165,0,0,0,0,0,91,0,32,0,212,0,108,0,178,0,0,0,75,0,219,0,134,0,164,0,214,0,0,0,227,0,165,0,174,0,99,0,144,0,7,0,100,0,0,0,0,0,160,0,131,0,26,0,81,0,132,0,50,0,190,0,166,0,0,0,119,0,0,0,0,0,0,0,154,0,0,0,0,0,209,0,255,0,241,0,15,0,154,0,99,0,143,0,227,0,80,0,143,0,169,0,0,0,43,0,131,0,166,0,92,0,20,0,113,0,86,0,14,0,188,0,194,0,254,0,0,0,123,0,200,0,119,0,126,0,17,0,109,0,0,0,30,0,229,0,28,0,174,0,29,0,0,0,211,0,0,0,147,0,0,0,0,0,60,0,107,0,130,0,64,0,228,0,22,0,0,0,229,0,0,0,123,0,254,0,208,0,162,0,90,0,65,0,199,0,102,0,216,0,0,0,219,0,0,0,82,0,200,0,0,0,0,0,0,0,11,0,0,0,0,0,0,0,194,0,0,0,62,0,68,0,0,0,111,0,54,0,115,0,0,0,157,0,53,0,176,0,15,0,129,0,76,0,187,0,193,0,194,0,73,0,216,0,59,0,73,0,54,0,146,0,88,0,190,0,5,0,141,0,156,0,201,0,13,0,109,0,121,0,0,0,204,0,0,0,0,0,0,0,0,0,161,0,0,0,149,0,0,0,243,0,177,0,99,0,243,0,80,0,239,0,77,0,34,0,227,0,90,0,9,0,214,0,68,0,151,0,235,0,238,0,247,0,0,0,19,0,210,0,79,0,0,0,0,0,23,0,186,0,20,0,0,0,39,0,0,0,154,0,151,0,229,0,179,0,62,0,59,0,170,0,45,0,101,0,0,0,0,0,0,0,136,0,90,0,100,0,164,0,0,0,226,0,126,0,0,0,197,0,161,0,151,0,82,0,244,0,77,0,0,0,154,0,0,0,158,0,24,0,0,0,20,0,33,0,207,0,246,0,147,0,172,0,138,0,88,0,210,0,135,0,22,0,232,0,123,0,54,0,239,0,0,0,22,0,218,0,0,0,30,0,0,0,129,0,0,0,217,0,167,0,12,0,0,0,148,0,131,0,233,0,84,0,0,0,231,0,36,0,49,0,183,0,232,0,79,0,186,0,158,0,194,0,130,0,0,0,228,0,51,0,227,0,195,0,0,0,211,0,0,0,174,0,0,0,0,0,0,0,7,0,0,0,104,0,235,0,206,0,0,0,0,0,242,0,0,0,62,0,0,0,134,0,0,0,0,0,199,0,0,0,42,0,25,0,0,0,195,0,112,0,137,0,56,0,0,0,4,0,126,0,101,0,40,0,195,0,222,0,243,0,0,0,166,0,161,0,47,0,75,0,217,0,0,0,89,0,163,0,32,0,72,0,190,0,232,0,0,0,107,0,186,0,163,0,199,0,76,0,192,0,195,0,156,0,146,0,104,0,37,0,216,0,138,0,203,0,63,0,210,0,119,0,72,0,159,0,7,0,70,0,240,0,226,0,92,0,246,0,205,0,94,0,91,0,113,0,0,0,3,0,0,0,0,0,0,0,240,0,39,0,94,0,133,0,0,0,56,0,173,0,0,0,0,0,18,0,63,0,246,0,173,0,3,0,148,0,0,0,0,0,242,0,177,0,42,0,158,0,214,0,0,0,235,0,169,0,130,0,167,0,185,0,184,0,0,0,19,0,137,0,180,0,111,0,30,0,167,0,234,0,0,0,10,0,186,0,29,0,53,0,0,0,183,0,64,0,30,0,0,0,130,0,167,0,251,0,53,0,249,0,0,0,202,0,114,0,190,0,130,0,108,0,13,0,113,0,233,0,25,0,0,0,41,0,108,0,160,0,0,0,0,0,12,0,127,0,0,0,46,0,167,0,204,0,114,0,241,0,3,0,0,0,168,0,111,0,0,0,184,0,37,0,202,0,0,0,113,0,0,0,219,0,231,0,237,0,112,0,94,0,199,0,78,0,148,0,122,0,0,0,0,0,22,0,160,0,0,0,58,0,104,0,26,0,0,0,101,0,17,0,77,0,169,0,8,0,92,0,21,0,202,0,85,0,95,0,236,0,6,0,13,0,10,0,129,0,115,0,0,0,26,0,0,0,131,0,97,0,0,0,38,0,232,0,214,0,15,0,191,0,0,0,0,0,238,0,0,0,240,0,0,0,213,0,0,0,0,0,76,0,56,0,160,0,213,0,0,0,164,0,78,0,247,0,228,0,150,0,35,0,115,0,64,0,0,0,97,0,0,0,0,0,110,0,51,0,254,0,174,0,183,0,240,0,122,0,200,0,1,0,0,0,22,0,127,0,182,0,85,0,110,0,86,0,7,0,169,0,143,0,91,0,117,0,0,0,28,0,202,0,127,0,75,0,114,0,209,0,171,0,144,0,58,0,69,0,30,0,91,0,255,0,0,0,0,0,0,0,0,0,211,0,0,0,49,0,154,0,152,0,29,0,195,0,104,0,0,0,162,0,237,0,221,0,0,0,241,0,0,0,123,0,205,0,127,0,39,0,0,0,147,0,13,0,177,0,188,0,90,0,40,0,237,0,0,0,197,0,0,0,0,0,15,0,200,0,61,0,251,0,85,0,218,0,99,0,211,0,0,0,221,0,120,0,159,0,77,0,186,0,18,0,0,0,0,0,0,0,0,0,201,0,176,0,1,0,242,0,153,0,0,0,5,0,0,0,161,0,221,0,80,0,239,0,96,0,122,0,0,0,90,0,122,0,0,0,141,0,243,0,125,0,0,0,194,0,141,0,122,0,0,0,0,0,166,0,88,0,90,0,213,0,0,0,51,0,118,0,16,0,88,0,178,0,231,0,186,0,6,0,127,0,174,0,176,0,99,0,64,0,121,0,92,0,184,0,194,0,93,0,171,0,23,0,0,0,27,0,179,0,159,0,60,0,138,0,62,0,0,0,255,0,254,0,10,0,0,0,209,0,20,0,19,0,0,0,0,0,59,0,47,0,228,0,229,0,31,0,214,0,0,0,182,0,173,0,203,0,169,0,0,0,0,0,201,0,0,0,0,0,0,0,0,0,105,0,152,0,152,0,221,0,42,0,227,0,236,0,78,0,131,0,0,0,198,0,209,0,165,0,98,0,0,0,94,0,110,0,106,0,107,0,16,0,224,0,247,0,185,0,229,0,0,0,242,0,236,0,35,0,14,0,155,0,100,0,0,0,0,0,152,0,67,0,0,0,0,0,113,0,231,0,217,0,0,0,246,0,0,0,181,0,219,0,244,0,56,0,0,0,195,0,0,0,49,0,9,0,0,0,27,0,51,0,200,0,0,0,17,0,225,0,2,0,142,0,0,0,183,0,132,0,161,0,0,0,36,0,222,0,232,0,113,0,62,0,102,0,51,0,205,0,93,0,224,0,168,0,0,0,0,0,172,0,0,0,0,0,22,0,112,0,206,0,170,0,137,0,244,0,153,0,0,0,186,0,74,0,67,0,154,0,135,0,2,0,159,0,211,0,221,0,196,0,0,0,102,0,96,0,8,0,0,0,161,0,15,0,0,0,92,0,180,0,97,0,34,0,0,0,93,0,83,0,203,0,186,0,35,0,200,0,0,0,0,0,136,0,89,0,40,0,167,0,20,0,0,0,79,0,0,0,214,0,0,0,24,0,22,0,193,0,76,0,216,0,18,0,213,0,255,0,34,0,6,0,202,0,0,0,34,0,0,0,236,0,43,0,57,0,155,0,245,0,126,0,0,0,54,0,120,0,0,0,79,0,91,0,0,0,106,0,156,0,0,0,172,0,47,0,235,0,42,0,164,0,0,0,0,0,11,0,0,0,184,0,231,0,29,0,4,0,0,0,0,0,0,0,145,0,0,0,0,0,145,0,105,0,204,0,246,0,0,0,0,0,105,0,10,0,122,0,68,0,87,0,82,0,15,0,98,0,91,0,86,0,233,0,101,0,237,0,174,0,44,0,112,0,119,0,0,0,143,0,166,0,87,0,111,0,61,0,86,0,93,0,207,0,98,0,184,0,173,0,36,0,211,0,0,0,7,0,130,0,78,0,240,0,133,0,60,0,0,0,83,0,132,0,218,0,71,0,0,0,0,0,253,0,241,0,171,0,7,0,65,0,31,0,77,0,148,0,73,0,0,0,107,0,64,0,177,0,0,0,48,0,0,0,149,0,142,0,3,0,85,0,0,0,193,0,67,0,164,0,109,0,0,0);
signal scenario_full  : scenario_type := (172,31,231,31,167,31,238,31,231,31,184,31,228,31,197,31,197,30,165,31,165,30,165,29,91,31,32,31,212,31,108,31,178,31,178,30,75,31,219,31,134,31,164,31,214,31,214,30,227,31,165,31,174,31,99,31,144,31,7,31,100,31,100,30,100,29,160,31,131,31,26,31,81,31,132,31,50,31,190,31,166,31,166,30,119,31,119,30,119,29,119,28,154,31,154,30,154,29,209,31,255,31,241,31,15,31,154,31,99,31,143,31,227,31,80,31,143,31,169,31,169,30,43,31,131,31,166,31,92,31,20,31,113,31,86,31,14,31,188,31,194,31,254,31,254,30,123,31,200,31,119,31,126,31,17,31,109,31,109,30,30,31,229,31,28,31,174,31,29,31,29,30,211,31,211,30,147,31,147,30,147,29,60,31,107,31,130,31,64,31,228,31,22,31,22,30,229,31,229,30,123,31,254,31,208,31,162,31,90,31,65,31,199,31,102,31,216,31,216,30,219,31,219,30,82,31,200,31,200,30,200,29,200,28,11,31,11,30,11,29,11,28,194,31,194,30,62,31,68,31,68,30,111,31,54,31,115,31,115,30,157,31,53,31,176,31,15,31,129,31,76,31,187,31,193,31,194,31,73,31,216,31,59,31,73,31,54,31,146,31,88,31,190,31,5,31,141,31,156,31,201,31,13,31,109,31,121,31,121,30,204,31,204,30,204,29,204,28,204,27,161,31,161,30,149,31,149,30,243,31,177,31,99,31,243,31,80,31,239,31,77,31,34,31,227,31,90,31,9,31,214,31,68,31,151,31,235,31,238,31,247,31,247,30,19,31,210,31,79,31,79,30,79,29,23,31,186,31,20,31,20,30,39,31,39,30,154,31,151,31,229,31,179,31,62,31,59,31,170,31,45,31,101,31,101,30,101,29,101,28,136,31,90,31,100,31,164,31,164,30,226,31,126,31,126,30,197,31,161,31,151,31,82,31,244,31,77,31,77,30,154,31,154,30,158,31,24,31,24,30,20,31,33,31,207,31,246,31,147,31,172,31,138,31,88,31,210,31,135,31,22,31,232,31,123,31,54,31,239,31,239,30,22,31,218,31,218,30,30,31,30,30,129,31,129,30,217,31,167,31,12,31,12,30,148,31,131,31,233,31,84,31,84,30,231,31,36,31,49,31,183,31,232,31,79,31,186,31,158,31,194,31,130,31,130,30,228,31,51,31,227,31,195,31,195,30,211,31,211,30,174,31,174,30,174,29,174,28,7,31,7,30,104,31,235,31,206,31,206,30,206,29,242,31,242,30,62,31,62,30,134,31,134,30,134,29,199,31,199,30,42,31,25,31,25,30,195,31,112,31,137,31,56,31,56,30,4,31,126,31,101,31,40,31,195,31,222,31,243,31,243,30,166,31,161,31,47,31,75,31,217,31,217,30,89,31,163,31,32,31,72,31,190,31,232,31,232,30,107,31,186,31,163,31,199,31,76,31,192,31,195,31,156,31,146,31,104,31,37,31,216,31,138,31,203,31,63,31,210,31,119,31,72,31,159,31,7,31,70,31,240,31,226,31,92,31,246,31,205,31,94,31,91,31,113,31,113,30,3,31,3,30,3,29,3,28,240,31,39,31,94,31,133,31,133,30,56,31,173,31,173,30,173,29,18,31,63,31,246,31,173,31,3,31,148,31,148,30,148,29,242,31,177,31,42,31,158,31,214,31,214,30,235,31,169,31,130,31,167,31,185,31,184,31,184,30,19,31,137,31,180,31,111,31,30,31,167,31,234,31,234,30,10,31,186,31,29,31,53,31,53,30,183,31,64,31,30,31,30,30,130,31,167,31,251,31,53,31,249,31,249,30,202,31,114,31,190,31,130,31,108,31,13,31,113,31,233,31,25,31,25,30,41,31,108,31,160,31,160,30,160,29,12,31,127,31,127,30,46,31,167,31,204,31,114,31,241,31,3,31,3,30,168,31,111,31,111,30,184,31,37,31,202,31,202,30,113,31,113,30,219,31,231,31,237,31,112,31,94,31,199,31,78,31,148,31,122,31,122,30,122,29,22,31,160,31,160,30,58,31,104,31,26,31,26,30,101,31,17,31,77,31,169,31,8,31,92,31,21,31,202,31,85,31,95,31,236,31,6,31,13,31,10,31,129,31,115,31,115,30,26,31,26,30,131,31,97,31,97,30,38,31,232,31,214,31,15,31,191,31,191,30,191,29,238,31,238,30,240,31,240,30,213,31,213,30,213,29,76,31,56,31,160,31,213,31,213,30,164,31,78,31,247,31,228,31,150,31,35,31,115,31,64,31,64,30,97,31,97,30,97,29,110,31,51,31,254,31,174,31,183,31,240,31,122,31,200,31,1,31,1,30,22,31,127,31,182,31,85,31,110,31,86,31,7,31,169,31,143,31,91,31,117,31,117,30,28,31,202,31,127,31,75,31,114,31,209,31,171,31,144,31,58,31,69,31,30,31,91,31,255,31,255,30,255,29,255,28,255,27,211,31,211,30,49,31,154,31,152,31,29,31,195,31,104,31,104,30,162,31,237,31,221,31,221,30,241,31,241,30,123,31,205,31,127,31,39,31,39,30,147,31,13,31,177,31,188,31,90,31,40,31,237,31,237,30,197,31,197,30,197,29,15,31,200,31,61,31,251,31,85,31,218,31,99,31,211,31,211,30,221,31,120,31,159,31,77,31,186,31,18,31,18,30,18,29,18,28,18,27,201,31,176,31,1,31,242,31,153,31,153,30,5,31,5,30,161,31,221,31,80,31,239,31,96,31,122,31,122,30,90,31,122,31,122,30,141,31,243,31,125,31,125,30,194,31,141,31,122,31,122,30,122,29,166,31,88,31,90,31,213,31,213,30,51,31,118,31,16,31,88,31,178,31,231,31,186,31,6,31,127,31,174,31,176,31,99,31,64,31,121,31,92,31,184,31,194,31,93,31,171,31,23,31,23,30,27,31,179,31,159,31,60,31,138,31,62,31,62,30,255,31,254,31,10,31,10,30,209,31,20,31,19,31,19,30,19,29,59,31,47,31,228,31,229,31,31,31,214,31,214,30,182,31,173,31,203,31,169,31,169,30,169,29,201,31,201,30,201,29,201,28,201,27,105,31,152,31,152,31,221,31,42,31,227,31,236,31,78,31,131,31,131,30,198,31,209,31,165,31,98,31,98,30,94,31,110,31,106,31,107,31,16,31,224,31,247,31,185,31,229,31,229,30,242,31,236,31,35,31,14,31,155,31,100,31,100,30,100,29,152,31,67,31,67,30,67,29,113,31,231,31,217,31,217,30,246,31,246,30,181,31,219,31,244,31,56,31,56,30,195,31,195,30,49,31,9,31,9,30,27,31,51,31,200,31,200,30,17,31,225,31,2,31,142,31,142,30,183,31,132,31,161,31,161,30,36,31,222,31,232,31,113,31,62,31,102,31,51,31,205,31,93,31,224,31,168,31,168,30,168,29,172,31,172,30,172,29,22,31,112,31,206,31,170,31,137,31,244,31,153,31,153,30,186,31,74,31,67,31,154,31,135,31,2,31,159,31,211,31,221,31,196,31,196,30,102,31,96,31,8,31,8,30,161,31,15,31,15,30,92,31,180,31,97,31,34,31,34,30,93,31,83,31,203,31,186,31,35,31,200,31,200,30,200,29,136,31,89,31,40,31,167,31,20,31,20,30,79,31,79,30,214,31,214,30,24,31,22,31,193,31,76,31,216,31,18,31,213,31,255,31,34,31,6,31,202,31,202,30,34,31,34,30,236,31,43,31,57,31,155,31,245,31,126,31,126,30,54,31,120,31,120,30,79,31,91,31,91,30,106,31,156,31,156,30,172,31,47,31,235,31,42,31,164,31,164,30,164,29,11,31,11,30,184,31,231,31,29,31,4,31,4,30,4,29,4,28,145,31,145,30,145,29,145,31,105,31,204,31,246,31,246,30,246,29,105,31,10,31,122,31,68,31,87,31,82,31,15,31,98,31,91,31,86,31,233,31,101,31,237,31,174,31,44,31,112,31,119,31,119,30,143,31,166,31,87,31,111,31,61,31,86,31,93,31,207,31,98,31,184,31,173,31,36,31,211,31,211,30,7,31,130,31,78,31,240,31,133,31,60,31,60,30,83,31,132,31,218,31,71,31,71,30,71,29,253,31,241,31,171,31,7,31,65,31,31,31,77,31,148,31,73,31,73,30,107,31,64,31,177,31,177,30,48,31,48,30,149,31,142,31,3,31,85,31,85,30,193,31,67,31,164,31,109,31,109,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
