-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_760 is
end project_tb_760;

architecture project_tb_arch_760 of project_tb_760 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 980;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (197,0,91,0,29,0,0,0,0,0,81,0,195,0,156,0,176,0,0,0,188,0,186,0,248,0,177,0,37,0,193,0,19,0,0,0,109,0,224,0,10,0,0,0,165,0,0,0,171,0,201,0,33,0,238,0,91,0,0,0,124,0,71,0,150,0,0,0,138,0,2,0,65,0,226,0,22,0,221,0,158,0,0,0,0,0,114,0,135,0,0,0,120,0,179,0,0,0,0,0,0,0,0,0,131,0,57,0,165,0,42,0,0,0,5,0,142,0,31,0,18,0,130,0,135,0,134,0,188,0,41,0,70,0,0,0,39,0,0,0,0,0,66,0,71,0,110,0,0,0,0,0,47,0,36,0,12,0,247,0,0,0,178,0,143,0,254,0,94,0,0,0,0,0,0,0,240,0,114,0,0,0,134,0,160,0,0,0,136,0,7,0,123,0,200,0,18,0,0,0,50,0,24,0,0,0,126,0,55,0,190,0,228,0,24,0,0,0,92,0,0,0,55,0,70,0,151,0,16,0,1,0,245,0,0,0,0,0,43,0,11,0,87,0,210,0,54,0,85,0,9,0,141,0,102,0,105,0,42,0,24,0,246,0,250,0,45,0,0,0,0,0,66,0,203,0,147,0,156,0,0,0,94,0,0,0,222,0,160,0,192,0,223,0,220,0,31,0,123,0,36,0,240,0,20,0,24,0,254,0,0,0,0,0,251,0,77,0,161,0,182,0,54,0,0,0,129,0,242,0,215,0,192,0,17,0,105,0,24,0,22,0,0,0,44,0,124,0,0,0,113,0,222,0,81,0,39,0,59,0,79,0,8,0,0,0,22,0,0,0,254,0,45,0,95,0,112,0,19,0,116,0,113,0,184,0,34,0,151,0,134,0,0,0,223,0,114,0,211,0,166,0,0,0,42,0,90,0,178,0,223,0,133,0,0,0,108,0,162,0,228,0,236,0,204,0,73,0,223,0,0,0,196,0,195,0,91,0,0,0,188,0,79,0,30,0,0,0,222,0,0,0,188,0,92,0,126,0,61,0,164,0,57,0,0,0,157,0,50,0,209,0,188,0,175,0,246,0,0,0,59,0,159,0,248,0,107,0,237,0,216,0,217,0,151,0,82,0,218,0,21,0,92,0,0,0,207,0,180,0,71,0,0,0,253,0,255,0,57,0,120,0,0,0,49,0,245,0,221,0,204,0,39,0,154,0,122,0,0,0,27,0,21,0,206,0,0,0,207,0,202,0,0,0,121,0,169,0,0,0,27,0,154,0,253,0,57,0,209,0,179,0,229,0,0,0,0,0,83,0,112,0,69,0,0,0,52,0,106,0,17,0,0,0,200,0,20,0,159,0,0,0,71,0,31,0,0,0,0,0,0,0,24,0,99,0,0,0,157,0,0,0,64,0,124,0,8,0,211,0,220,0,182,0,90,0,6,0,58,0,22,0,215,0,141,0,213,0,249,0,140,0,0,0,57,0,67,0,113,0,37,0,35,0,234,0,21,0,227,0,119,0,0,0,61,0,227,0,0,0,49,0,224,0,217,0,0,0,76,0,51,0,159,0,0,0,237,0,178,0,177,0,30,0,78,0,0,0,116,0,240,0,78,0,0,0,164,0,147,0,119,0,107,0,169,0,60,0,105,0,3,0,170,0,76,0,156,0,185,0,18,0,123,0,149,0,70,0,2,0,73,0,168,0,0,0,0,0,47,0,86,0,189,0,206,0,34,0,129,0,53,0,27,0,44,0,230,0,0,0,49,0,57,0,104,0,0,0,57,0,35,0,133,0,252,0,183,0,209,0,206,0,135,0,96,0,97,0,50,0,245,0,76,0,34,0,0,0,209,0,245,0,4,0,1,0,232,0,175,0,175,0,0,0,24,0,0,0,176,0,236,0,47,0,61,0,213,0,18,0,166,0,0,0,230,0,0,0,13,0,44,0,183,0,110,0,204,0,0,0,0,0,174,0,0,0,156,0,0,0,211,0,141,0,0,0,0,0,22,0,39,0,0,0,137,0,92,0,0,0,177,0,131,0,214,0,230,0,0,0,241,0,116,0,78,0,33,0,230,0,0,0,188,0,0,0,120,0,84,0,154,0,0,0,238,0,81,0,82,0,106,0,173,0,216,0,186,0,83,0,183,0,96,0,26,0,146,0,227,0,97,0,45,0,90,0,0,0,106,0,194,0,74,0,151,0,144,0,0,0,92,0,80,0,0,0,112,0,198,0,182,0,253,0,245,0,0,0,253,0,0,0,0,0,187,0,28,0,141,0,185,0,148,0,141,0,78,0,52,0,236,0,130,0,129,0,242,0,187,0,0,0,255,0,77,0,167,0,0,0,170,0,84,0,74,0,138,0,0,0,118,0,150,0,162,0,120,0,0,0,250,0,139,0,59,0,0,0,0,0,141,0,0,0,174,0,66,0,0,0,163,0,129,0,148,0,253,0,20,0,0,0,0,0,94,0,9,0,123,0,0,0,173,0,25,0,133,0,0,0,204,0,27,0,0,0,0,0,247,0,129,0,54,0,166,0,48,0,10,0,202,0,0,0,0,0,153,0,0,0,80,0,0,0,18,0,60,0,208,0,0,0,120,0,0,0,159,0,111,0,84,0,44,0,49,0,234,0,0,0,93,0,0,0,245,0,95,0,44,0,11,0,241,0,65,0,248,0,129,0,196,0,71,0,15,0,168,0,108,0,136,0,47,0,0,0,72,0,229,0,243,0,0,0,127,0,20,0,124,0,179,0,216,0,85,0,0,0,31,0,71,0,219,0,0,0,83,0,103,0,139,0,0,0,0,0,217,0,226,0,46,0,63,0,79,0,227,0,217,0,192,0,0,0,225,0,0,0,174,0,9,0,210,0,63,0,0,0,129,0,0,0,236,0,124,0,0,0,0,0,106,0,0,0,67,0,177,0,139,0,102,0,0,0,227,0,0,0,19,0,0,0,109,0,18,0,0,0,0,0,26,0,50,0,24,0,0,0,160,0,57,0,51,0,101,0,18,0,47,0,150,0,104,0,173,0,193,0,77,0,0,0,151,0,237,0,252,0,113,0,52,0,178,0,127,0,42,0,0,0,162,0,43,0,65,0,148,0,0,0,68,0,20,0,0,0,132,0,0,0,47,0,0,0,18,0,203,0,0,0,0,0,189,0,140,0,213,0,48,0,176,0,244,0,0,0,148,0,229,0,251,0,201,0,75,0,109,0,242,0,205,0,11,0,178,0,205,0,41,0,39,0,161,0,252,0,27,0,54,0,225,0,144,0,36,0,0,0,0,0,46,0,203,0,60,0,122,0,202,0,63,0,125,0,228,0,0,0,81,0,119,0,106,0,116,0,38,0,8,0,0,0,179,0,211,0,0,0,77,0,152,0,117,0,219,0,81,0,0,0,20,0,0,0,245,0,142,0,227,0,117,0,71,0,108,0,233,0,120,0,0,0,117,0,184,0,166,0,97,0,106,0,174,0,241,0,47,0,142,0,105,0,20,0,0,0,137,0,0,0,0,0,41,0,144,0,87,0,240,0,0,0,5,0,174,0,26,0,146,0,58,0,214,0,49,0,223,0,0,0,136,0,112,0,74,0,149,0,57,0,243,0,0,0,66,0,176,0,180,0,0,0,66,0,63,0,207,0,254,0,97,0,174,0,219,0,203,0,222,0,230,0,0,0,110,0,189,0,49,0,212,0,131,0,120,0,249,0,226,0,0,0,0,0,191,0,73,0,143,0,101,0,206,0,161,0,221,0,0,0,242,0,125,0,110,0,177,0,149,0,143,0,79,0,43,0,215,0,13,0,248,0,243,0,0,0,0,0,0,0,200,0,185,0,212,0,192,0,122,0,0,0,89,0,136,0,85,0,210,0,0,0,248,0,0,0,97,0,227,0,53,0,164,0,254,0,0,0,69,0,191,0,0,0,193,0,24,0,0,0,19,0,196,0,0,0,109,0,59,0,0,0,66,0,151,0,21,0,154,0,0,0,249,0,247,0,114,0,59,0,0,0,43,0,73,0,175,0,0,0,0,0,175,0,12,0,117,0,135,0,154,0,0,0,10,0,29,0,0,0,0,0,219,0,75,0,12,0,66,0,170,0,0,0,91,0,158,0,183,0,227,0,202,0,239,0,239,0,47,0,170,0,25,0,55,0,0,0,250,0,0,0,0,0,195,0,17,0,0,0,228,0,9,0,81,0,0,0,3,0,206,0,131,0,105,0,216,0,216,0,228,0,196,0,165,0,5,0,69,0,172,0,81,0,169,0,124,0,21,0,181,0,92,0,36,0,249,0,191,0,201,0,7,0,28,0,242,0,65,0,61,0,247,0,220,0,193,0,252,0,194,0,180,0,0,0,0,0,128,0,203,0,108,0,169,0,183,0,0,0,0,0,0,0,102,0,40,0,112,0);
signal scenario_full  : scenario_type := (197,31,91,31,29,31,29,30,29,29,81,31,195,31,156,31,176,31,176,30,188,31,186,31,248,31,177,31,37,31,193,31,19,31,19,30,109,31,224,31,10,31,10,30,165,31,165,30,171,31,201,31,33,31,238,31,91,31,91,30,124,31,71,31,150,31,150,30,138,31,2,31,65,31,226,31,22,31,221,31,158,31,158,30,158,29,114,31,135,31,135,30,120,31,179,31,179,30,179,29,179,28,179,27,131,31,57,31,165,31,42,31,42,30,5,31,142,31,31,31,18,31,130,31,135,31,134,31,188,31,41,31,70,31,70,30,39,31,39,30,39,29,66,31,71,31,110,31,110,30,110,29,47,31,36,31,12,31,247,31,247,30,178,31,143,31,254,31,94,31,94,30,94,29,94,28,240,31,114,31,114,30,134,31,160,31,160,30,136,31,7,31,123,31,200,31,18,31,18,30,50,31,24,31,24,30,126,31,55,31,190,31,228,31,24,31,24,30,92,31,92,30,55,31,70,31,151,31,16,31,1,31,245,31,245,30,245,29,43,31,11,31,87,31,210,31,54,31,85,31,9,31,141,31,102,31,105,31,42,31,24,31,246,31,250,31,45,31,45,30,45,29,66,31,203,31,147,31,156,31,156,30,94,31,94,30,222,31,160,31,192,31,223,31,220,31,31,31,123,31,36,31,240,31,20,31,24,31,254,31,254,30,254,29,251,31,77,31,161,31,182,31,54,31,54,30,129,31,242,31,215,31,192,31,17,31,105,31,24,31,22,31,22,30,44,31,124,31,124,30,113,31,222,31,81,31,39,31,59,31,79,31,8,31,8,30,22,31,22,30,254,31,45,31,95,31,112,31,19,31,116,31,113,31,184,31,34,31,151,31,134,31,134,30,223,31,114,31,211,31,166,31,166,30,42,31,90,31,178,31,223,31,133,31,133,30,108,31,162,31,228,31,236,31,204,31,73,31,223,31,223,30,196,31,195,31,91,31,91,30,188,31,79,31,30,31,30,30,222,31,222,30,188,31,92,31,126,31,61,31,164,31,57,31,57,30,157,31,50,31,209,31,188,31,175,31,246,31,246,30,59,31,159,31,248,31,107,31,237,31,216,31,217,31,151,31,82,31,218,31,21,31,92,31,92,30,207,31,180,31,71,31,71,30,253,31,255,31,57,31,120,31,120,30,49,31,245,31,221,31,204,31,39,31,154,31,122,31,122,30,27,31,21,31,206,31,206,30,207,31,202,31,202,30,121,31,169,31,169,30,27,31,154,31,253,31,57,31,209,31,179,31,229,31,229,30,229,29,83,31,112,31,69,31,69,30,52,31,106,31,17,31,17,30,200,31,20,31,159,31,159,30,71,31,31,31,31,30,31,29,31,28,24,31,99,31,99,30,157,31,157,30,64,31,124,31,8,31,211,31,220,31,182,31,90,31,6,31,58,31,22,31,215,31,141,31,213,31,249,31,140,31,140,30,57,31,67,31,113,31,37,31,35,31,234,31,21,31,227,31,119,31,119,30,61,31,227,31,227,30,49,31,224,31,217,31,217,30,76,31,51,31,159,31,159,30,237,31,178,31,177,31,30,31,78,31,78,30,116,31,240,31,78,31,78,30,164,31,147,31,119,31,107,31,169,31,60,31,105,31,3,31,170,31,76,31,156,31,185,31,18,31,123,31,149,31,70,31,2,31,73,31,168,31,168,30,168,29,47,31,86,31,189,31,206,31,34,31,129,31,53,31,27,31,44,31,230,31,230,30,49,31,57,31,104,31,104,30,57,31,35,31,133,31,252,31,183,31,209,31,206,31,135,31,96,31,97,31,50,31,245,31,76,31,34,31,34,30,209,31,245,31,4,31,1,31,232,31,175,31,175,31,175,30,24,31,24,30,176,31,236,31,47,31,61,31,213,31,18,31,166,31,166,30,230,31,230,30,13,31,44,31,183,31,110,31,204,31,204,30,204,29,174,31,174,30,156,31,156,30,211,31,141,31,141,30,141,29,22,31,39,31,39,30,137,31,92,31,92,30,177,31,131,31,214,31,230,31,230,30,241,31,116,31,78,31,33,31,230,31,230,30,188,31,188,30,120,31,84,31,154,31,154,30,238,31,81,31,82,31,106,31,173,31,216,31,186,31,83,31,183,31,96,31,26,31,146,31,227,31,97,31,45,31,90,31,90,30,106,31,194,31,74,31,151,31,144,31,144,30,92,31,80,31,80,30,112,31,198,31,182,31,253,31,245,31,245,30,253,31,253,30,253,29,187,31,28,31,141,31,185,31,148,31,141,31,78,31,52,31,236,31,130,31,129,31,242,31,187,31,187,30,255,31,77,31,167,31,167,30,170,31,84,31,74,31,138,31,138,30,118,31,150,31,162,31,120,31,120,30,250,31,139,31,59,31,59,30,59,29,141,31,141,30,174,31,66,31,66,30,163,31,129,31,148,31,253,31,20,31,20,30,20,29,94,31,9,31,123,31,123,30,173,31,25,31,133,31,133,30,204,31,27,31,27,30,27,29,247,31,129,31,54,31,166,31,48,31,10,31,202,31,202,30,202,29,153,31,153,30,80,31,80,30,18,31,60,31,208,31,208,30,120,31,120,30,159,31,111,31,84,31,44,31,49,31,234,31,234,30,93,31,93,30,245,31,95,31,44,31,11,31,241,31,65,31,248,31,129,31,196,31,71,31,15,31,168,31,108,31,136,31,47,31,47,30,72,31,229,31,243,31,243,30,127,31,20,31,124,31,179,31,216,31,85,31,85,30,31,31,71,31,219,31,219,30,83,31,103,31,139,31,139,30,139,29,217,31,226,31,46,31,63,31,79,31,227,31,217,31,192,31,192,30,225,31,225,30,174,31,9,31,210,31,63,31,63,30,129,31,129,30,236,31,124,31,124,30,124,29,106,31,106,30,67,31,177,31,139,31,102,31,102,30,227,31,227,30,19,31,19,30,109,31,18,31,18,30,18,29,26,31,50,31,24,31,24,30,160,31,57,31,51,31,101,31,18,31,47,31,150,31,104,31,173,31,193,31,77,31,77,30,151,31,237,31,252,31,113,31,52,31,178,31,127,31,42,31,42,30,162,31,43,31,65,31,148,31,148,30,68,31,20,31,20,30,132,31,132,30,47,31,47,30,18,31,203,31,203,30,203,29,189,31,140,31,213,31,48,31,176,31,244,31,244,30,148,31,229,31,251,31,201,31,75,31,109,31,242,31,205,31,11,31,178,31,205,31,41,31,39,31,161,31,252,31,27,31,54,31,225,31,144,31,36,31,36,30,36,29,46,31,203,31,60,31,122,31,202,31,63,31,125,31,228,31,228,30,81,31,119,31,106,31,116,31,38,31,8,31,8,30,179,31,211,31,211,30,77,31,152,31,117,31,219,31,81,31,81,30,20,31,20,30,245,31,142,31,227,31,117,31,71,31,108,31,233,31,120,31,120,30,117,31,184,31,166,31,97,31,106,31,174,31,241,31,47,31,142,31,105,31,20,31,20,30,137,31,137,30,137,29,41,31,144,31,87,31,240,31,240,30,5,31,174,31,26,31,146,31,58,31,214,31,49,31,223,31,223,30,136,31,112,31,74,31,149,31,57,31,243,31,243,30,66,31,176,31,180,31,180,30,66,31,63,31,207,31,254,31,97,31,174,31,219,31,203,31,222,31,230,31,230,30,110,31,189,31,49,31,212,31,131,31,120,31,249,31,226,31,226,30,226,29,191,31,73,31,143,31,101,31,206,31,161,31,221,31,221,30,242,31,125,31,110,31,177,31,149,31,143,31,79,31,43,31,215,31,13,31,248,31,243,31,243,30,243,29,243,28,200,31,185,31,212,31,192,31,122,31,122,30,89,31,136,31,85,31,210,31,210,30,248,31,248,30,97,31,227,31,53,31,164,31,254,31,254,30,69,31,191,31,191,30,193,31,24,31,24,30,19,31,196,31,196,30,109,31,59,31,59,30,66,31,151,31,21,31,154,31,154,30,249,31,247,31,114,31,59,31,59,30,43,31,73,31,175,31,175,30,175,29,175,31,12,31,117,31,135,31,154,31,154,30,10,31,29,31,29,30,29,29,219,31,75,31,12,31,66,31,170,31,170,30,91,31,158,31,183,31,227,31,202,31,239,31,239,31,47,31,170,31,25,31,55,31,55,30,250,31,250,30,250,29,195,31,17,31,17,30,228,31,9,31,81,31,81,30,3,31,206,31,131,31,105,31,216,31,216,31,228,31,196,31,165,31,5,31,69,31,172,31,81,31,169,31,124,31,21,31,181,31,92,31,36,31,249,31,191,31,201,31,7,31,28,31,242,31,65,31,61,31,247,31,220,31,193,31,252,31,194,31,180,31,180,30,180,29,128,31,203,31,108,31,169,31,183,31,183,30,183,29,183,28,102,31,40,31,112,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
