-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 919;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (70,0,164,0,157,0,244,0,116,0,30,0,33,0,0,0,212,0,172,0,46,0,35,0,177,0,0,0,166,0,166,0,0,0,29,0,168,0,227,0,8,0,17,0,233,0,106,0,0,0,0,0,141,0,55,0,111,0,76,0,0,0,248,0,98,0,0,0,140,0,11,0,248,0,69,0,179,0,31,0,232,0,0,0,0,0,176,0,4,0,231,0,38,0,107,0,212,0,9,0,176,0,228,0,122,0,197,0,0,0,38,0,37,0,228,0,14,0,0,0,208,0,100,0,215,0,158,0,39,0,39,0,201,0,125,0,57,0,244,0,219,0,21,0,144,0,228,0,157,0,10,0,115,0,0,0,201,0,0,0,0,0,0,0,199,0,188,0,134,0,23,0,214,0,214,0,155,0,126,0,227,0,0,0,128,0,189,0,0,0,70,0,25,0,0,0,232,0,0,0,169,0,194,0,137,0,60,0,0,0,89,0,113,0,159,0,203,0,78,0,0,0,0,0,37,0,53,0,167,0,148,0,0,0,150,0,214,0,7,0,212,0,0,0,0,0,104,0,0,0,197,0,175,0,111,0,218,0,83,0,247,0,0,0,217,0,57,0,191,0,138,0,0,0,158,0,46,0,108,0,170,0,57,0,202,0,188,0,111,0,0,0,105,0,168,0,40,0,241,0,110,0,40,0,249,0,162,0,0,0,150,0,136,0,38,0,157,0,182,0,126,0,0,0,92,0,49,0,192,0,254,0,254,0,33,0,70,0,32,0,0,0,49,0,149,0,0,0,254,0,20,0,244,0,234,0,0,0,123,0,0,0,90,0,122,0,122,0,79,0,41,0,98,0,219,0,176,0,151,0,0,0,188,0,111,0,0,0,126,0,227,0,100,0,95,0,46,0,0,0,104,0,187,0,22,0,49,0,100,0,52,0,0,0,15,0,129,0,0,0,60,0,157,0,92,0,48,0,4,0,223,0,189,0,152,0,224,0,0,0,0,0,137,0,0,0,103,0,50,0,169,0,154,0,24,0,27,0,0,0,81,0,120,0,127,0,14,0,89,0,128,0,38,0,0,0,124,0,254,0,39,0,146,0,236,0,80,0,0,0,251,0,0,0,183,0,189,0,0,0,126,0,41,0,212,0,0,0,0,0,0,0,0,0,0,0,50,0,239,0,152,0,0,0,251,0,174,0,19,0,51,0,186,0,153,0,85,0,230,0,80,0,0,0,0,0,106,0,134,0,200,0,214,0,91,0,124,0,204,0,32,0,0,0,203,0,217,0,242,0,170,0,138,0,41,0,94,0,151,0,198,0,104,0,109,0,188,0,109,0,7,0,223,0,138,0,234,0,211,0,129,0,124,0,0,0,0,0,0,0,21,0,164,0,0,0,25,0,0,0,0,0,184,0,0,0,12,0,96,0,199,0,0,0,154,0,157,0,0,0,227,0,207,0,150,0,0,0,40,0,146,0,21,0,71,0,0,0,6,0,17,0,129,0,22,0,0,0,223,0,91,0,3,0,114,0,230,0,141,0,0,0,166,0,49,0,0,0,73,0,70,0,11,0,228,0,146,0,0,0,0,0,103,0,75,0,0,0,101,0,37,0,0,0,230,0,166,0,249,0,92,0,0,0,165,0,20,0,19,0,27,0,0,0,128,0,111,0,0,0,24,0,68,0,0,0,163,0,176,0,55,0,56,0,0,0,92,0,57,0,16,0,39,0,0,0,228,0,0,0,127,0,219,0,47,0,86,0,205,0,115,0,38,0,0,0,220,0,226,0,180,0,75,0,172,0,89,0,40,0,232,0,47,0,39,0,69,0,224,0,4,0,198,0,0,0,239,0,254,0,34,0,218,0,221,0,250,0,100,0,49,0,133,0,3,0,11,0,0,0,248,0,211,0,7,0,76,0,205,0,180,0,0,0,0,0,47,0,181,0,61,0,158,0,0,0,37,0,75,0,238,0,97,0,46,0,68,0,132,0,49,0,61,0,0,0,167,0,28,0,152,0,0,0,128,0,114,0,211,0,120,0,217,0,114,0,0,0,208,0,0,0,26,0,121,0,0,0,181,0,246,0,8,0,0,0,209,0,247,0,166,0,0,0,37,0,123,0,163,0,150,0,33,0,0,0,32,0,138,0,110,0,204,0,79,0,0,0,167,0,183,0,16,0,19,0,69,0,131,0,190,0,0,0,5,0,0,0,163,0,151,0,116,0,44,0,34,0,115,0,0,0,0,0,0,0,0,0,47,0,96,0,199,0,216,0,169,0,185,0,151,0,230,0,100,0,0,0,197,0,0,0,0,0,101,0,99,0,13,0,174,0,95,0,74,0,0,0,243,0,194,0,201,0,222,0,3,0,235,0,119,0,203,0,98,0,233,0,136,0,208,0,34,0,85,0,30,0,179,0,155,0,244,0,200,0,121,0,0,0,146,0,170,0,206,0,78,0,97,0,34,0,20,0,63,0,25,0,182,0,134,0,145,0,163,0,178,0,245,0,29,0,45,0,0,0,229,0,220,0,140,0,118,0,49,0,199,0,247,0,34,0,171,0,114,0,169,0,209,0,105,0,236,0,184,0,180,0,0,0,71,0,41,0,229,0,98,0,197,0,0,0,216,0,219,0,41,0,197,0,49,0,205,0,254,0,27,0,0,0,212,0,105,0,36,0,195,0,232,0,253,0,31,0,189,0,194,0,48,0,234,0,0,0,226,0,238,0,151,0,114,0,0,0,122,0,140,0,55,0,222,0,118,0,255,0,213,0,60,0,13,0,162,0,168,0,20,0,123,0,0,0,83,0,199,0,233,0,193,0,232,0,255,0,224,0,0,0,120,0,223,0,143,0,221,0,0,0,231,0,0,0,187,0,251,0,243,0,27,0,91,0,37,0,24,0,134,0,0,0,115,0,148,0,254,0,144,0,0,0,0,0,155,0,46,0,162,0,129,0,84,0,4,0,247,0,215,0,158,0,185,0,60,0,0,0,75,0,143,0,38,0,0,0,78,0,249,0,0,0,154,0,87,0,254,0,211,0,143,0,181,0,3,0,22,0,108,0,204,0,139,0,74,0,201,0,157,0,23,0,100,0,0,0,203,0,251,0,44,0,52,0,21,0,53,0,0,0,0,0,0,0,85,0,19,0,0,0,254,0,210,0,21,0,62,0,0,0,11,0,227,0,22,0,23,0,0,0,0,0,136,0,108,0,25,0,189,0,0,0,179,0,48,0,0,0,244,0,217,0,9,0,0,0,107,0,153,0,0,0,127,0,207,0,23,0,210,0,202,0,27,0,183,0,198,0,231,0,101,0,146,0,60,0,127,0,9,0,220,0,48,0,134,0,0,0,29,0,28,0,67,0,0,0,183,0,0,0,147,0,124,0,224,0,123,0,221,0,0,0,0,0,185,0,241,0,212,0,40,0,152,0,46,0,77,0,0,0,244,0,0,0,129,0,49,0,0,0,47,0,240,0,51,0,244,0,50,0,5,0,18,0,40,0,0,0,148,0,0,0,235,0,254,0,0,0,152,0,0,0,13,0,110,0,149,0,30,0,249,0,20,0,40,0,140,0,24,0,149,0,196,0,88,0,145,0,0,0,154,0,80,0,88,0,216,0,198,0,211,0,60,0,0,0,175,0,57,0,148,0,0,0,193,0,0,0,0,0,193,0,0,0,0,0,185,0,101,0,114,0,0,0,51,0,123,0,232,0,70,0,179,0,57,0,171,0,0,0,0,0,100,0,246,0,103,0,19,0,0,0,102,0,0,0,0,0,68,0,25,0,48,0,0,0,15,0,76,0,153,0,238,0,0,0,0,0,107,0,22,0,114,0,116,0,170,0,0,0,0,0,0,0,200,0,207,0,181,0,166,0,130,0,16,0,109,0,231,0,198,0,189,0,1,0,217,0,0,0,34,0,91,0,67,0,18,0,162,0,0,0,19,0,152,0,83,0,247,0,173,0,0,0,0,0,220,0,147,0,139,0,0,0,169,0,62,0,227,0,151,0,152,0,88,0,97,0,206,0,123,0,81,0,152,0,0,0,135,0,159,0,0,0,0,0,172,0,193,0,202,0,39,0,0,0,127,0,0,0,116,0,69,0,0,0,102,0,100,0,6,0,159,0,0,0,132,0,153,0);
signal scenario_full  : scenario_type := (70,31,164,31,157,31,244,31,116,31,30,31,33,31,33,30,212,31,172,31,46,31,35,31,177,31,177,30,166,31,166,31,166,30,29,31,168,31,227,31,8,31,17,31,233,31,106,31,106,30,106,29,141,31,55,31,111,31,76,31,76,30,248,31,98,31,98,30,140,31,11,31,248,31,69,31,179,31,31,31,232,31,232,30,232,29,176,31,4,31,231,31,38,31,107,31,212,31,9,31,176,31,228,31,122,31,197,31,197,30,38,31,37,31,228,31,14,31,14,30,208,31,100,31,215,31,158,31,39,31,39,31,201,31,125,31,57,31,244,31,219,31,21,31,144,31,228,31,157,31,10,31,115,31,115,30,201,31,201,30,201,29,201,28,199,31,188,31,134,31,23,31,214,31,214,31,155,31,126,31,227,31,227,30,128,31,189,31,189,30,70,31,25,31,25,30,232,31,232,30,169,31,194,31,137,31,60,31,60,30,89,31,113,31,159,31,203,31,78,31,78,30,78,29,37,31,53,31,167,31,148,31,148,30,150,31,214,31,7,31,212,31,212,30,212,29,104,31,104,30,197,31,175,31,111,31,218,31,83,31,247,31,247,30,217,31,57,31,191,31,138,31,138,30,158,31,46,31,108,31,170,31,57,31,202,31,188,31,111,31,111,30,105,31,168,31,40,31,241,31,110,31,40,31,249,31,162,31,162,30,150,31,136,31,38,31,157,31,182,31,126,31,126,30,92,31,49,31,192,31,254,31,254,31,33,31,70,31,32,31,32,30,49,31,149,31,149,30,254,31,20,31,244,31,234,31,234,30,123,31,123,30,90,31,122,31,122,31,79,31,41,31,98,31,219,31,176,31,151,31,151,30,188,31,111,31,111,30,126,31,227,31,100,31,95,31,46,31,46,30,104,31,187,31,22,31,49,31,100,31,52,31,52,30,15,31,129,31,129,30,60,31,157,31,92,31,48,31,4,31,223,31,189,31,152,31,224,31,224,30,224,29,137,31,137,30,103,31,50,31,169,31,154,31,24,31,27,31,27,30,81,31,120,31,127,31,14,31,89,31,128,31,38,31,38,30,124,31,254,31,39,31,146,31,236,31,80,31,80,30,251,31,251,30,183,31,189,31,189,30,126,31,41,31,212,31,212,30,212,29,212,28,212,27,212,26,50,31,239,31,152,31,152,30,251,31,174,31,19,31,51,31,186,31,153,31,85,31,230,31,80,31,80,30,80,29,106,31,134,31,200,31,214,31,91,31,124,31,204,31,32,31,32,30,203,31,217,31,242,31,170,31,138,31,41,31,94,31,151,31,198,31,104,31,109,31,188,31,109,31,7,31,223,31,138,31,234,31,211,31,129,31,124,31,124,30,124,29,124,28,21,31,164,31,164,30,25,31,25,30,25,29,184,31,184,30,12,31,96,31,199,31,199,30,154,31,157,31,157,30,227,31,207,31,150,31,150,30,40,31,146,31,21,31,71,31,71,30,6,31,17,31,129,31,22,31,22,30,223,31,91,31,3,31,114,31,230,31,141,31,141,30,166,31,49,31,49,30,73,31,70,31,11,31,228,31,146,31,146,30,146,29,103,31,75,31,75,30,101,31,37,31,37,30,230,31,166,31,249,31,92,31,92,30,165,31,20,31,19,31,27,31,27,30,128,31,111,31,111,30,24,31,68,31,68,30,163,31,176,31,55,31,56,31,56,30,92,31,57,31,16,31,39,31,39,30,228,31,228,30,127,31,219,31,47,31,86,31,205,31,115,31,38,31,38,30,220,31,226,31,180,31,75,31,172,31,89,31,40,31,232,31,47,31,39,31,69,31,224,31,4,31,198,31,198,30,239,31,254,31,34,31,218,31,221,31,250,31,100,31,49,31,133,31,3,31,11,31,11,30,248,31,211,31,7,31,76,31,205,31,180,31,180,30,180,29,47,31,181,31,61,31,158,31,158,30,37,31,75,31,238,31,97,31,46,31,68,31,132,31,49,31,61,31,61,30,167,31,28,31,152,31,152,30,128,31,114,31,211,31,120,31,217,31,114,31,114,30,208,31,208,30,26,31,121,31,121,30,181,31,246,31,8,31,8,30,209,31,247,31,166,31,166,30,37,31,123,31,163,31,150,31,33,31,33,30,32,31,138,31,110,31,204,31,79,31,79,30,167,31,183,31,16,31,19,31,69,31,131,31,190,31,190,30,5,31,5,30,163,31,151,31,116,31,44,31,34,31,115,31,115,30,115,29,115,28,115,27,47,31,96,31,199,31,216,31,169,31,185,31,151,31,230,31,100,31,100,30,197,31,197,30,197,29,101,31,99,31,13,31,174,31,95,31,74,31,74,30,243,31,194,31,201,31,222,31,3,31,235,31,119,31,203,31,98,31,233,31,136,31,208,31,34,31,85,31,30,31,179,31,155,31,244,31,200,31,121,31,121,30,146,31,170,31,206,31,78,31,97,31,34,31,20,31,63,31,25,31,182,31,134,31,145,31,163,31,178,31,245,31,29,31,45,31,45,30,229,31,220,31,140,31,118,31,49,31,199,31,247,31,34,31,171,31,114,31,169,31,209,31,105,31,236,31,184,31,180,31,180,30,71,31,41,31,229,31,98,31,197,31,197,30,216,31,219,31,41,31,197,31,49,31,205,31,254,31,27,31,27,30,212,31,105,31,36,31,195,31,232,31,253,31,31,31,189,31,194,31,48,31,234,31,234,30,226,31,238,31,151,31,114,31,114,30,122,31,140,31,55,31,222,31,118,31,255,31,213,31,60,31,13,31,162,31,168,31,20,31,123,31,123,30,83,31,199,31,233,31,193,31,232,31,255,31,224,31,224,30,120,31,223,31,143,31,221,31,221,30,231,31,231,30,187,31,251,31,243,31,27,31,91,31,37,31,24,31,134,31,134,30,115,31,148,31,254,31,144,31,144,30,144,29,155,31,46,31,162,31,129,31,84,31,4,31,247,31,215,31,158,31,185,31,60,31,60,30,75,31,143,31,38,31,38,30,78,31,249,31,249,30,154,31,87,31,254,31,211,31,143,31,181,31,3,31,22,31,108,31,204,31,139,31,74,31,201,31,157,31,23,31,100,31,100,30,203,31,251,31,44,31,52,31,21,31,53,31,53,30,53,29,53,28,85,31,19,31,19,30,254,31,210,31,21,31,62,31,62,30,11,31,227,31,22,31,23,31,23,30,23,29,136,31,108,31,25,31,189,31,189,30,179,31,48,31,48,30,244,31,217,31,9,31,9,30,107,31,153,31,153,30,127,31,207,31,23,31,210,31,202,31,27,31,183,31,198,31,231,31,101,31,146,31,60,31,127,31,9,31,220,31,48,31,134,31,134,30,29,31,28,31,67,31,67,30,183,31,183,30,147,31,124,31,224,31,123,31,221,31,221,30,221,29,185,31,241,31,212,31,40,31,152,31,46,31,77,31,77,30,244,31,244,30,129,31,49,31,49,30,47,31,240,31,51,31,244,31,50,31,5,31,18,31,40,31,40,30,148,31,148,30,235,31,254,31,254,30,152,31,152,30,13,31,110,31,149,31,30,31,249,31,20,31,40,31,140,31,24,31,149,31,196,31,88,31,145,31,145,30,154,31,80,31,88,31,216,31,198,31,211,31,60,31,60,30,175,31,57,31,148,31,148,30,193,31,193,30,193,29,193,31,193,30,193,29,185,31,101,31,114,31,114,30,51,31,123,31,232,31,70,31,179,31,57,31,171,31,171,30,171,29,100,31,246,31,103,31,19,31,19,30,102,31,102,30,102,29,68,31,25,31,48,31,48,30,15,31,76,31,153,31,238,31,238,30,238,29,107,31,22,31,114,31,116,31,170,31,170,30,170,29,170,28,200,31,207,31,181,31,166,31,130,31,16,31,109,31,231,31,198,31,189,31,1,31,217,31,217,30,34,31,91,31,67,31,18,31,162,31,162,30,19,31,152,31,83,31,247,31,173,31,173,30,173,29,220,31,147,31,139,31,139,30,169,31,62,31,227,31,151,31,152,31,88,31,97,31,206,31,123,31,81,31,152,31,152,30,135,31,159,31,159,30,159,29,172,31,193,31,202,31,39,31,39,30,127,31,127,30,116,31,69,31,69,30,102,31,100,31,6,31,159,31,159,30,132,31,153,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
