-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 705;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (162,0,62,0,0,0,0,0,248,0,0,0,243,0,172,0,96,0,16,0,153,0,100,0,180,0,238,0,67,0,156,0,78,0,36,0,250,0,218,0,17,0,189,0,208,0,121,0,75,0,136,0,98,0,184,0,43,0,100,0,4,0,93,0,68,0,0,0,182,0,251,0,49,0,86,0,68,0,146,0,0,0,145,0,66,0,28,0,31,0,175,0,75,0,52,0,163,0,4,0,0,0,0,0,0,0,0,0,0,0,14,0,191,0,111,0,0,0,108,0,200,0,176,0,205,0,174,0,221,0,51,0,196,0,162,0,68,0,6,0,202,0,0,0,233,0,132,0,104,0,0,0,209,0,92,0,181,0,80,0,68,0,108,0,204,0,0,0,0,0,161,0,22,0,58,0,254,0,140,0,198,0,0,0,34,0,209,0,144,0,231,0,0,0,134,0,98,0,166,0,0,0,117,0,237,0,228,0,224,0,249,0,102,0,161,0,26,0,175,0,239,0,0,0,152,0,0,0,51,0,23,0,241,0,62,0,115,0,100,0,0,0,71,0,238,0,241,0,54,0,0,0,178,0,169,0,131,0,197,0,188,0,237,0,15,0,130,0,168,0,39,0,31,0,0,0,38,0,66,0,62,0,253,0,227,0,151,0,219,0,154,0,190,0,179,0,0,0,16,0,29,0,191,0,189,0,107,0,125,0,221,0,0,0,180,0,112,0,52,0,37,0,52,0,172,0,154,0,21,0,0,0,173,0,145,0,173,0,38,0,220,0,0,0,54,0,223,0,77,0,42,0,233,0,54,0,0,0,95,0,156,0,121,0,24,0,146,0,116,0,0,0,129,0,186,0,5,0,0,0,99,0,0,0,202,0,229,0,22,0,0,0,221,0,187,0,23,0,2,0,245,0,0,0,0,0,248,0,217,0,95,0,224,0,0,0,0,0,0,0,0,0,145,0,64,0,176,0,119,0,0,0,139,0,156,0,150,0,220,0,181,0,92,0,91,0,0,0,17,0,95,0,19,0,0,0,209,0,0,0,230,0,136,0,0,0,97,0,187,0,0,0,209,0,151,0,88,0,165,0,176,0,141,0,100,0,163,0,19,0,0,0,150,0,78,0,13,0,194,0,37,0,253,0,15,0,0,0,220,0,86,0,164,0,179,0,14,0,0,0,134,0,229,0,0,0,173,0,115,0,229,0,174,0,229,0,129,0,0,0,62,0,167,0,235,0,192,0,170,0,250,0,97,0,0,0,0,0,0,0,250,0,244,0,138,0,46,0,27,0,33,0,205,0,0,0,223,0,0,0,226,0,220,0,0,0,201,0,166,0,233,0,29,0,74,0,182,0,20,0,253,0,80,0,62,0,28,0,37,0,203,0,90,0,51,0,200,0,31,0,14,0,20,0,149,0,125,0,62,0,28,0,121,0,102,0,159,0,141,0,76,0,0,0,167,0,0,0,0,0,24,0,158,0,24,0,0,0,147,0,71,0,22,0,0,0,0,0,0,0,125,0,101,0,78,0,3,0,14,0,180,0,0,0,209,0,0,0,171,0,136,0,0,0,86,0,0,0,116,0,13,0,8,0,108,0,207,0,128,0,0,0,0,0,214,0,70,0,85,0,161,0,204,0,120,0,213,0,87,0,153,0,98,0,111,0,244,0,91,0,247,0,0,0,164,0,144,0,31,0,103,0,182,0,62,0,152,0,190,0,215,0,11,0,15,0,84,0,239,0,117,0,145,0,0,0,202,0,0,0,0,0,0,0,255,0,56,0,52,0,82,0,0,0,34,0,0,0,211,0,245,0,44,0,10,0,40,0,101,0,18,0,0,0,204,0,8,0,209,0,59,0,84,0,17,0,145,0,231,0,136,0,64,0,0,0,196,0,96,0,248,0,0,0,177,0,58,0,238,0,196,0,22,0,168,0,0,0,181,0,0,0,105,0,167,0,65,0,0,0,0,0,115,0,0,0,0,0,249,0,34,0,20,0,41,0,248,0,138,0,3,0,78,0,84,0,244,0,109,0,241,0,231,0,254,0,106,0,113,0,252,0,0,0,60,0,212,0,69,0,0,0,215,0,154,0,218,0,92,0,20,0,133,0,16,0,242,0,175,0,75,0,220,0,215,0,0,0,13,0,21,0,87,0,57,0,198,0,44,0,180,0,98,0,0,0,130,0,60,0,158,0,8,0,249,0,0,0,158,0,0,0,3,0,0,0,0,0,51,0,170,0,0,0,0,0,237,0,0,0,214,0,0,0,142,0,173,0,202,0,246,0,0,0,0,0,195,0,0,0,141,0,0,0,169,0,241,0,71,0,141,0,0,0,0,0,236,0,7,0,38,0,0,0,148,0,8,0,44,0,182,0,163,0,0,0,1,0,128,0,3,0,169,0,0,0,0,0,68,0,4,0,0,0,113,0,0,0,119,0,163,0,139,0,42,0,196,0,0,0,148,0,190,0,0,0,0,0,4,0,133,0,171,0,83,0,167,0,128,0,69,0,163,0,164,0,204,0,200,0,208,0,253,0,138,0,83,0,39,0,72,0,0,0,252,0,0,0,187,0,0,0,0,0,71,0,144,0,199,0,0,0,12,0,137,0,0,0,89,0,107,0,35,0,180,0,141,0,0,0,206,0,42,0,159,0,152,0,230,0,122,0,0,0,0,0,217,0,113,0,123,0,195,0,100,0,0,0,0,0,228,0,199,0,71,0,57,0,196,0,70,0,255,0,192,0,11,0,127,0,249,0,183,0,10,0,93,0,81,0,133,0,213,0,0,0,0,0,186,0,44,0,47,0,44,0,2,0,169,0,0,0,64,0,89,0,13,0,0,0,0,0,195,0,0,0,99,0,29,0,162,0,149,0,199,0,154,0,144,0,0,0,111,0,0,0,68,0,0,0,0,0,142,0,0,0,2,0,229,0,0,0,22,0,183,0,37,0,85,0,107,0,92,0,0,0,134,0,0,0,0,0,9,0,51,0,111,0,166,0,0,0,0,0,0,0,138,0,48,0,190,0,76,0,66,0,223,0,72,0,131,0,255,0,112,0,133,0,156,0,244,0,46,0,210,0,136,0,213,0,216,0,177,0,24,0,209,0,0,0,82,0,214,0,232,0,0,0,221,0,0,0,211,0,89,0,0,0,0,0,11,0,238,0,0,0,113,0,172,0);
signal scenario_full  : scenario_type := (162,31,62,31,62,30,62,29,248,31,248,30,243,31,172,31,96,31,16,31,153,31,100,31,180,31,238,31,67,31,156,31,78,31,36,31,250,31,218,31,17,31,189,31,208,31,121,31,75,31,136,31,98,31,184,31,43,31,100,31,4,31,93,31,68,31,68,30,182,31,251,31,49,31,86,31,68,31,146,31,146,30,145,31,66,31,28,31,31,31,175,31,75,31,52,31,163,31,4,31,4,30,4,29,4,28,4,27,4,26,14,31,191,31,111,31,111,30,108,31,200,31,176,31,205,31,174,31,221,31,51,31,196,31,162,31,68,31,6,31,202,31,202,30,233,31,132,31,104,31,104,30,209,31,92,31,181,31,80,31,68,31,108,31,204,31,204,30,204,29,161,31,22,31,58,31,254,31,140,31,198,31,198,30,34,31,209,31,144,31,231,31,231,30,134,31,98,31,166,31,166,30,117,31,237,31,228,31,224,31,249,31,102,31,161,31,26,31,175,31,239,31,239,30,152,31,152,30,51,31,23,31,241,31,62,31,115,31,100,31,100,30,71,31,238,31,241,31,54,31,54,30,178,31,169,31,131,31,197,31,188,31,237,31,15,31,130,31,168,31,39,31,31,31,31,30,38,31,66,31,62,31,253,31,227,31,151,31,219,31,154,31,190,31,179,31,179,30,16,31,29,31,191,31,189,31,107,31,125,31,221,31,221,30,180,31,112,31,52,31,37,31,52,31,172,31,154,31,21,31,21,30,173,31,145,31,173,31,38,31,220,31,220,30,54,31,223,31,77,31,42,31,233,31,54,31,54,30,95,31,156,31,121,31,24,31,146,31,116,31,116,30,129,31,186,31,5,31,5,30,99,31,99,30,202,31,229,31,22,31,22,30,221,31,187,31,23,31,2,31,245,31,245,30,245,29,248,31,217,31,95,31,224,31,224,30,224,29,224,28,224,27,145,31,64,31,176,31,119,31,119,30,139,31,156,31,150,31,220,31,181,31,92,31,91,31,91,30,17,31,95,31,19,31,19,30,209,31,209,30,230,31,136,31,136,30,97,31,187,31,187,30,209,31,151,31,88,31,165,31,176,31,141,31,100,31,163,31,19,31,19,30,150,31,78,31,13,31,194,31,37,31,253,31,15,31,15,30,220,31,86,31,164,31,179,31,14,31,14,30,134,31,229,31,229,30,173,31,115,31,229,31,174,31,229,31,129,31,129,30,62,31,167,31,235,31,192,31,170,31,250,31,97,31,97,30,97,29,97,28,250,31,244,31,138,31,46,31,27,31,33,31,205,31,205,30,223,31,223,30,226,31,220,31,220,30,201,31,166,31,233,31,29,31,74,31,182,31,20,31,253,31,80,31,62,31,28,31,37,31,203,31,90,31,51,31,200,31,31,31,14,31,20,31,149,31,125,31,62,31,28,31,121,31,102,31,159,31,141,31,76,31,76,30,167,31,167,30,167,29,24,31,158,31,24,31,24,30,147,31,71,31,22,31,22,30,22,29,22,28,125,31,101,31,78,31,3,31,14,31,180,31,180,30,209,31,209,30,171,31,136,31,136,30,86,31,86,30,116,31,13,31,8,31,108,31,207,31,128,31,128,30,128,29,214,31,70,31,85,31,161,31,204,31,120,31,213,31,87,31,153,31,98,31,111,31,244,31,91,31,247,31,247,30,164,31,144,31,31,31,103,31,182,31,62,31,152,31,190,31,215,31,11,31,15,31,84,31,239,31,117,31,145,31,145,30,202,31,202,30,202,29,202,28,255,31,56,31,52,31,82,31,82,30,34,31,34,30,211,31,245,31,44,31,10,31,40,31,101,31,18,31,18,30,204,31,8,31,209,31,59,31,84,31,17,31,145,31,231,31,136,31,64,31,64,30,196,31,96,31,248,31,248,30,177,31,58,31,238,31,196,31,22,31,168,31,168,30,181,31,181,30,105,31,167,31,65,31,65,30,65,29,115,31,115,30,115,29,249,31,34,31,20,31,41,31,248,31,138,31,3,31,78,31,84,31,244,31,109,31,241,31,231,31,254,31,106,31,113,31,252,31,252,30,60,31,212,31,69,31,69,30,215,31,154,31,218,31,92,31,20,31,133,31,16,31,242,31,175,31,75,31,220,31,215,31,215,30,13,31,21,31,87,31,57,31,198,31,44,31,180,31,98,31,98,30,130,31,60,31,158,31,8,31,249,31,249,30,158,31,158,30,3,31,3,30,3,29,51,31,170,31,170,30,170,29,237,31,237,30,214,31,214,30,142,31,173,31,202,31,246,31,246,30,246,29,195,31,195,30,141,31,141,30,169,31,241,31,71,31,141,31,141,30,141,29,236,31,7,31,38,31,38,30,148,31,8,31,44,31,182,31,163,31,163,30,1,31,128,31,3,31,169,31,169,30,169,29,68,31,4,31,4,30,113,31,113,30,119,31,163,31,139,31,42,31,196,31,196,30,148,31,190,31,190,30,190,29,4,31,133,31,171,31,83,31,167,31,128,31,69,31,163,31,164,31,204,31,200,31,208,31,253,31,138,31,83,31,39,31,72,31,72,30,252,31,252,30,187,31,187,30,187,29,71,31,144,31,199,31,199,30,12,31,137,31,137,30,89,31,107,31,35,31,180,31,141,31,141,30,206,31,42,31,159,31,152,31,230,31,122,31,122,30,122,29,217,31,113,31,123,31,195,31,100,31,100,30,100,29,228,31,199,31,71,31,57,31,196,31,70,31,255,31,192,31,11,31,127,31,249,31,183,31,10,31,93,31,81,31,133,31,213,31,213,30,213,29,186,31,44,31,47,31,44,31,2,31,169,31,169,30,64,31,89,31,13,31,13,30,13,29,195,31,195,30,99,31,29,31,162,31,149,31,199,31,154,31,144,31,144,30,111,31,111,30,68,31,68,30,68,29,142,31,142,30,2,31,229,31,229,30,22,31,183,31,37,31,85,31,107,31,92,31,92,30,134,31,134,30,134,29,9,31,51,31,111,31,166,31,166,30,166,29,166,28,138,31,48,31,190,31,76,31,66,31,223,31,72,31,131,31,255,31,112,31,133,31,156,31,244,31,46,31,210,31,136,31,213,31,216,31,177,31,24,31,209,31,209,30,82,31,214,31,232,31,232,30,221,31,221,30,211,31,89,31,89,30,89,29,11,31,238,31,238,30,113,31,172,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
