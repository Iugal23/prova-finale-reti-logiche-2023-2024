-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 362;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,143,0,0,0,0,0,0,0,27,0,13,0,184,0,231,0,0,0,0,0,244,0,14,0,119,0,93,0,216,0,0,0,217,0,106,0,74,0,16,0,31,0,139,0,39,0,237,0,0,0,156,0,139,0,41,0,229,0,240,0,87,0,89,0,64,0,79,0,118,0,0,0,0,0,111,0,174,0,32,0,158,0,245,0,229,0,172,0,165,0,194,0,62,0,94,0,49,0,47,0,216,0,20,0,90,0,232,0,238,0,50,0,192,0,115,0,203,0,44,0,129,0,15,0,8,0,0,0,0,0,222,0,99,0,0,0,0,0,0,0,0,0,125,0,0,0,67,0,183,0,128,0,244,0,74,0,93,0,6,0,0,0,34,0,0,0,164,0,172,0,46,0,120,0,231,0,157,0,0,0,0,0,228,0,133,0,83,0,231,0,67,0,180,0,35,0,198,0,46,0,0,0,248,0,201,0,3,0,207,0,42,0,166,0,100,0,173,0,231,0,186,0,0,0,149,0,0,0,0,0,200,0,107,0,254,0,96,0,211,0,0,0,165,0,185,0,185,0,125,0,44,0,107,0,119,0,220,0,120,0,211,0,204,0,57,0,0,0,95,0,1,0,225,0,178,0,248,0,74,0,2,0,9,0,144,0,63,0,111,0,164,0,77,0,0,0,15,0,0,0,173,0,237,0,85,0,208,0,35,0,3,0,247,0,0,0,75,0,50,0,43,0,182,0,201,0,31,0,177,0,174,0,158,0,31,0,96,0,120,0,0,0,146,0,21,0,47,0,252,0,0,0,0,0,120,0,0,0,0,0,0,0,27,0,201,0,56,0,64,0,160,0,134,0,86,0,119,0,0,0,120,0,0,0,23,0,0,0,0,0,0,0,13,0,205,0,225,0,157,0,0,0,0,0,201,0,239,0,0,0,237,0,0,0,82,0,113,0,94,0,212,0,18,0,0,0,55,0,0,0,0,0,96,0,68,0,126,0,102,0,64,0,111,0,241,0,0,0,251,0,4,0,208,0,174,0,9,0,146,0,136,0,0,0,62,0,154,0,0,0,211,0,0,0,0,0,0,0,136,0,51,0,19,0,108,0,35,0,141,0,19,0,0,0,18,0,196,0,247,0,0,0,45,0,144,0,114,0,62,0,26,0,14,0,16,0,131,0,230,0,17,0,115,0,58,0,5,0,126,0,218,0,232,0,0,0,157,0,147,0,179,0,0,0,79,0,95,0,58,0,153,0,0,0,85,0,130,0,172,0,167,0,167,0,183,0,32,0,240,0,104,0,158,0,0,0,222,0,254,0,227,0,15,0,177,0,0,0,106,0,59,0,142,0,0,0,0,0,91,0,29,0,52,0,0,0,173,0,107,0,84,0,69,0,244,0,0,0,0,0,26,0,251,0,0,0,84,0,181,0,60,0,0,0,185,0,119,0,34,0,44,0,0,0,73,0,132,0,91,0,8,0,86,0,30,0,241,0,0,0,92,0,23,0,0,0,203,0,120,0,0,0,131,0,29,0,144,0,66,0,179,0,193,0,45,0,0,0,220,0,221,0,72,0,207,0,0,0,46,0,204,0,197,0,128,0,47,0,0,0,0,0,149,0,73,0,0,0,42,0,115,0);
signal scenario_full  : scenario_type := (0,0,143,31,143,30,143,29,143,28,27,31,13,31,184,31,231,31,231,30,231,29,244,31,14,31,119,31,93,31,216,31,216,30,217,31,106,31,74,31,16,31,31,31,139,31,39,31,237,31,237,30,156,31,139,31,41,31,229,31,240,31,87,31,89,31,64,31,79,31,118,31,118,30,118,29,111,31,174,31,32,31,158,31,245,31,229,31,172,31,165,31,194,31,62,31,94,31,49,31,47,31,216,31,20,31,90,31,232,31,238,31,50,31,192,31,115,31,203,31,44,31,129,31,15,31,8,31,8,30,8,29,222,31,99,31,99,30,99,29,99,28,99,27,125,31,125,30,67,31,183,31,128,31,244,31,74,31,93,31,6,31,6,30,34,31,34,30,164,31,172,31,46,31,120,31,231,31,157,31,157,30,157,29,228,31,133,31,83,31,231,31,67,31,180,31,35,31,198,31,46,31,46,30,248,31,201,31,3,31,207,31,42,31,166,31,100,31,173,31,231,31,186,31,186,30,149,31,149,30,149,29,200,31,107,31,254,31,96,31,211,31,211,30,165,31,185,31,185,31,125,31,44,31,107,31,119,31,220,31,120,31,211,31,204,31,57,31,57,30,95,31,1,31,225,31,178,31,248,31,74,31,2,31,9,31,144,31,63,31,111,31,164,31,77,31,77,30,15,31,15,30,173,31,237,31,85,31,208,31,35,31,3,31,247,31,247,30,75,31,50,31,43,31,182,31,201,31,31,31,177,31,174,31,158,31,31,31,96,31,120,31,120,30,146,31,21,31,47,31,252,31,252,30,252,29,120,31,120,30,120,29,120,28,27,31,201,31,56,31,64,31,160,31,134,31,86,31,119,31,119,30,120,31,120,30,23,31,23,30,23,29,23,28,13,31,205,31,225,31,157,31,157,30,157,29,201,31,239,31,239,30,237,31,237,30,82,31,113,31,94,31,212,31,18,31,18,30,55,31,55,30,55,29,96,31,68,31,126,31,102,31,64,31,111,31,241,31,241,30,251,31,4,31,208,31,174,31,9,31,146,31,136,31,136,30,62,31,154,31,154,30,211,31,211,30,211,29,211,28,136,31,51,31,19,31,108,31,35,31,141,31,19,31,19,30,18,31,196,31,247,31,247,30,45,31,144,31,114,31,62,31,26,31,14,31,16,31,131,31,230,31,17,31,115,31,58,31,5,31,126,31,218,31,232,31,232,30,157,31,147,31,179,31,179,30,79,31,95,31,58,31,153,31,153,30,85,31,130,31,172,31,167,31,167,31,183,31,32,31,240,31,104,31,158,31,158,30,222,31,254,31,227,31,15,31,177,31,177,30,106,31,59,31,142,31,142,30,142,29,91,31,29,31,52,31,52,30,173,31,107,31,84,31,69,31,244,31,244,30,244,29,26,31,251,31,251,30,84,31,181,31,60,31,60,30,185,31,119,31,34,31,44,31,44,30,73,31,132,31,91,31,8,31,86,31,30,31,241,31,241,30,92,31,23,31,23,30,203,31,120,31,120,30,131,31,29,31,144,31,66,31,179,31,193,31,45,31,45,30,220,31,221,31,72,31,207,31,207,30,46,31,204,31,197,31,128,31,47,31,47,30,47,29,149,31,73,31,73,30,42,31,115,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
