-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_214 is
end project_tb_214;

architecture project_tb_arch_214 of project_tb_214 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 457;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,182,0,188,0,141,0,0,0,246,0,150,0,58,0,0,0,74,0,224,0,0,0,113,0,0,0,145,0,220,0,210,0,228,0,0,0,0,0,97,0,210,0,42,0,129,0,0,0,138,0,218,0,127,0,129,0,0,0,179,0,214,0,222,0,0,0,237,0,217,0,121,0,0,0,220,0,209,0,109,0,147,0,8,0,131,0,0,0,0,0,186,0,245,0,90,0,37,0,67,0,226,0,147,0,154,0,53,0,20,0,0,0,243,0,189,0,100,0,247,0,162,0,0,0,122,0,28,0,13,0,215,0,118,0,0,0,14,0,98,0,128,0,152,0,0,0,252,0,149,0,57,0,247,0,0,0,18,0,252,0,67,0,0,0,103,0,255,0,201,0,35,0,148,0,143,0,148,0,0,0,0,0,137,0,186,0,0,0,202,0,0,0,201,0,185,0,33,0,176,0,240,0,32,0,10,0,0,0,246,0,101,0,141,0,0,0,177,0,169,0,165,0,90,0,209,0,247,0,104,0,244,0,164,0,120,0,249,0,186,0,249,0,186,0,0,0,228,0,26,0,102,0,0,0,152,0,150,0,182,0,239,0,236,0,234,0,0,0,186,0,60,0,0,0,0,0,72,0,22,0,8,0,110,0,66,0,74,0,160,0,11,0,55,0,25,0,0,0,9,0,0,0,179,0,0,0,11,0,240,0,46,0,226,0,107,0,187,0,103,0,0,0,104,0,27,0,45,0,245,0,255,0,209,0,0,0,173,0,239,0,102,0,50,0,56,0,0,0,0,0,242,0,0,0,75,0,26,0,172,0,0,0,43,0,132,0,38,0,148,0,0,0,144,0,171,0,0,0,121,0,136,0,139,0,0,0,0,0,177,0,111,0,38,0,98,0,145,0,80,0,0,0,0,0,93,0,0,0,13,0,64,0,165,0,110,0,14,0,0,0,0,0,73,0,179,0,155,0,38,0,178,0,42,0,121,0,0,0,165,0,74,0,0,0,151,0,70,0,198,0,0,0,26,0,0,0,186,0,0,0,219,0,165,0,0,0,0,0,196,0,0,0,102,0,215,0,29,0,35,0,100,0,30,0,92,0,0,0,188,0,227,0,228,0,0,0,42,0,0,0,0,0,89,0,226,0,0,0,214,0,219,0,222,0,91,0,0,0,230,0,9,0,66,0,0,0,184,0,188,0,0,0,213,0,0,0,0,0,202,0,21,0,124,0,254,0,15,0,216,0,90,0,233,0,0,0,44,0,14,0,110,0,65,0,0,0,97,0,0,0,152,0,172,0,222,0,140,0,60,0,240,0,115,0,65,0,35,0,125,0,139,0,221,0,19,0,181,0,0,0,0,0,0,0,0,0,215,0,90,0,193,0,128,0,14,0,0,0,185,0,0,0,0,0,115,0,0,0,158,0,130,0,214,0,123,0,56,0,0,0,142,0,0,0,200,0,236,0,251,0,0,0,0,0,61,0,46,0,0,0,237,0,138,0,0,0,0,0,40,0,0,0,0,0,134,0,24,0,215,0,72,0,7,0,184,0,31,0,177,0,169,0,137,0,0,0,0,0,0,0,163,0,0,0,6,0,85,0,165,0,211,0,155,0,86,0,73,0,222,0,0,0,11,0,124,0,198,0,0,0,52,0,114,0,27,0,174,0,237,0,0,0,0,0,166,0,0,0,26,0,109,0,0,0,165,0,199,0,74,0,99,0,0,0,233,0,158,0,88,0,172,0,0,0,145,0,0,0,96,0,220,0,0,0,45,0,90,0,17,0,170,0,239,0,0,0,194,0,236,0,0,0,233,0,103,0,42,0,23,0,0,0,251,0,5,0,131,0,170,0,238,0,78,0,46,0,128,0,160,0,13,0,241,0,87,0,81,0,166,0,170,0,0,0,0,0,143,0,202,0,5,0,0,0,0,0,17,0,237,0,166,0,106,0,142,0,142,0,149,0,0,0,0,0,0,0,0,0,120,0,83,0,40,0,30,0,21,0,0,0,120,0,47,0,175,0,0,0,143,0,181,0,178,0,66,0,150,0,26,0,20,0);
signal scenario_full  : scenario_type := (0,0,182,31,188,31,141,31,141,30,246,31,150,31,58,31,58,30,74,31,224,31,224,30,113,31,113,30,145,31,220,31,210,31,228,31,228,30,228,29,97,31,210,31,42,31,129,31,129,30,138,31,218,31,127,31,129,31,129,30,179,31,214,31,222,31,222,30,237,31,217,31,121,31,121,30,220,31,209,31,109,31,147,31,8,31,131,31,131,30,131,29,186,31,245,31,90,31,37,31,67,31,226,31,147,31,154,31,53,31,20,31,20,30,243,31,189,31,100,31,247,31,162,31,162,30,122,31,28,31,13,31,215,31,118,31,118,30,14,31,98,31,128,31,152,31,152,30,252,31,149,31,57,31,247,31,247,30,18,31,252,31,67,31,67,30,103,31,255,31,201,31,35,31,148,31,143,31,148,31,148,30,148,29,137,31,186,31,186,30,202,31,202,30,201,31,185,31,33,31,176,31,240,31,32,31,10,31,10,30,246,31,101,31,141,31,141,30,177,31,169,31,165,31,90,31,209,31,247,31,104,31,244,31,164,31,120,31,249,31,186,31,249,31,186,31,186,30,228,31,26,31,102,31,102,30,152,31,150,31,182,31,239,31,236,31,234,31,234,30,186,31,60,31,60,30,60,29,72,31,22,31,8,31,110,31,66,31,74,31,160,31,11,31,55,31,25,31,25,30,9,31,9,30,179,31,179,30,11,31,240,31,46,31,226,31,107,31,187,31,103,31,103,30,104,31,27,31,45,31,245,31,255,31,209,31,209,30,173,31,239,31,102,31,50,31,56,31,56,30,56,29,242,31,242,30,75,31,26,31,172,31,172,30,43,31,132,31,38,31,148,31,148,30,144,31,171,31,171,30,121,31,136,31,139,31,139,30,139,29,177,31,111,31,38,31,98,31,145,31,80,31,80,30,80,29,93,31,93,30,13,31,64,31,165,31,110,31,14,31,14,30,14,29,73,31,179,31,155,31,38,31,178,31,42,31,121,31,121,30,165,31,74,31,74,30,151,31,70,31,198,31,198,30,26,31,26,30,186,31,186,30,219,31,165,31,165,30,165,29,196,31,196,30,102,31,215,31,29,31,35,31,100,31,30,31,92,31,92,30,188,31,227,31,228,31,228,30,42,31,42,30,42,29,89,31,226,31,226,30,214,31,219,31,222,31,91,31,91,30,230,31,9,31,66,31,66,30,184,31,188,31,188,30,213,31,213,30,213,29,202,31,21,31,124,31,254,31,15,31,216,31,90,31,233,31,233,30,44,31,14,31,110,31,65,31,65,30,97,31,97,30,152,31,172,31,222,31,140,31,60,31,240,31,115,31,65,31,35,31,125,31,139,31,221,31,19,31,181,31,181,30,181,29,181,28,181,27,215,31,90,31,193,31,128,31,14,31,14,30,185,31,185,30,185,29,115,31,115,30,158,31,130,31,214,31,123,31,56,31,56,30,142,31,142,30,200,31,236,31,251,31,251,30,251,29,61,31,46,31,46,30,237,31,138,31,138,30,138,29,40,31,40,30,40,29,134,31,24,31,215,31,72,31,7,31,184,31,31,31,177,31,169,31,137,31,137,30,137,29,137,28,163,31,163,30,6,31,85,31,165,31,211,31,155,31,86,31,73,31,222,31,222,30,11,31,124,31,198,31,198,30,52,31,114,31,27,31,174,31,237,31,237,30,237,29,166,31,166,30,26,31,109,31,109,30,165,31,199,31,74,31,99,31,99,30,233,31,158,31,88,31,172,31,172,30,145,31,145,30,96,31,220,31,220,30,45,31,90,31,17,31,170,31,239,31,239,30,194,31,236,31,236,30,233,31,103,31,42,31,23,31,23,30,251,31,5,31,131,31,170,31,238,31,78,31,46,31,128,31,160,31,13,31,241,31,87,31,81,31,166,31,170,31,170,30,170,29,143,31,202,31,5,31,5,30,5,29,17,31,237,31,166,31,106,31,142,31,142,31,149,31,149,30,149,29,149,28,149,27,120,31,83,31,40,31,30,31,21,31,21,30,120,31,47,31,175,31,175,30,143,31,181,31,178,31,66,31,150,31,26,31,20,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
