-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 958;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (127,0,230,0,207,0,34,0,53,0,82,0,156,0,204,0,0,0,249,0,129,0,18,0,85,0,0,0,172,0,200,0,0,0,79,0,0,0,0,0,52,0,244,0,0,0,82,0,0,0,238,0,142,0,39,0,32,0,235,0,46,0,110,0,0,0,240,0,99,0,197,0,46,0,224,0,198,0,213,0,0,0,0,0,96,0,14,0,104,0,178,0,0,0,152,0,11,0,179,0,84,0,44,0,180,0,0,0,0,0,0,0,153,0,0,0,171,0,32,0,157,0,14,0,0,0,129,0,0,0,0,0,24,0,159,0,217,0,241,0,98,0,56,0,32,0,0,0,53,0,67,0,208,0,87,0,236,0,49,0,181,0,0,0,121,0,118,0,164,0,213,0,77,0,188,0,221,0,181,0,77,0,74,0,0,0,0,0,123,0,76,0,241,0,182,0,71,0,0,0,167,0,126,0,46,0,64,0,91,0,82,0,0,0,107,0,56,0,106,0,103,0,38,0,219,0,184,0,231,0,232,0,94,0,0,0,74,0,121,0,14,0,193,0,173,0,99,0,192,0,244,0,112,0,151,0,233,0,0,0,116,0,209,0,0,0,171,0,217,0,0,0,192,0,8,0,0,0,188,0,210,0,86,0,146,0,27,0,190,0,201,0,0,0,31,0,179,0,168,0,27,0,86,0,184,0,1,0,230,0,220,0,147,0,173,0,22,0,153,0,187,0,0,0,188,0,188,0,35,0,58,0,115,0,122,0,197,0,9,0,117,0,210,0,49,0,80,0,218,0,148,0,144,0,231,0,0,0,165,0,26,0,0,0,80,0,205,0,156,0,111,0,1,0,0,0,130,0,0,0,53,0,141,0,185,0,20,0,195,0,248,0,216,0,86,0,0,0,14,0,157,0,164,0,60,0,141,0,86,0,214,0,131,0,0,0,76,0,229,0,0,0,5,0,25,0,180,0,0,0,0,0,218,0,0,0,147,0,0,0,75,0,131,0,187,0,252,0,173,0,0,0,117,0,137,0,0,0,213,0,113,0,184,0,170,0,171,0,212,0,103,0,202,0,251,0,0,0,60,0,181,0,193,0,118,0,95,0,19,0,249,0,149,0,229,0,53,0,99,0,245,0,94,0,209,0,95,0,0,0,0,0,0,0,97,0,37,0,0,0,105,0,0,0,77,0,31,0,93,0,179,0,136,0,149,0,73,0,61,0,249,0,172,0,0,0,35,0,27,0,211,0,0,0,2,0,74,0,3,0,65,0,48,0,91,0,207,0,46,0,60,0,0,0,65,0,45,0,194,0,29,0,23,0,0,0,171,0,151,0,140,0,192,0,0,0,4,0,0,0,3,0,0,0,0,0,130,0,0,0,105,0,174,0,0,0,0,0,128,0,53,0,0,0,0,0,243,0,6,0,178,0,153,0,163,0,220,0,14,0,0,0,173,0,117,0,145,0,208,0,0,0,180,0,226,0,174,0,0,0,254,0,0,0,0,0,164,0,49,0,188,0,105,0,76,0,236,0,0,0,244,0,0,0,0,0,8,0,171,0,27,0,188,0,146,0,67,0,94,0,0,0,240,0,0,0,191,0,196,0,253,0,116,0,249,0,171,0,0,0,178,0,122,0,0,0,148,0,0,0,0,0,158,0,0,0,190,0,0,0,20,0,147,0,165,0,225,0,191,0,214,0,188,0,234,0,80,0,173,0,47,0,36,0,212,0,34,0,1,0,176,0,0,0,125,0,11,0,244,0,0,0,73,0,201,0,119,0,48,0,161,0,237,0,21,0,0,0,186,0,121,0,0,0,26,0,215,0,31,0,128,0,167,0,231,0,0,0,8,0,8,0,114,0,0,0,127,0,178,0,74,0,200,0,95,0,241,0,0,0,221,0,86,0,106,0,17,0,192,0,229,0,233,0,208,0,117,0,85,0,143,0,0,0,159,0,0,0,119,0,0,0,50,0,18,0,156,0,225,0,65,0,0,0,108,0,53,0,100,0,114,0,70,0,141,0,147,0,128,0,0,0,131,0,0,0,195,0,208,0,210,0,226,0,116,0,195,0,0,0,207,0,0,0,15,0,106,0,81,0,0,0,161,0,90,0,0,0,56,0,73,0,173,0,160,0,36,0,138,0,188,0,22,0,0,0,181,0,201,0,125,0,132,0,0,0,128,0,136,0,198,0,99,0,151,0,0,0,207,0,0,0,0,0,0,0,220,0,183,0,0,0,92,0,106,0,101,0,241,0,161,0,115,0,204,0,0,0,0,0,84,0,130,0,116,0,218,0,59,0,4,0,214,0,181,0,105,0,102,0,202,0,18,0,164,0,129,0,0,0,125,0,107,0,0,0,0,0,226,0,0,0,114,0,191,0,43,0,192,0,30,0,218,0,62,0,70,0,76,0,0,0,73,0,99,0,38,0,179,0,0,0,161,0,182,0,97,0,148,0,238,0,108,0,55,0,216,0,0,0,0,0,193,0,238,0,227,0,234,0,37,0,1,0,0,0,149,0,138,0,250,0,208,0,7,0,105,0,6,0,185,0,71,0,208,0,39,0,0,0,25,0,0,0,0,0,38,0,101,0,8,0,137,0,231,0,0,0,136,0,136,0,42,0,0,0,119,0,17,0,218,0,22,0,24,0,65,0,30,0,0,0,0,0,174,0,52,0,218,0,170,0,205,0,0,0,0,0,109,0,220,0,0,0,168,0,82,0,98,0,20,0,0,0,0,0,88,0,154,0,125,0,181,0,0,0,87,0,11,0,0,0,133,0,65,0,55,0,0,0,27,0,114,0,128,0,200,0,155,0,79,0,0,0,251,0,0,0,90,0,177,0,82,0,218,0,43,0,27,0,142,0,195,0,60,0,45,0,174,0,87,0,249,0,169,0,101,0,32,0,251,0,0,0,216,0,0,0,28,0,0,0,22,0,215,0,121,0,156,0,109,0,177,0,90,0,122,0,40,0,90,0,0,0,0,0,184,0,104,0,20,0,219,0,0,0,19,0,31,0,19,0,108,0,0,0,218,0,149,0,230,0,0,0,200,0,154,0,95,0,170,0,58,0,5,0,226,0,128,0,54,0,113,0,59,0,49,0,217,0,135,0,245,0,0,0,0,0,0,0,0,0,254,0,95,0,64,0,20,0,145,0,213,0,46,0,64,0,93,0,194,0,29,0,208,0,0,0,176,0,0,0,0,0,236,0,172,0,20,0,151,0,254,0,47,0,133,0,0,0,75,0,28,0,127,0,29,0,16,0,131,0,5,0,124,0,196,0,22,0,0,0,217,0,146,0,192,0,0,0,40,0,16,0,43,0,45,0,240,0,0,0,51,0,240,0,17,0,0,0,20,0,41,0,224,0,88,0,230,0,0,0,83,0,10,0,175,0,0,0,186,0,230,0,222,0,183,0,255,0,255,0,210,0,89,0,0,0,240,0,251,0,0,0,0,0,172,0,11,0,149,0,83,0,0,0,131,0,0,0,242,0,0,0,0,0,201,0,0,0,0,0,190,0,12,0,192,0,114,0,129,0,212,0,212,0,5,0,0,0,96,0,51,0,0,0,33,0,0,0,0,0,32,0,213,0,166,0,125,0,0,0,134,0,61,0,75,0,81,0,0,0,157,0,212,0,0,0,74,0,0,0,164,0,31,0,0,0,0,0,0,0,164,0,141,0,78,0,0,0,0,0,62,0,0,0,221,0,0,0,63,0,0,0,0,0,223,0,205,0,175,0,0,0,0,0,106,0,86,0,178,0,12,0,0,0,0,0,164,0,0,0,117,0,221,0,0,0,90,0,70,0,240,0,65,0,54,0,73,0,56,0,0,0,230,0,176,0,252,0,252,0,217,0,19,0,118,0,103,0,237,0,174,0,162,0,0,0,61,0,123,0,13,0,205,0,0,0,112,0,0,0,135,0,11,0,124,0,66,0,243,0,70,0,68,0,101,0,41,0,107,0,129,0,10,0,129,0,33,0,18,0,131,0,0,0,219,0,48,0,206,0,152,0,11,0,77,0,228,0,171,0,99,0,0,0,241,0,0,0,118,0,133,0,7,0,0,0,0,0,82,0,168,0,196,0,112,0,15,0,139,0,0,0,11,0,112,0,115,0,186,0,24,0,120,0,0,0,53,0,9,0,91,0,86,0,133,0,0,0,0,0,82,0,93,0,90,0,45,0,136,0,179,0,17,0,145,0,205,0,160,0,0,0,118,0,110,0,217,0,26,0,171,0,104,0,253,0,207,0,57,0,220,0,171,0,6,0,0,0,96,0,98,0,0,0,8,0,156,0,247,0,17,0,244,0);
signal scenario_full  : scenario_type := (127,31,230,31,207,31,34,31,53,31,82,31,156,31,204,31,204,30,249,31,129,31,18,31,85,31,85,30,172,31,200,31,200,30,79,31,79,30,79,29,52,31,244,31,244,30,82,31,82,30,238,31,142,31,39,31,32,31,235,31,46,31,110,31,110,30,240,31,99,31,197,31,46,31,224,31,198,31,213,31,213,30,213,29,96,31,14,31,104,31,178,31,178,30,152,31,11,31,179,31,84,31,44,31,180,31,180,30,180,29,180,28,153,31,153,30,171,31,32,31,157,31,14,31,14,30,129,31,129,30,129,29,24,31,159,31,217,31,241,31,98,31,56,31,32,31,32,30,53,31,67,31,208,31,87,31,236,31,49,31,181,31,181,30,121,31,118,31,164,31,213,31,77,31,188,31,221,31,181,31,77,31,74,31,74,30,74,29,123,31,76,31,241,31,182,31,71,31,71,30,167,31,126,31,46,31,64,31,91,31,82,31,82,30,107,31,56,31,106,31,103,31,38,31,219,31,184,31,231,31,232,31,94,31,94,30,74,31,121,31,14,31,193,31,173,31,99,31,192,31,244,31,112,31,151,31,233,31,233,30,116,31,209,31,209,30,171,31,217,31,217,30,192,31,8,31,8,30,188,31,210,31,86,31,146,31,27,31,190,31,201,31,201,30,31,31,179,31,168,31,27,31,86,31,184,31,1,31,230,31,220,31,147,31,173,31,22,31,153,31,187,31,187,30,188,31,188,31,35,31,58,31,115,31,122,31,197,31,9,31,117,31,210,31,49,31,80,31,218,31,148,31,144,31,231,31,231,30,165,31,26,31,26,30,80,31,205,31,156,31,111,31,1,31,1,30,130,31,130,30,53,31,141,31,185,31,20,31,195,31,248,31,216,31,86,31,86,30,14,31,157,31,164,31,60,31,141,31,86,31,214,31,131,31,131,30,76,31,229,31,229,30,5,31,25,31,180,31,180,30,180,29,218,31,218,30,147,31,147,30,75,31,131,31,187,31,252,31,173,31,173,30,117,31,137,31,137,30,213,31,113,31,184,31,170,31,171,31,212,31,103,31,202,31,251,31,251,30,60,31,181,31,193,31,118,31,95,31,19,31,249,31,149,31,229,31,53,31,99,31,245,31,94,31,209,31,95,31,95,30,95,29,95,28,97,31,37,31,37,30,105,31,105,30,77,31,31,31,93,31,179,31,136,31,149,31,73,31,61,31,249,31,172,31,172,30,35,31,27,31,211,31,211,30,2,31,74,31,3,31,65,31,48,31,91,31,207,31,46,31,60,31,60,30,65,31,45,31,194,31,29,31,23,31,23,30,171,31,151,31,140,31,192,31,192,30,4,31,4,30,3,31,3,30,3,29,130,31,130,30,105,31,174,31,174,30,174,29,128,31,53,31,53,30,53,29,243,31,6,31,178,31,153,31,163,31,220,31,14,31,14,30,173,31,117,31,145,31,208,31,208,30,180,31,226,31,174,31,174,30,254,31,254,30,254,29,164,31,49,31,188,31,105,31,76,31,236,31,236,30,244,31,244,30,244,29,8,31,171,31,27,31,188,31,146,31,67,31,94,31,94,30,240,31,240,30,191,31,196,31,253,31,116,31,249,31,171,31,171,30,178,31,122,31,122,30,148,31,148,30,148,29,158,31,158,30,190,31,190,30,20,31,147,31,165,31,225,31,191,31,214,31,188,31,234,31,80,31,173,31,47,31,36,31,212,31,34,31,1,31,176,31,176,30,125,31,11,31,244,31,244,30,73,31,201,31,119,31,48,31,161,31,237,31,21,31,21,30,186,31,121,31,121,30,26,31,215,31,31,31,128,31,167,31,231,31,231,30,8,31,8,31,114,31,114,30,127,31,178,31,74,31,200,31,95,31,241,31,241,30,221,31,86,31,106,31,17,31,192,31,229,31,233,31,208,31,117,31,85,31,143,31,143,30,159,31,159,30,119,31,119,30,50,31,18,31,156,31,225,31,65,31,65,30,108,31,53,31,100,31,114,31,70,31,141,31,147,31,128,31,128,30,131,31,131,30,195,31,208,31,210,31,226,31,116,31,195,31,195,30,207,31,207,30,15,31,106,31,81,31,81,30,161,31,90,31,90,30,56,31,73,31,173,31,160,31,36,31,138,31,188,31,22,31,22,30,181,31,201,31,125,31,132,31,132,30,128,31,136,31,198,31,99,31,151,31,151,30,207,31,207,30,207,29,207,28,220,31,183,31,183,30,92,31,106,31,101,31,241,31,161,31,115,31,204,31,204,30,204,29,84,31,130,31,116,31,218,31,59,31,4,31,214,31,181,31,105,31,102,31,202,31,18,31,164,31,129,31,129,30,125,31,107,31,107,30,107,29,226,31,226,30,114,31,191,31,43,31,192,31,30,31,218,31,62,31,70,31,76,31,76,30,73,31,99,31,38,31,179,31,179,30,161,31,182,31,97,31,148,31,238,31,108,31,55,31,216,31,216,30,216,29,193,31,238,31,227,31,234,31,37,31,1,31,1,30,149,31,138,31,250,31,208,31,7,31,105,31,6,31,185,31,71,31,208,31,39,31,39,30,25,31,25,30,25,29,38,31,101,31,8,31,137,31,231,31,231,30,136,31,136,31,42,31,42,30,119,31,17,31,218,31,22,31,24,31,65,31,30,31,30,30,30,29,174,31,52,31,218,31,170,31,205,31,205,30,205,29,109,31,220,31,220,30,168,31,82,31,98,31,20,31,20,30,20,29,88,31,154,31,125,31,181,31,181,30,87,31,11,31,11,30,133,31,65,31,55,31,55,30,27,31,114,31,128,31,200,31,155,31,79,31,79,30,251,31,251,30,90,31,177,31,82,31,218,31,43,31,27,31,142,31,195,31,60,31,45,31,174,31,87,31,249,31,169,31,101,31,32,31,251,31,251,30,216,31,216,30,28,31,28,30,22,31,215,31,121,31,156,31,109,31,177,31,90,31,122,31,40,31,90,31,90,30,90,29,184,31,104,31,20,31,219,31,219,30,19,31,31,31,19,31,108,31,108,30,218,31,149,31,230,31,230,30,200,31,154,31,95,31,170,31,58,31,5,31,226,31,128,31,54,31,113,31,59,31,49,31,217,31,135,31,245,31,245,30,245,29,245,28,245,27,254,31,95,31,64,31,20,31,145,31,213,31,46,31,64,31,93,31,194,31,29,31,208,31,208,30,176,31,176,30,176,29,236,31,172,31,20,31,151,31,254,31,47,31,133,31,133,30,75,31,28,31,127,31,29,31,16,31,131,31,5,31,124,31,196,31,22,31,22,30,217,31,146,31,192,31,192,30,40,31,16,31,43,31,45,31,240,31,240,30,51,31,240,31,17,31,17,30,20,31,41,31,224,31,88,31,230,31,230,30,83,31,10,31,175,31,175,30,186,31,230,31,222,31,183,31,255,31,255,31,210,31,89,31,89,30,240,31,251,31,251,30,251,29,172,31,11,31,149,31,83,31,83,30,131,31,131,30,242,31,242,30,242,29,201,31,201,30,201,29,190,31,12,31,192,31,114,31,129,31,212,31,212,31,5,31,5,30,96,31,51,31,51,30,33,31,33,30,33,29,32,31,213,31,166,31,125,31,125,30,134,31,61,31,75,31,81,31,81,30,157,31,212,31,212,30,74,31,74,30,164,31,31,31,31,30,31,29,31,28,164,31,141,31,78,31,78,30,78,29,62,31,62,30,221,31,221,30,63,31,63,30,63,29,223,31,205,31,175,31,175,30,175,29,106,31,86,31,178,31,12,31,12,30,12,29,164,31,164,30,117,31,221,31,221,30,90,31,70,31,240,31,65,31,54,31,73,31,56,31,56,30,230,31,176,31,252,31,252,31,217,31,19,31,118,31,103,31,237,31,174,31,162,31,162,30,61,31,123,31,13,31,205,31,205,30,112,31,112,30,135,31,11,31,124,31,66,31,243,31,70,31,68,31,101,31,41,31,107,31,129,31,10,31,129,31,33,31,18,31,131,31,131,30,219,31,48,31,206,31,152,31,11,31,77,31,228,31,171,31,99,31,99,30,241,31,241,30,118,31,133,31,7,31,7,30,7,29,82,31,168,31,196,31,112,31,15,31,139,31,139,30,11,31,112,31,115,31,186,31,24,31,120,31,120,30,53,31,9,31,91,31,86,31,133,31,133,30,133,29,82,31,93,31,90,31,45,31,136,31,179,31,17,31,145,31,205,31,160,31,160,30,118,31,110,31,217,31,26,31,171,31,104,31,253,31,207,31,57,31,220,31,171,31,6,31,6,30,96,31,98,31,98,30,8,31,156,31,247,31,17,31,244,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
