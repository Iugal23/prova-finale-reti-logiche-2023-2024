-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 918;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,91,0,197,0,12,0,255,0,237,0,0,0,210,0,0,0,37,0,0,0,107,0,79,0,213,0,61,0,167,0,0,0,226,0,0,0,10,0,51,0,141,0,21,0,74,0,5,0,51,0,115,0,0,0,12,0,183,0,224,0,159,0,86,0,91,0,26,0,23,0,164,0,38,0,29,0,0,0,119,0,0,0,75,0,158,0,177,0,0,0,86,0,44,0,52,0,85,0,0,0,56,0,0,0,194,0,0,0,88,0,41,0,231,0,200,0,62,0,50,0,114,0,154,0,0,0,185,0,174,0,143,0,133,0,97,0,18,0,230,0,141,0,13,0,120,0,117,0,249,0,69,0,247,0,93,0,0,0,66,0,0,0,15,0,184,0,211,0,22,0,144,0,102,0,47,0,111,0,211,0,26,0,220,0,0,0,217,0,169,0,141,0,97,0,245,0,0,0,249,0,75,0,104,0,227,0,203,0,11,0,63,0,252,0,141,0,58,0,0,0,199,0,221,0,79,0,0,0,55,0,17,0,127,0,0,0,18,0,111,0,149,0,121,0,0,0,40,0,0,0,68,0,0,0,0,0,0,0,204,0,58,0,131,0,30,0,206,0,45,0,203,0,127,0,61,0,135,0,237,0,170,0,219,0,86,0,9,0,0,0,13,0,0,0,59,0,23,0,227,0,38,0,89,0,64,0,0,0,178,0,199,0,222,0,0,0,93,0,254,0,209,0,136,0,13,0,177,0,191,0,238,0,33,0,156,0,72,0,0,0,36,0,0,0,0,0,185,0,255,0,54,0,220,0,0,0,240,0,38,0,16,0,151,0,47,0,106,0,92,0,34,0,102,0,234,0,0,0,177,0,65,0,227,0,245,0,132,0,155,0,38,0,248,0,43,0,239,0,146,0,158,0,233,0,123,0,102,0,41,0,0,0,190,0,81,0,187,0,154,0,51,0,22,0,241,0,68,0,86,0,238,0,45,0,70,0,0,0,38,0,209,0,197,0,0,0,199,0,36,0,67,0,17,0,229,0,43,0,135,0,0,0,205,0,0,0,0,0,208,0,0,0,0,0,226,0,28,0,168,0,121,0,27,0,69,0,28,0,0,0,206,0,28,0,101,0,227,0,0,0,178,0,22,0,134,0,185,0,0,0,0,0,213,0,39,0,54,0,32,0,158,0,129,0,1,0,37,0,166,0,143,0,34,0,67,0,38,0,160,0,153,0,0,0,141,0,85,0,85,0,242,0,4,0,203,0,247,0,81,0,84,0,254,0,120,0,90,0,105,0,240,0,162,0,97,0,0,0,145,0,58,0,202,0,29,0,147,0,180,0,0,0,0,0,111,0,0,0,0,0,0,0,231,0,192,0,157,0,208,0,164,0,0,0,60,0,82,0,210,0,238,0,211,0,149,0,149,0,245,0,126,0,248,0,0,0,0,0,248,0,63,0,119,0,225,0,191,0,7,0,32,0,170,0,42,0,168,0,151,0,245,0,0,0,5,0,192,0,121,0,162,0,229,0,152,0,55,0,182,0,117,0,55,0,69,0,0,0,77,0,213,0,11,0,111,0,228,0,50,0,245,0,115,0,30,0,2,0,108,0,136,0,122,0,65,0,155,0,205,0,63,0,84,0,230,0,120,0,99,0,0,0,148,0,0,0,81,0,38,0,251,0,127,0,116,0,113,0,170,0,19,0,49,0,109,0,0,0,9,0,136,0,247,0,240,0,189,0,166,0,134,0,0,0,234,0,201,0,170,0,72,0,239,0,16,0,111,0,122,0,85,0,228,0,0,0,36,0,182,0,191,0,66,0,0,0,11,0,120,0,4,0,0,0,38,0,175,0,202,0,184,0,233,0,127,0,239,0,167,0,166,0,0,0,12,0,242,0,20,0,0,0,116,0,131,0,112,0,255,0,0,0,250,0,104,0,26,0,42,0,108,0,158,0,63,0,225,0,0,0,0,0,60,0,207,0,148,0,5,0,248,0,247,0,194,0,41,0,159,0,184,0,105,0,115,0,0,0,0,0,0,0,203,0,209,0,137,0,37,0,56,0,89,0,0,0,195,0,156,0,151,0,0,0,149,0,169,0,218,0,194,0,113,0,248,0,0,0,103,0,249,0,224,0,187,0,98,0,178,0,6,0,151,0,170,0,0,0,239,0,201,0,203,0,251,0,96,0,0,0,64,0,116,0,213,0,68,0,176,0,147,0,186,0,154,0,103,0,252,0,20,0,185,0,141,0,198,0,0,0,180,0,0,0,217,0,64,0,0,0,222,0,121,0,5,0,87,0,123,0,16,0,105,0,116,0,0,0,126,0,238,0,0,0,170,0,45,0,0,0,38,0,107,0,106,0,142,0,0,0,0,0,231,0,64,0,251,0,162,0,87,0,193,0,43,0,0,0,0,0,24,0,32,0,142,0,0,0,141,0,241,0,191,0,53,0,0,0,160,0,232,0,121,0,112,0,0,0,41,0,69,0,250,0,101,0,59,0,240,0,0,0,13,0,94,0,231,0,0,0,28,0,0,0,75,0,0,0,33,0,0,0,50,0,197,0,255,0,177,0,246,0,7,0,99,0,18,0,58,0,36,0,0,0,251,0,197,0,164,0,224,0,194,0,11,0,0,0,36,0,0,0,0,0,33,0,143,0,32,0,222,0,88,0,0,0,92,0,233,0,117,0,37,0,0,0,64,0,87,0,183,0,11,0,0,0,0,0,0,0,0,0,0,0,18,0,77,0,99,0,221,0,14,0,123,0,231,0,21,0,90,0,207,0,0,0,195,0,0,0,166,0,212,0,0,0,0,0,11,0,138,0,77,0,43,0,80,0,61,0,203,0,177,0,0,0,251,0,217,0,30,0,0,0,42,0,100,0,230,0,0,0,230,0,214,0,213,0,87,0,154,0,92,0,97,0,190,0,0,0,55,0,254,0,0,0,173,0,18,0,58,0,178,0,112,0,92,0,50,0,206,0,219,0,111,0,25,0,231,0,59,0,172,0,189,0,0,0,26,0,244,0,106,0,106,0,19,0,200,0,0,0,193,0,99,0,168,0,138,0,42,0,36,0,25,0,0,0,0,0,0,0,166,0,115,0,0,0,161,0,33,0,134,0,31,0,162,0,0,0,40,0,127,0,107,0,62,0,110,0,0,0,42,0,60,0,31,0,244,0,54,0,41,0,0,0,0,0,197,0,238,0,119,0,93,0,0,0,199,0,144,0,0,0,58,0,85,0,237,0,160,0,46,0,177,0,210,0,251,0,140,0,0,0,182,0,148,0,92,0,242,0,246,0,0,0,150,0,0,0,57,0,120,0,239,0,204,0,12,0,143,0,41,0,10,0,119,0,165,0,249,0,202,0,254,0,174,0,230,0,176,0,242,0,245,0,48,0,8,0,106,0,28,0,41,0,28,0,238,0,175,0,67,0,3,0,54,0,119,0,99,0,83,0,180,0,109,0,0,0,0,0,0,0,41,0,78,0,0,0,195,0,84,0,173,0,235,0,168,0,117,0,0,0,0,0,54,0,249,0,95,0,203,0,159,0,32,0,0,0,0,0,0,0,133,0,196,0,42,0,248,0,225,0,187,0,42,0,206,0,28,0,0,0,181,0,101,0,226,0,161,0,206,0,22,0,3,0,78,0,223,0,90,0,129,0,204,0,54,0,168,0,192,0,24,0,0,0,14,0,10,0,214,0,220,0,177,0,116,0,61,0,71,0,147,0,0,0,182,0,3,0,76,0,239,0,254,0,95,0,43,0,191,0,211,0,53,0,0,0,59,0,58,0,192,0,0,0,0,0,161,0,6,0,0,0,0,0,159,0,206,0,0,0,229,0,194,0,0,0,0,0,69,0,157,0,213,0,0,0,221,0,85,0,0,0,97,0,45,0,179,0,190,0,156,0,181,0,197,0,0,0,0,0,157,0,152,0,168,0,130,0,115,0,0,0,213,0,68,0,241,0,0,0,213,0,0,0,250,0,0,0,0,0,61,0,59,0,137,0,155,0,128,0,253,0,6,0,46,0,138,0,125,0,72,0,41,0,104,0,83,0,115,0,150,0,240,0,212,0,195,0,98,0,213,0,233,0,86,0,40,0,150,0,0,0,0,0,0,0,161,0,16,0);
signal scenario_full  : scenario_type := (0,0,91,31,197,31,12,31,255,31,237,31,237,30,210,31,210,30,37,31,37,30,107,31,79,31,213,31,61,31,167,31,167,30,226,31,226,30,10,31,51,31,141,31,21,31,74,31,5,31,51,31,115,31,115,30,12,31,183,31,224,31,159,31,86,31,91,31,26,31,23,31,164,31,38,31,29,31,29,30,119,31,119,30,75,31,158,31,177,31,177,30,86,31,44,31,52,31,85,31,85,30,56,31,56,30,194,31,194,30,88,31,41,31,231,31,200,31,62,31,50,31,114,31,154,31,154,30,185,31,174,31,143,31,133,31,97,31,18,31,230,31,141,31,13,31,120,31,117,31,249,31,69,31,247,31,93,31,93,30,66,31,66,30,15,31,184,31,211,31,22,31,144,31,102,31,47,31,111,31,211,31,26,31,220,31,220,30,217,31,169,31,141,31,97,31,245,31,245,30,249,31,75,31,104,31,227,31,203,31,11,31,63,31,252,31,141,31,58,31,58,30,199,31,221,31,79,31,79,30,55,31,17,31,127,31,127,30,18,31,111,31,149,31,121,31,121,30,40,31,40,30,68,31,68,30,68,29,68,28,204,31,58,31,131,31,30,31,206,31,45,31,203,31,127,31,61,31,135,31,237,31,170,31,219,31,86,31,9,31,9,30,13,31,13,30,59,31,23,31,227,31,38,31,89,31,64,31,64,30,178,31,199,31,222,31,222,30,93,31,254,31,209,31,136,31,13,31,177,31,191,31,238,31,33,31,156,31,72,31,72,30,36,31,36,30,36,29,185,31,255,31,54,31,220,31,220,30,240,31,38,31,16,31,151,31,47,31,106,31,92,31,34,31,102,31,234,31,234,30,177,31,65,31,227,31,245,31,132,31,155,31,38,31,248,31,43,31,239,31,146,31,158,31,233,31,123,31,102,31,41,31,41,30,190,31,81,31,187,31,154,31,51,31,22,31,241,31,68,31,86,31,238,31,45,31,70,31,70,30,38,31,209,31,197,31,197,30,199,31,36,31,67,31,17,31,229,31,43,31,135,31,135,30,205,31,205,30,205,29,208,31,208,30,208,29,226,31,28,31,168,31,121,31,27,31,69,31,28,31,28,30,206,31,28,31,101,31,227,31,227,30,178,31,22,31,134,31,185,31,185,30,185,29,213,31,39,31,54,31,32,31,158,31,129,31,1,31,37,31,166,31,143,31,34,31,67,31,38,31,160,31,153,31,153,30,141,31,85,31,85,31,242,31,4,31,203,31,247,31,81,31,84,31,254,31,120,31,90,31,105,31,240,31,162,31,97,31,97,30,145,31,58,31,202,31,29,31,147,31,180,31,180,30,180,29,111,31,111,30,111,29,111,28,231,31,192,31,157,31,208,31,164,31,164,30,60,31,82,31,210,31,238,31,211,31,149,31,149,31,245,31,126,31,248,31,248,30,248,29,248,31,63,31,119,31,225,31,191,31,7,31,32,31,170,31,42,31,168,31,151,31,245,31,245,30,5,31,192,31,121,31,162,31,229,31,152,31,55,31,182,31,117,31,55,31,69,31,69,30,77,31,213,31,11,31,111,31,228,31,50,31,245,31,115,31,30,31,2,31,108,31,136,31,122,31,65,31,155,31,205,31,63,31,84,31,230,31,120,31,99,31,99,30,148,31,148,30,81,31,38,31,251,31,127,31,116,31,113,31,170,31,19,31,49,31,109,31,109,30,9,31,136,31,247,31,240,31,189,31,166,31,134,31,134,30,234,31,201,31,170,31,72,31,239,31,16,31,111,31,122,31,85,31,228,31,228,30,36,31,182,31,191,31,66,31,66,30,11,31,120,31,4,31,4,30,38,31,175,31,202,31,184,31,233,31,127,31,239,31,167,31,166,31,166,30,12,31,242,31,20,31,20,30,116,31,131,31,112,31,255,31,255,30,250,31,104,31,26,31,42,31,108,31,158,31,63,31,225,31,225,30,225,29,60,31,207,31,148,31,5,31,248,31,247,31,194,31,41,31,159,31,184,31,105,31,115,31,115,30,115,29,115,28,203,31,209,31,137,31,37,31,56,31,89,31,89,30,195,31,156,31,151,31,151,30,149,31,169,31,218,31,194,31,113,31,248,31,248,30,103,31,249,31,224,31,187,31,98,31,178,31,6,31,151,31,170,31,170,30,239,31,201,31,203,31,251,31,96,31,96,30,64,31,116,31,213,31,68,31,176,31,147,31,186,31,154,31,103,31,252,31,20,31,185,31,141,31,198,31,198,30,180,31,180,30,217,31,64,31,64,30,222,31,121,31,5,31,87,31,123,31,16,31,105,31,116,31,116,30,126,31,238,31,238,30,170,31,45,31,45,30,38,31,107,31,106,31,142,31,142,30,142,29,231,31,64,31,251,31,162,31,87,31,193,31,43,31,43,30,43,29,24,31,32,31,142,31,142,30,141,31,241,31,191,31,53,31,53,30,160,31,232,31,121,31,112,31,112,30,41,31,69,31,250,31,101,31,59,31,240,31,240,30,13,31,94,31,231,31,231,30,28,31,28,30,75,31,75,30,33,31,33,30,50,31,197,31,255,31,177,31,246,31,7,31,99,31,18,31,58,31,36,31,36,30,251,31,197,31,164,31,224,31,194,31,11,31,11,30,36,31,36,30,36,29,33,31,143,31,32,31,222,31,88,31,88,30,92,31,233,31,117,31,37,31,37,30,64,31,87,31,183,31,11,31,11,30,11,29,11,28,11,27,11,26,18,31,77,31,99,31,221,31,14,31,123,31,231,31,21,31,90,31,207,31,207,30,195,31,195,30,166,31,212,31,212,30,212,29,11,31,138,31,77,31,43,31,80,31,61,31,203,31,177,31,177,30,251,31,217,31,30,31,30,30,42,31,100,31,230,31,230,30,230,31,214,31,213,31,87,31,154,31,92,31,97,31,190,31,190,30,55,31,254,31,254,30,173,31,18,31,58,31,178,31,112,31,92,31,50,31,206,31,219,31,111,31,25,31,231,31,59,31,172,31,189,31,189,30,26,31,244,31,106,31,106,31,19,31,200,31,200,30,193,31,99,31,168,31,138,31,42,31,36,31,25,31,25,30,25,29,25,28,166,31,115,31,115,30,161,31,33,31,134,31,31,31,162,31,162,30,40,31,127,31,107,31,62,31,110,31,110,30,42,31,60,31,31,31,244,31,54,31,41,31,41,30,41,29,197,31,238,31,119,31,93,31,93,30,199,31,144,31,144,30,58,31,85,31,237,31,160,31,46,31,177,31,210,31,251,31,140,31,140,30,182,31,148,31,92,31,242,31,246,31,246,30,150,31,150,30,57,31,120,31,239,31,204,31,12,31,143,31,41,31,10,31,119,31,165,31,249,31,202,31,254,31,174,31,230,31,176,31,242,31,245,31,48,31,8,31,106,31,28,31,41,31,28,31,238,31,175,31,67,31,3,31,54,31,119,31,99,31,83,31,180,31,109,31,109,30,109,29,109,28,41,31,78,31,78,30,195,31,84,31,173,31,235,31,168,31,117,31,117,30,117,29,54,31,249,31,95,31,203,31,159,31,32,31,32,30,32,29,32,28,133,31,196,31,42,31,248,31,225,31,187,31,42,31,206,31,28,31,28,30,181,31,101,31,226,31,161,31,206,31,22,31,3,31,78,31,223,31,90,31,129,31,204,31,54,31,168,31,192,31,24,31,24,30,14,31,10,31,214,31,220,31,177,31,116,31,61,31,71,31,147,31,147,30,182,31,3,31,76,31,239,31,254,31,95,31,43,31,191,31,211,31,53,31,53,30,59,31,58,31,192,31,192,30,192,29,161,31,6,31,6,30,6,29,159,31,206,31,206,30,229,31,194,31,194,30,194,29,69,31,157,31,213,31,213,30,221,31,85,31,85,30,97,31,45,31,179,31,190,31,156,31,181,31,197,31,197,30,197,29,157,31,152,31,168,31,130,31,115,31,115,30,213,31,68,31,241,31,241,30,213,31,213,30,250,31,250,30,250,29,61,31,59,31,137,31,155,31,128,31,253,31,6,31,46,31,138,31,125,31,72,31,41,31,104,31,83,31,115,31,150,31,240,31,212,31,195,31,98,31,213,31,233,31,86,31,40,31,150,31,150,30,150,29,150,28,161,31,16,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
