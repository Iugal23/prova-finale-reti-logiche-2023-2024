-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 543;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,180,0,56,0,231,0,236,0,0,0,112,0,70,0,0,0,134,0,242,0,198,0,107,0,238,0,57,0,0,0,166,0,49,0,207,0,0,0,119,0,255,0,24,0,250,0,217,0,95,0,96,0,54,0,29,0,0,0,96,0,163,0,239,0,200,0,0,0,132,0,179,0,0,0,150,0,0,0,41,0,0,0,134,0,149,0,14,0,69,0,0,0,190,0,184,0,213,0,229,0,0,0,0,0,0,0,82,0,0,0,232,0,101,0,43,0,16,0,136,0,189,0,87,0,27,0,115,0,106,0,62,0,227,0,99,0,0,0,0,0,148,0,113,0,20,0,112,0,171,0,0,0,141,0,0,0,0,0,216,0,0,0,237,0,197,0,185,0,227,0,247,0,249,0,0,0,252,0,102,0,110,0,5,0,51,0,194,0,172,0,86,0,106,0,0,0,69,0,0,0,96,0,203,0,121,0,14,0,126,0,66,0,190,0,175,0,253,0,155,0,170,0,174,0,0,0,207,0,182,0,136,0,0,0,76,0,61,0,198,0,84,0,122,0,154,0,0,0,52,0,195,0,34,0,0,0,32,0,223,0,88,0,0,0,94,0,23,0,168,0,61,0,28,0,105,0,0,0,0,0,233,0,205,0,143,0,193,0,234,0,231,0,179,0,1,0,161,0,132,0,0,0,198,0,130,0,102,0,0,0,11,0,253,0,7,0,192,0,158,0,92,0,0,0,44,0,78,0,129,0,116,0,114,0,172,0,0,0,36,0,243,0,39,0,205,0,108,0,222,0,70,0,99,0,166,0,254,0,0,0,13,0,177,0,18,0,238,0,0,0,210,0,152,0,242,0,151,0,179,0,36,0,76,0,147,0,150,0,96,0,0,0,216,0,25,0,246,0,242,0,244,0,164,0,0,0,0,0,0,0,66,0,0,0,68,0,116,0,177,0,0,0,156,0,60,0,5,0,11,0,126,0,162,0,0,0,136,0,208,0,165,0,178,0,138,0,247,0,132,0,22,0,117,0,70,0,210,0,198,0,145,0,0,0,34,0,34,0,248,0,228,0,247,0,191,0,0,0,82,0,70,0,0,0,103,0,8,0,231,0,231,0,0,0,53,0,7,0,193,0,153,0,108,0,196,0,93,0,26,0,3,0,194,0,8,0,204,0,0,0,156,0,0,0,219,0,0,0,49,0,186,0,64,0,29,0,68,0,65,0,92,0,101,0,251,0,47,0,202,0,220,0,222,0,130,0,81,0,235,0,95,0,13,0,176,0,230,0,90,0,70,0,0,0,0,0,0,0,220,0,211,0,209,0,46,0,238,0,61,0,84,0,0,0,42,0,208,0,150,0,154,0,148,0,194,0,190,0,0,0,236,0,0,0,98,0,70,0,240,0,51,0,179,0,237,0,189,0,161,0,245,0,227,0,123,0,77,0,0,0,200,0,229,0,233,0,219,0,0,0,100,0,0,0,64,0,116,0,0,0,69,0,50,0,153,0,0,0,171,0,3,0,146,0,79,0,165,0,73,0,31,0,146,0,105,0,104,0,147,0,180,0,246,0,0,0,22,0,173,0,0,0,242,0,31,0,69,0,85,0,62,0,0,0,0,0,49,0,25,0,0,0,184,0,0,0,170,0,223,0,213,0,14,0,171,0,179,0,148,0,17,0,254,0,0,0,21,0,222,0,219,0,0,0,217,0,0,0,0,0,0,0,233,0,233,0,23,0,117,0,0,0,253,0,171,0,55,0,201,0,0,0,119,0,48,0,223,0,4,0,99,0,207,0,72,0,230,0,0,0,206,0,0,0,243,0,181,0,125,0,141,0,81,0,243,0,137,0,221,0,95,0,40,0,0,0,166,0,163,0,0,0,169,0,80,0,0,0,85,0,100,0,121,0,79,0,9,0,1,0,39,0,70,0,0,0,0,0,189,0,216,0,41,0,187,0,233,0,46,0,224,0,124,0,240,0,167,0,0,0,231,0,116,0,227,0,207,0,140,0,231,0,204,0,0,0,0,0,118,0,205,0,176,0,168,0,14,0,61,0,252,0,50,0,240,0,37,0,84,0,5,0,169,0,68,0,0,0,189,0,240,0,0,0,161,0,172,0,72,0,248,0,134,0,162,0,208,0,0,0,47,0,164,0,0,0,6,0,222,0,152,0,149,0,155,0,114,0,78,0,30,0,123,0,207,0,168,0,187,0,0,0,106,0,137,0,79,0,0,0,225,0,243,0,0,0,34,0,37,0,8,0,123,0,99,0,94,0,149,0,131,0,99,0,220,0,24,0,10,0,0,0,231,0,184,0,190,0,51,0,129,0,34,0,116,0,207,0,173,0,120,0,234,0,0,0,111,0,187,0,216,0,235,0,144,0,193,0,62,0,0,0,66,0,100,0,43,0,152,0,5,0,26,0,0,0,0,0,0,0,0,0,133,0);
signal scenario_full  : scenario_type := (0,0,180,31,56,31,231,31,236,31,236,30,112,31,70,31,70,30,134,31,242,31,198,31,107,31,238,31,57,31,57,30,166,31,49,31,207,31,207,30,119,31,255,31,24,31,250,31,217,31,95,31,96,31,54,31,29,31,29,30,96,31,163,31,239,31,200,31,200,30,132,31,179,31,179,30,150,31,150,30,41,31,41,30,134,31,149,31,14,31,69,31,69,30,190,31,184,31,213,31,229,31,229,30,229,29,229,28,82,31,82,30,232,31,101,31,43,31,16,31,136,31,189,31,87,31,27,31,115,31,106,31,62,31,227,31,99,31,99,30,99,29,148,31,113,31,20,31,112,31,171,31,171,30,141,31,141,30,141,29,216,31,216,30,237,31,197,31,185,31,227,31,247,31,249,31,249,30,252,31,102,31,110,31,5,31,51,31,194,31,172,31,86,31,106,31,106,30,69,31,69,30,96,31,203,31,121,31,14,31,126,31,66,31,190,31,175,31,253,31,155,31,170,31,174,31,174,30,207,31,182,31,136,31,136,30,76,31,61,31,198,31,84,31,122,31,154,31,154,30,52,31,195,31,34,31,34,30,32,31,223,31,88,31,88,30,94,31,23,31,168,31,61,31,28,31,105,31,105,30,105,29,233,31,205,31,143,31,193,31,234,31,231,31,179,31,1,31,161,31,132,31,132,30,198,31,130,31,102,31,102,30,11,31,253,31,7,31,192,31,158,31,92,31,92,30,44,31,78,31,129,31,116,31,114,31,172,31,172,30,36,31,243,31,39,31,205,31,108,31,222,31,70,31,99,31,166,31,254,31,254,30,13,31,177,31,18,31,238,31,238,30,210,31,152,31,242,31,151,31,179,31,36,31,76,31,147,31,150,31,96,31,96,30,216,31,25,31,246,31,242,31,244,31,164,31,164,30,164,29,164,28,66,31,66,30,68,31,116,31,177,31,177,30,156,31,60,31,5,31,11,31,126,31,162,31,162,30,136,31,208,31,165,31,178,31,138,31,247,31,132,31,22,31,117,31,70,31,210,31,198,31,145,31,145,30,34,31,34,31,248,31,228,31,247,31,191,31,191,30,82,31,70,31,70,30,103,31,8,31,231,31,231,31,231,30,53,31,7,31,193,31,153,31,108,31,196,31,93,31,26,31,3,31,194,31,8,31,204,31,204,30,156,31,156,30,219,31,219,30,49,31,186,31,64,31,29,31,68,31,65,31,92,31,101,31,251,31,47,31,202,31,220,31,222,31,130,31,81,31,235,31,95,31,13,31,176,31,230,31,90,31,70,31,70,30,70,29,70,28,220,31,211,31,209,31,46,31,238,31,61,31,84,31,84,30,42,31,208,31,150,31,154,31,148,31,194,31,190,31,190,30,236,31,236,30,98,31,70,31,240,31,51,31,179,31,237,31,189,31,161,31,245,31,227,31,123,31,77,31,77,30,200,31,229,31,233,31,219,31,219,30,100,31,100,30,64,31,116,31,116,30,69,31,50,31,153,31,153,30,171,31,3,31,146,31,79,31,165,31,73,31,31,31,146,31,105,31,104,31,147,31,180,31,246,31,246,30,22,31,173,31,173,30,242,31,31,31,69,31,85,31,62,31,62,30,62,29,49,31,25,31,25,30,184,31,184,30,170,31,223,31,213,31,14,31,171,31,179,31,148,31,17,31,254,31,254,30,21,31,222,31,219,31,219,30,217,31,217,30,217,29,217,28,233,31,233,31,23,31,117,31,117,30,253,31,171,31,55,31,201,31,201,30,119,31,48,31,223,31,4,31,99,31,207,31,72,31,230,31,230,30,206,31,206,30,243,31,181,31,125,31,141,31,81,31,243,31,137,31,221,31,95,31,40,31,40,30,166,31,163,31,163,30,169,31,80,31,80,30,85,31,100,31,121,31,79,31,9,31,1,31,39,31,70,31,70,30,70,29,189,31,216,31,41,31,187,31,233,31,46,31,224,31,124,31,240,31,167,31,167,30,231,31,116,31,227,31,207,31,140,31,231,31,204,31,204,30,204,29,118,31,205,31,176,31,168,31,14,31,61,31,252,31,50,31,240,31,37,31,84,31,5,31,169,31,68,31,68,30,189,31,240,31,240,30,161,31,172,31,72,31,248,31,134,31,162,31,208,31,208,30,47,31,164,31,164,30,6,31,222,31,152,31,149,31,155,31,114,31,78,31,30,31,123,31,207,31,168,31,187,31,187,30,106,31,137,31,79,31,79,30,225,31,243,31,243,30,34,31,37,31,8,31,123,31,99,31,94,31,149,31,131,31,99,31,220,31,24,31,10,31,10,30,231,31,184,31,190,31,51,31,129,31,34,31,116,31,207,31,173,31,120,31,234,31,234,30,111,31,187,31,216,31,235,31,144,31,193,31,62,31,62,30,66,31,100,31,43,31,152,31,5,31,26,31,26,30,26,29,26,28,26,27,133,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
