-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 258;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (93,0,0,0,16,0,148,0,41,0,84,0,107,0,220,0,105,0,0,0,35,0,98,0,0,0,133,0,63,0,128,0,251,0,152,0,36,0,30,0,0,0,105,0,128,0,16,0,57,0,150,0,0,0,80,0,11,0,0,0,187,0,247,0,0,0,40,0,145,0,0,0,160,0,245,0,2,0,140,0,0,0,21,0,12,0,241,0,172,0,127,0,1,0,21,0,68,0,128,0,64,0,215,0,0,0,251,0,152,0,117,0,144,0,64,0,96,0,31,0,114,0,80,0,0,0,0,0,0,0,23,0,161,0,203,0,84,0,101,0,107,0,7,0,0,0,49,0,203,0,81,0,135,0,124,0,0,0,107,0,99,0,192,0,79,0,0,0,55,0,0,0,175,0,229,0,142,0,79,0,47,0,27,0,10,0,194,0,91,0,0,0,99,0,182,0,140,0,0,0,141,0,129,0,0,0,51,0,0,0,188,0,148,0,204,0,0,0,94,0,0,0,200,0,13,0,161,0,244,0,0,0,78,0,0,0,220,0,190,0,193,0,12,0,111,0,0,0,0,0,110,0,0,0,13,0,105,0,0,0,216,0,35,0,71,0,0,0,183,0,15,0,155,0,0,0,207,0,172,0,0,0,124,0,138,0,89,0,2,0,0,0,202,0,75,0,236,0,105,0,239,0,206,0,106,0,147,0,202,0,0,0,52,0,175,0,249,0,0,0,0,0,34,0,167,0,136,0,69,0,112,0,233,0,201,0,90,0,237,0,135,0,0,0,55,0,84,0,204,0,0,0,0,0,77,0,219,0,0,0,220,0,38,0,0,0,198,0,145,0,175,0,90,0,19,0,0,0,225,0,140,0,159,0,25,0,227,0,239,0,151,0,151,0,121,0,67,0,109,0,231,0,6,0,181,0,111,0,143,0,136,0,250,0,144,0,39,0,165,0,242,0,234,0,153,0,92,0,19,0,0,0,250,0,14,0,104,0,146,0,210,0,100,0,56,0,112,0,0,0,110,0,35,0,43,0,218,0,242,0,236,0,4,0,79,0,0,0,0,0,5,0,96,0,30,0,224,0,77,0,13,0,82,0,221,0,79,0,11,0,73,0,201,0,193,0,101,0,228,0,102,0,95,0,0,0,102,0,0,0,233,0,19,0,69,0);
signal scenario_full  : scenario_type := (93,31,93,30,16,31,148,31,41,31,84,31,107,31,220,31,105,31,105,30,35,31,98,31,98,30,133,31,63,31,128,31,251,31,152,31,36,31,30,31,30,30,105,31,128,31,16,31,57,31,150,31,150,30,80,31,11,31,11,30,187,31,247,31,247,30,40,31,145,31,145,30,160,31,245,31,2,31,140,31,140,30,21,31,12,31,241,31,172,31,127,31,1,31,21,31,68,31,128,31,64,31,215,31,215,30,251,31,152,31,117,31,144,31,64,31,96,31,31,31,114,31,80,31,80,30,80,29,80,28,23,31,161,31,203,31,84,31,101,31,107,31,7,31,7,30,49,31,203,31,81,31,135,31,124,31,124,30,107,31,99,31,192,31,79,31,79,30,55,31,55,30,175,31,229,31,142,31,79,31,47,31,27,31,10,31,194,31,91,31,91,30,99,31,182,31,140,31,140,30,141,31,129,31,129,30,51,31,51,30,188,31,148,31,204,31,204,30,94,31,94,30,200,31,13,31,161,31,244,31,244,30,78,31,78,30,220,31,190,31,193,31,12,31,111,31,111,30,111,29,110,31,110,30,13,31,105,31,105,30,216,31,35,31,71,31,71,30,183,31,15,31,155,31,155,30,207,31,172,31,172,30,124,31,138,31,89,31,2,31,2,30,202,31,75,31,236,31,105,31,239,31,206,31,106,31,147,31,202,31,202,30,52,31,175,31,249,31,249,30,249,29,34,31,167,31,136,31,69,31,112,31,233,31,201,31,90,31,237,31,135,31,135,30,55,31,84,31,204,31,204,30,204,29,77,31,219,31,219,30,220,31,38,31,38,30,198,31,145,31,175,31,90,31,19,31,19,30,225,31,140,31,159,31,25,31,227,31,239,31,151,31,151,31,121,31,67,31,109,31,231,31,6,31,181,31,111,31,143,31,136,31,250,31,144,31,39,31,165,31,242,31,234,31,153,31,92,31,19,31,19,30,250,31,14,31,104,31,146,31,210,31,100,31,56,31,112,31,112,30,110,31,35,31,43,31,218,31,242,31,236,31,4,31,79,31,79,30,79,29,5,31,96,31,30,31,224,31,77,31,13,31,82,31,221,31,79,31,11,31,73,31,201,31,193,31,101,31,228,31,102,31,95,31,95,30,102,31,102,30,233,31,19,31,69,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
