-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 540;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (205,0,0,0,0,0,18,0,0,0,183,0,213,0,170,0,136,0,137,0,32,0,234,0,0,0,69,0,33,0,191,0,234,0,216,0,0,0,127,0,199,0,17,0,0,0,138,0,181,0,84,0,86,0,108,0,219,0,141,0,72,0,245,0,0,0,69,0,184,0,0,0,40,0,194,0,83,0,190,0,237,0,11,0,0,0,12,0,229,0,0,0,0,0,190,0,77,0,159,0,132,0,103,0,0,0,55,0,0,0,155,0,31,0,0,0,73,0,120,0,0,0,0,0,104,0,173,0,0,0,185,0,81,0,111,0,59,0,111,0,0,0,53,0,28,0,0,0,174,0,112,0,151,0,47,0,0,0,0,0,160,0,0,0,26,0,0,0,10,0,132,0,0,0,74,0,218,0,173,0,113,0,0,0,12,0,108,0,149,0,102,0,46,0,0,0,222,0,132,0,160,0,0,0,151,0,123,0,151,0,143,0,62,0,54,0,83,0,176,0,56,0,67,0,177,0,71,0,84,0,93,0,193,0,80,0,14,0,223,0,0,0,197,0,0,0,0,0,162,0,29,0,0,0,0,0,0,0,0,0,25,0,96,0,88,0,99,0,169,0,44,0,119,0,0,0,13,0,187,0,37,0,13,0,93,0,113,0,211,0,224,0,99,0,208,0,171,0,115,0,185,0,248,0,78,0,165,0,25,0,56,0,62,0,42,0,229,0,26,0,0,0,84,0,202,0,168,0,0,0,121,0,39,0,202,0,8,0,0,0,63,0,58,0,93,0,21,0,29,0,186,0,5,0,0,0,0,0,109,0,31,0,120,0,85,0,38,0,0,0,254,0,0,0,186,0,230,0,58,0,3,0,8,0,255,0,232,0,140,0,0,0,29,0,65,0,234,0,0,0,0,0,0,0,203,0,210,0,16,0,224,0,77,0,122,0,124,0,97,0,50,0,207,0,0,0,53,0,220,0,183,0,188,0,141,0,0,0,46,0,0,0,121,0,0,0,242,0,146,0,67,0,204,0,248,0,3,0,213,0,0,0,68,0,184,0,220,0,0,0,84,0,0,0,18,0,24,0,106,0,166,0,109,0,225,0,177,0,38,0,183,0,0,0,157,0,243,0,196,0,127,0,48,0,59,0,0,0,177,0,100,0,6,0,98,0,226,0,0,0,251,0,137,0,139,0,181,0,0,0,198,0,210,0,76,0,243,0,0,0,156,0,24,0,0,0,231,0,34,0,102,0,69,0,0,0,55,0,0,0,126,0,120,0,171,0,0,0,34,0,72,0,210,0,219,0,27,0,68,0,179,0,0,0,204,0,172,0,186,0,232,0,47,0,4,0,98,0,18,0,77,0,0,0,18,0,197,0,97,0,41,0,98,0,215,0,145,0,229,0,52,0,40,0,144,0,102,0,175,0,145,0,177,0,173,0,172,0,214,0,122,0,113,0,0,0,86,0,87,0,163,0,0,0,109,0,115,0,180,0,0,0,1,0,243,0,106,0,0,0,0,0,198,0,0,0,68,0,48,0,0,0,160,0,0,0,45,0,26,0,221,0,0,0,55,0,37,0,0,0,38,0,14,0,100,0,30,0,225,0,0,0,132,0,0,0,0,0,214,0,54,0,97,0,0,0,2,0,140,0,186,0,0,0,226,0,228,0,120,0,251,0,253,0,165,0,227,0,11,0,27,0,2,0,0,0,245,0,70,0,187,0,10,0,79,0,179,0,231,0,218,0,145,0,228,0,249,0,179,0,0,0,240,0,0,0,240,0,0,0,86,0,232,0,242,0,1,0,138,0,79,0,95,0,0,0,28,0,163,0,244,0,243,0,241,0,113,0,179,0,0,0,171,0,77,0,0,0,82,0,30,0,71,0,0,0,160,0,142,0,207,0,12,0,66,0,32,0,6,0,0,0,27,0,107,0,182,0,167,0,110,0,125,0,180,0,51,0,77,0,111,0,0,0,176,0,0,0,34,0,124,0,168,0,21,0,90,0,144,0,135,0,226,0,239,0,0,0,69,0,171,0,220,0,49,0,25,0,73,0,0,0,223,0,124,0,22,0,56,0,212,0,249,0,42,0,124,0,118,0,66,0,228,0,53,0,198,0,250,0,102,0,134,0,125,0,147,0,148,0,116,0,141,0,149,0,48,0,249,0,164,0,0,0,23,0,84,0,0,0,0,0,136,0,91,0,142,0,49,0,193,0,132,0,118,0,76,0,90,0,134,0,184,0,50,0,0,0,0,0,0,0,23,0,140,0,48,0,1,0,199,0,0,0,134,0,153,0,210,0,221,0,82,0,150,0,185,0,0,0,0,0,0,0,67,0,0,0,242,0,0,0,121,0,30,0,0,0,89,0,55,0,236,0,73,0,36,0,85,0,215,0,221,0,0,0,253,0,117,0,132,0,0,0,189,0,107,0,0,0);
signal scenario_full  : scenario_type := (205,31,205,30,205,29,18,31,18,30,183,31,213,31,170,31,136,31,137,31,32,31,234,31,234,30,69,31,33,31,191,31,234,31,216,31,216,30,127,31,199,31,17,31,17,30,138,31,181,31,84,31,86,31,108,31,219,31,141,31,72,31,245,31,245,30,69,31,184,31,184,30,40,31,194,31,83,31,190,31,237,31,11,31,11,30,12,31,229,31,229,30,229,29,190,31,77,31,159,31,132,31,103,31,103,30,55,31,55,30,155,31,31,31,31,30,73,31,120,31,120,30,120,29,104,31,173,31,173,30,185,31,81,31,111,31,59,31,111,31,111,30,53,31,28,31,28,30,174,31,112,31,151,31,47,31,47,30,47,29,160,31,160,30,26,31,26,30,10,31,132,31,132,30,74,31,218,31,173,31,113,31,113,30,12,31,108,31,149,31,102,31,46,31,46,30,222,31,132,31,160,31,160,30,151,31,123,31,151,31,143,31,62,31,54,31,83,31,176,31,56,31,67,31,177,31,71,31,84,31,93,31,193,31,80,31,14,31,223,31,223,30,197,31,197,30,197,29,162,31,29,31,29,30,29,29,29,28,29,27,25,31,96,31,88,31,99,31,169,31,44,31,119,31,119,30,13,31,187,31,37,31,13,31,93,31,113,31,211,31,224,31,99,31,208,31,171,31,115,31,185,31,248,31,78,31,165,31,25,31,56,31,62,31,42,31,229,31,26,31,26,30,84,31,202,31,168,31,168,30,121,31,39,31,202,31,8,31,8,30,63,31,58,31,93,31,21,31,29,31,186,31,5,31,5,30,5,29,109,31,31,31,120,31,85,31,38,31,38,30,254,31,254,30,186,31,230,31,58,31,3,31,8,31,255,31,232,31,140,31,140,30,29,31,65,31,234,31,234,30,234,29,234,28,203,31,210,31,16,31,224,31,77,31,122,31,124,31,97,31,50,31,207,31,207,30,53,31,220,31,183,31,188,31,141,31,141,30,46,31,46,30,121,31,121,30,242,31,146,31,67,31,204,31,248,31,3,31,213,31,213,30,68,31,184,31,220,31,220,30,84,31,84,30,18,31,24,31,106,31,166,31,109,31,225,31,177,31,38,31,183,31,183,30,157,31,243,31,196,31,127,31,48,31,59,31,59,30,177,31,100,31,6,31,98,31,226,31,226,30,251,31,137,31,139,31,181,31,181,30,198,31,210,31,76,31,243,31,243,30,156,31,24,31,24,30,231,31,34,31,102,31,69,31,69,30,55,31,55,30,126,31,120,31,171,31,171,30,34,31,72,31,210,31,219,31,27,31,68,31,179,31,179,30,204,31,172,31,186,31,232,31,47,31,4,31,98,31,18,31,77,31,77,30,18,31,197,31,97,31,41,31,98,31,215,31,145,31,229,31,52,31,40,31,144,31,102,31,175,31,145,31,177,31,173,31,172,31,214,31,122,31,113,31,113,30,86,31,87,31,163,31,163,30,109,31,115,31,180,31,180,30,1,31,243,31,106,31,106,30,106,29,198,31,198,30,68,31,48,31,48,30,160,31,160,30,45,31,26,31,221,31,221,30,55,31,37,31,37,30,38,31,14,31,100,31,30,31,225,31,225,30,132,31,132,30,132,29,214,31,54,31,97,31,97,30,2,31,140,31,186,31,186,30,226,31,228,31,120,31,251,31,253,31,165,31,227,31,11,31,27,31,2,31,2,30,245,31,70,31,187,31,10,31,79,31,179,31,231,31,218,31,145,31,228,31,249,31,179,31,179,30,240,31,240,30,240,31,240,30,86,31,232,31,242,31,1,31,138,31,79,31,95,31,95,30,28,31,163,31,244,31,243,31,241,31,113,31,179,31,179,30,171,31,77,31,77,30,82,31,30,31,71,31,71,30,160,31,142,31,207,31,12,31,66,31,32,31,6,31,6,30,27,31,107,31,182,31,167,31,110,31,125,31,180,31,51,31,77,31,111,31,111,30,176,31,176,30,34,31,124,31,168,31,21,31,90,31,144,31,135,31,226,31,239,31,239,30,69,31,171,31,220,31,49,31,25,31,73,31,73,30,223,31,124,31,22,31,56,31,212,31,249,31,42,31,124,31,118,31,66,31,228,31,53,31,198,31,250,31,102,31,134,31,125,31,147,31,148,31,116,31,141,31,149,31,48,31,249,31,164,31,164,30,23,31,84,31,84,30,84,29,136,31,91,31,142,31,49,31,193,31,132,31,118,31,76,31,90,31,134,31,184,31,50,31,50,30,50,29,50,28,23,31,140,31,48,31,1,31,199,31,199,30,134,31,153,31,210,31,221,31,82,31,150,31,185,31,185,30,185,29,185,28,67,31,67,30,242,31,242,30,121,31,30,31,30,30,89,31,55,31,236,31,73,31,36,31,85,31,215,31,221,31,221,30,253,31,117,31,132,31,132,30,189,31,107,31,107,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
