-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_467 is
end project_tb_467;

architecture project_tb_arch_467 of project_tb_467 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 346;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (240,0,0,0,29,0,120,0,248,0,151,0,38,0,160,0,122,0,117,0,112,0,4,0,0,0,0,0,7,0,6,0,126,0,224,0,33,0,207,0,217,0,0,0,174,0,0,0,215,0,143,0,0,0,46,0,173,0,128,0,208,0,72,0,43,0,0,0,0,0,56,0,0,0,0,0,114,0,58,0,56,0,188,0,161,0,177,0,0,0,121,0,45,0,15,0,88,0,71,0,168,0,0,0,180,0,7,0,7,0,98,0,0,0,75,0,0,0,158,0,47,0,0,0,0,0,0,0,80,0,106,0,160,0,188,0,35,0,0,0,66,0,121,0,0,0,176,0,101,0,241,0,10,0,0,0,88,0,0,0,219,0,131,0,0,0,71,0,0,0,213,0,221,0,0,0,130,0,149,0,0,0,180,0,14,0,111,0,229,0,53,0,102,0,76,0,53,0,38,0,0,0,40,0,57,0,6,0,0,0,188,0,184,0,72,0,221,0,0,0,166,0,0,0,0,0,0,0,0,0,63,0,73,0,0,0,95,0,78,0,103,0,14,0,64,0,84,0,246,0,0,0,252,0,69,0,197,0,255,0,0,0,238,0,53,0,0,0,0,0,88,0,141,0,213,0,0,0,161,0,191,0,94,0,151,0,27,0,116,0,0,0,97,0,169,0,155,0,168,0,53,0,240,0,37,0,0,0,186,0,91,0,11,0,133,0,41,0,0,0,184,0,95,0,228,0,233,0,75,0,0,0,146,0,226,0,0,0,113,0,52,0,64,0,98,0,135,0,178,0,202,0,191,0,0,0,107,0,57,0,0,0,177,0,171,0,179,0,0,0,141,0,129,0,0,0,72,0,169,0,208,0,244,0,40,0,42,0,135,0,110,0,0,0,7,0,252,0,193,0,10,0,251,0,117,0,0,0,182,0,161,0,89,0,192,0,213,0,159,0,30,0,31,0,206,0,0,0,178,0,91,0,127,0,124,0,9,0,169,0,79,0,55,0,203,0,201,0,70,0,93,0,62,0,239,0,142,0,244,0,234,0,0,0,0,0,127,0,73,0,82,0,69,0,109,0,36,0,147,0,76,0,226,0,0,0,0,0,229,0,166,0,72,0,127,0,197,0,0,0,177,0,88,0,33,0,11,0,55,0,199,0,133,0,216,0,58,0,0,0,141,0,231,0,45,0,245,0,0,0,92,0,0,0,194,0,106,0,14,0,232,0,158,0,111,0,228,0,104,0,70,0,71,0,125,0,30,0,0,0,134,0,20,0,208,0,47,0,72,0,55,0,0,0,249,0,150,0,0,0,0,0,243,0,0,0,236,0,0,0,90,0,0,0,57,0,0,0,229,0,0,0,0,0,0,0,93,0,225,0,200,0,46,0,0,0,49,0,185,0,99,0,83,0,151,0,31,0,0,0,136,0,135,0,66,0,183,0,0,0,243,0,15,0,0,0,254,0,0,0,202,0,66,0,238,0,54,0,43,0,0,0,18,0,152,0,180,0,250,0,151,0,0,0,0,0,0,0,255,0,178,0,157,0,2,0,50,0,173,0,254,0);
signal scenario_full  : scenario_type := (240,31,240,30,29,31,120,31,248,31,151,31,38,31,160,31,122,31,117,31,112,31,4,31,4,30,4,29,7,31,6,31,126,31,224,31,33,31,207,31,217,31,217,30,174,31,174,30,215,31,143,31,143,30,46,31,173,31,128,31,208,31,72,31,43,31,43,30,43,29,56,31,56,30,56,29,114,31,58,31,56,31,188,31,161,31,177,31,177,30,121,31,45,31,15,31,88,31,71,31,168,31,168,30,180,31,7,31,7,31,98,31,98,30,75,31,75,30,158,31,47,31,47,30,47,29,47,28,80,31,106,31,160,31,188,31,35,31,35,30,66,31,121,31,121,30,176,31,101,31,241,31,10,31,10,30,88,31,88,30,219,31,131,31,131,30,71,31,71,30,213,31,221,31,221,30,130,31,149,31,149,30,180,31,14,31,111,31,229,31,53,31,102,31,76,31,53,31,38,31,38,30,40,31,57,31,6,31,6,30,188,31,184,31,72,31,221,31,221,30,166,31,166,30,166,29,166,28,166,27,63,31,73,31,73,30,95,31,78,31,103,31,14,31,64,31,84,31,246,31,246,30,252,31,69,31,197,31,255,31,255,30,238,31,53,31,53,30,53,29,88,31,141,31,213,31,213,30,161,31,191,31,94,31,151,31,27,31,116,31,116,30,97,31,169,31,155,31,168,31,53,31,240,31,37,31,37,30,186,31,91,31,11,31,133,31,41,31,41,30,184,31,95,31,228,31,233,31,75,31,75,30,146,31,226,31,226,30,113,31,52,31,64,31,98,31,135,31,178,31,202,31,191,31,191,30,107,31,57,31,57,30,177,31,171,31,179,31,179,30,141,31,129,31,129,30,72,31,169,31,208,31,244,31,40,31,42,31,135,31,110,31,110,30,7,31,252,31,193,31,10,31,251,31,117,31,117,30,182,31,161,31,89,31,192,31,213,31,159,31,30,31,31,31,206,31,206,30,178,31,91,31,127,31,124,31,9,31,169,31,79,31,55,31,203,31,201,31,70,31,93,31,62,31,239,31,142,31,244,31,234,31,234,30,234,29,127,31,73,31,82,31,69,31,109,31,36,31,147,31,76,31,226,31,226,30,226,29,229,31,166,31,72,31,127,31,197,31,197,30,177,31,88,31,33,31,11,31,55,31,199,31,133,31,216,31,58,31,58,30,141,31,231,31,45,31,245,31,245,30,92,31,92,30,194,31,106,31,14,31,232,31,158,31,111,31,228,31,104,31,70,31,71,31,125,31,30,31,30,30,134,31,20,31,208,31,47,31,72,31,55,31,55,30,249,31,150,31,150,30,150,29,243,31,243,30,236,31,236,30,90,31,90,30,57,31,57,30,229,31,229,30,229,29,229,28,93,31,225,31,200,31,46,31,46,30,49,31,185,31,99,31,83,31,151,31,31,31,31,30,136,31,135,31,66,31,183,31,183,30,243,31,15,31,15,30,254,31,254,30,202,31,66,31,238,31,54,31,43,31,43,30,18,31,152,31,180,31,250,31,151,31,151,30,151,29,151,28,255,31,178,31,157,31,2,31,50,31,173,31,254,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
