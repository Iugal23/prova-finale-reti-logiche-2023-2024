-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_158 is
end project_tb_158;

architecture project_tb_arch_158 of project_tb_158 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 889;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (241,0,29,0,50,0,104,0,63,0,223,0,0,0,0,0,183,0,110,0,244,0,153,0,9,0,93,0,231,0,246,0,10,0,72,0,241,0,0,0,252,0,239,0,107,0,55,0,0,0,0,0,59,0,133,0,251,0,0,0,211,0,223,0,129,0,185,0,0,0,81,0,3,0,0,0,155,0,105,0,132,0,124,0,174,0,196,0,124,0,154,0,0,0,38,0,86,0,162,0,196,0,62,0,165,0,35,0,221,0,5,0,178,0,0,0,120,0,121,0,11,0,131,0,79,0,149,0,231,0,154,0,64,0,6,0,226,0,198,0,215,0,59,0,197,0,73,0,2,0,166,0,101,0,162,0,157,0,120,0,62,0,0,0,164,0,230,0,154,0,11,0,251,0,0,0,121,0,148,0,81,0,43,0,167,0,37,0,63,0,0,0,210,0,105,0,232,0,181,0,187,0,105,0,114,0,46,0,77,0,0,0,103,0,0,0,121,0,56,0,80,0,175,0,250,0,3,0,228,0,98,0,82,0,91,0,0,0,0,0,44,0,43,0,5,0,50,0,195,0,14,0,99,0,151,0,193,0,96,0,85,0,229,0,222,0,0,0,119,0,192,0,212,0,133,0,125,0,0,0,0,0,192,0,55,0,93,0,0,0,95,0,199,0,0,0,0,0,0,0,0,0,0,0,122,0,175,0,187,0,64,0,121,0,188,0,104,0,217,0,146,0,105,0,39,0,226,0,138,0,0,0,0,0,191,0,79,0,6,0,20,0,190,0,0,0,120,0,0,0,0,0,0,0,2,0,0,0,236,0,0,0,0,0,44,0,224,0,97,0,113,0,193,0,132,0,47,0,82,0,241,0,0,0,202,0,112,0,199,0,204,0,44,0,0,0,238,0,227,0,88,0,206,0,2,0,235,0,223,0,0,0,0,0,240,0,197,0,161,0,117,0,27,0,39,0,136,0,135,0,39,0,118,0,164,0,0,0,0,0,186,0,0,0,58,0,50,0,87,0,175,0,221,0,0,0,52,0,0,0,45,0,193,0,236,0,141,0,248,0,79,0,0,0,197,0,150,0,85,0,57,0,45,0,112,0,0,0,74,0,102,0,253,0,184,0,0,0,138,0,73,0,159,0,97,0,214,0,132,0,236,0,159,0,0,0,241,0,204,0,117,0,0,0,227,0,0,0,0,0,12,0,0,0,188,0,182,0,0,0,219,0,88,0,0,0,57,0,164,0,228,0,214,0,0,0,45,0,0,0,223,0,0,0,173,0,173,0,0,0,156,0,173,0,12,0,177,0,149,0,189,0,162,0,82,0,0,0,14,0,143,0,0,0,35,0,10,0,255,0,142,0,211,0,159,0,66,0,163,0,0,0,211,0,163,0,248,0,0,0,116,0,9,0,232,0,0,0,0,0,231,0,165,0,223,0,56,0,0,0,99,0,2,0,143,0,88,0,46,0,91,0,210,0,69,0,251,0,76,0,19,0,153,0,247,0,144,0,0,0,0,0,130,0,0,0,86,0,212,0,138,0,0,0,186,0,143,0,87,0,48,0,133,0,144,0,230,0,0,0,122,0,0,0,119,0,0,0,92,0,113,0,123,0,0,0,26,0,249,0,74,0,178,0,50,0,0,0,67,0,208,0,113,0,156,0,172,0,0,0,44,0,174,0,110,0,126,0,59,0,152,0,121,0,216,0,104,0,223,0,196,0,81,0,123,0,0,0,75,0,152,0,80,0,0,0,0,0,64,0,29,0,53,0,200,0,0,0,170,0,203,0,0,0,9,0,184,0,0,0,0,0,145,0,35,0,219,0,207,0,30,0,238,0,0,0,101,0,23,0,0,0,2,0,0,0,25,0,230,0,0,0,0,0,57,0,30,0,104,0,0,0,28,0,45,0,0,0,117,0,123,0,52,0,87,0,157,0,54,0,248,0,0,0,85,0,131,0,0,0,0,0,231,0,171,0,157,0,192,0,161,0,215,0,143,0,0,0,112,0,0,0,217,0,17,0,112,0,44,0,118,0,95,0,48,0,44,0,184,0,190,0,82,0,239,0,195,0,27,0,73,0,0,0,73,0,119,0,213,0,0,0,0,0,185,0,153,0,0,0,120,0,103,0,0,0,152,0,68,0,173,0,65,0,0,0,0,0,162,0,4,0,98,0,89,0,226,0,83,0,0,0,214,0,238,0,51,0,97,0,73,0,0,0,36,0,186,0,241,0,37,0,23,0,0,0,0,0,46,0,21,0,222,0,0,0,109,0,137,0,0,0,162,0,142,0,87,0,0,0,0,0,19,0,0,0,10,0,41,0,27,0,238,0,41,0,238,0,203,0,58,0,105,0,101,0,117,0,187,0,191,0,11,0,93,0,89,0,242,0,190,0,45,0,0,0,244,0,137,0,221,0,7,0,243,0,162,0,0,0,183,0,250,0,212,0,84,0,4,0,0,0,135,0,196,0,69,0,148,0,142,0,0,0,255,0,154,0,178,0,22,0,215,0,243,0,155,0,47,0,0,0,64,0,191,0,119,0,12,0,0,0,3,0,62,0,181,0,171,0,219,0,0,0,9,0,0,0,56,0,0,0,0,0,145,0,200,0,56,0,0,0,138,0,187,0,59,0,0,0,148,0,121,0,148,0,0,0,38,0,0,0,172,0,0,0,0,0,89,0,217,0,244,0,211,0,133,0,242,0,96,0,106,0,0,0,0,0,244,0,240,0,91,0,97,0,133,0,57,0,0,0,19,0,0,0,105,0,39,0,69,0,0,0,0,0,109,0,0,0,118,0,0,0,44,0,89,0,49,0,69,0,238,0,0,0,0,0,0,0,192,0,61,0,114,0,103,0,217,0,39,0,105,0,0,0,105,0,0,0,119,0,21,0,65,0,136,0,108,0,0,0,59,0,0,0,80,0,241,0,68,0,39,0,247,0,33,0,200,0,191,0,0,0,241,0,19,0,241,0,0,0,215,0,0,0,230,0,0,0,0,0,87,0,136,0,153,0,25,0,216,0,144,0,60,0,166,0,79,0,229,0,252,0,146,0,120,0,216,0,177,0,165,0,0,0,65,0,246,0,225,0,167,0,73,0,110,0,0,0,105,0,0,0,0,0,120,0,0,0,114,0,129,0,105,0,60,0,83,0,1,0,139,0,55,0,0,0,171,0,24,0,224,0,121,0,0,0,131,0,0,0,218,0,37,0,178,0,21,0,150,0,136,0,0,0,2,0,223,0,144,0,0,0,192,0,170,0,11,0,70,0,163,0,54,0,0,0,34,0,165,0,58,0,190,0,0,0,0,0,175,0,67,0,0,0,240,0,245,0,100,0,54,0,80,0,152,0,229,0,224,0,228,0,67,0,0,0,183,0,48,0,93,0,0,0,231,0,10,0,196,0,35,0,138,0,231,0,42,0,28,0,123,0,6,0,75,0,218,0,146,0,152,0,24,0,155,0,64,0,225,0,177,0,171,0,26,0,157,0,0,0,213,0,0,0,59,0,55,0,196,0,3,0,63,0,223,0,220,0,71,0,125,0,48,0,80,0,17,0,214,0,0,0,0,0,0,0,147,0,0,0,43,0,95,0,14,0,0,0,120,0,12,0,214,0,0,0,213,0,233,0,0,0,35,0,0,0,156,0,51,0,119,0,113,0,0,0,0,0,59,0,186,0,53,0,59,0,3,0,247,0,92,0,0,0,139,0,0,0,8,0,169,0,0,0,28,0,182,0,0,0,232,0,178,0,157,0,109,0,28,0,0,0,53,0,0,0,0,0,138,0,0,0,66,0,164,0,195,0,34,0,140,0,34,0,32,0,133,0,205,0,0,0,0,0,217,0,0,0,67,0,23,0,53,0,232,0,0,0,0,0,0,0,16,0,0,0,0,0,16,0,0,0,32,0,83,0,84,0,59,0,209,0,0,0,228,0,148,0,178,0,239,0,90,0,59,0,90,0,108,0,105,0,129,0,181,0,214,0,21,0,101,0,112,0,227,0);
signal scenario_full  : scenario_type := (241,31,29,31,50,31,104,31,63,31,223,31,223,30,223,29,183,31,110,31,244,31,153,31,9,31,93,31,231,31,246,31,10,31,72,31,241,31,241,30,252,31,239,31,107,31,55,31,55,30,55,29,59,31,133,31,251,31,251,30,211,31,223,31,129,31,185,31,185,30,81,31,3,31,3,30,155,31,105,31,132,31,124,31,174,31,196,31,124,31,154,31,154,30,38,31,86,31,162,31,196,31,62,31,165,31,35,31,221,31,5,31,178,31,178,30,120,31,121,31,11,31,131,31,79,31,149,31,231,31,154,31,64,31,6,31,226,31,198,31,215,31,59,31,197,31,73,31,2,31,166,31,101,31,162,31,157,31,120,31,62,31,62,30,164,31,230,31,154,31,11,31,251,31,251,30,121,31,148,31,81,31,43,31,167,31,37,31,63,31,63,30,210,31,105,31,232,31,181,31,187,31,105,31,114,31,46,31,77,31,77,30,103,31,103,30,121,31,56,31,80,31,175,31,250,31,3,31,228,31,98,31,82,31,91,31,91,30,91,29,44,31,43,31,5,31,50,31,195,31,14,31,99,31,151,31,193,31,96,31,85,31,229,31,222,31,222,30,119,31,192,31,212,31,133,31,125,31,125,30,125,29,192,31,55,31,93,31,93,30,95,31,199,31,199,30,199,29,199,28,199,27,199,26,122,31,175,31,187,31,64,31,121,31,188,31,104,31,217,31,146,31,105,31,39,31,226,31,138,31,138,30,138,29,191,31,79,31,6,31,20,31,190,31,190,30,120,31,120,30,120,29,120,28,2,31,2,30,236,31,236,30,236,29,44,31,224,31,97,31,113,31,193,31,132,31,47,31,82,31,241,31,241,30,202,31,112,31,199,31,204,31,44,31,44,30,238,31,227,31,88,31,206,31,2,31,235,31,223,31,223,30,223,29,240,31,197,31,161,31,117,31,27,31,39,31,136,31,135,31,39,31,118,31,164,31,164,30,164,29,186,31,186,30,58,31,50,31,87,31,175,31,221,31,221,30,52,31,52,30,45,31,193,31,236,31,141,31,248,31,79,31,79,30,197,31,150,31,85,31,57,31,45,31,112,31,112,30,74,31,102,31,253,31,184,31,184,30,138,31,73,31,159,31,97,31,214,31,132,31,236,31,159,31,159,30,241,31,204,31,117,31,117,30,227,31,227,30,227,29,12,31,12,30,188,31,182,31,182,30,219,31,88,31,88,30,57,31,164,31,228,31,214,31,214,30,45,31,45,30,223,31,223,30,173,31,173,31,173,30,156,31,173,31,12,31,177,31,149,31,189,31,162,31,82,31,82,30,14,31,143,31,143,30,35,31,10,31,255,31,142,31,211,31,159,31,66,31,163,31,163,30,211,31,163,31,248,31,248,30,116,31,9,31,232,31,232,30,232,29,231,31,165,31,223,31,56,31,56,30,99,31,2,31,143,31,88,31,46,31,91,31,210,31,69,31,251,31,76,31,19,31,153,31,247,31,144,31,144,30,144,29,130,31,130,30,86,31,212,31,138,31,138,30,186,31,143,31,87,31,48,31,133,31,144,31,230,31,230,30,122,31,122,30,119,31,119,30,92,31,113,31,123,31,123,30,26,31,249,31,74,31,178,31,50,31,50,30,67,31,208,31,113,31,156,31,172,31,172,30,44,31,174,31,110,31,126,31,59,31,152,31,121,31,216,31,104,31,223,31,196,31,81,31,123,31,123,30,75,31,152,31,80,31,80,30,80,29,64,31,29,31,53,31,200,31,200,30,170,31,203,31,203,30,9,31,184,31,184,30,184,29,145,31,35,31,219,31,207,31,30,31,238,31,238,30,101,31,23,31,23,30,2,31,2,30,25,31,230,31,230,30,230,29,57,31,30,31,104,31,104,30,28,31,45,31,45,30,117,31,123,31,52,31,87,31,157,31,54,31,248,31,248,30,85,31,131,31,131,30,131,29,231,31,171,31,157,31,192,31,161,31,215,31,143,31,143,30,112,31,112,30,217,31,17,31,112,31,44,31,118,31,95,31,48,31,44,31,184,31,190,31,82,31,239,31,195,31,27,31,73,31,73,30,73,31,119,31,213,31,213,30,213,29,185,31,153,31,153,30,120,31,103,31,103,30,152,31,68,31,173,31,65,31,65,30,65,29,162,31,4,31,98,31,89,31,226,31,83,31,83,30,214,31,238,31,51,31,97,31,73,31,73,30,36,31,186,31,241,31,37,31,23,31,23,30,23,29,46,31,21,31,222,31,222,30,109,31,137,31,137,30,162,31,142,31,87,31,87,30,87,29,19,31,19,30,10,31,41,31,27,31,238,31,41,31,238,31,203,31,58,31,105,31,101,31,117,31,187,31,191,31,11,31,93,31,89,31,242,31,190,31,45,31,45,30,244,31,137,31,221,31,7,31,243,31,162,31,162,30,183,31,250,31,212,31,84,31,4,31,4,30,135,31,196,31,69,31,148,31,142,31,142,30,255,31,154,31,178,31,22,31,215,31,243,31,155,31,47,31,47,30,64,31,191,31,119,31,12,31,12,30,3,31,62,31,181,31,171,31,219,31,219,30,9,31,9,30,56,31,56,30,56,29,145,31,200,31,56,31,56,30,138,31,187,31,59,31,59,30,148,31,121,31,148,31,148,30,38,31,38,30,172,31,172,30,172,29,89,31,217,31,244,31,211,31,133,31,242,31,96,31,106,31,106,30,106,29,244,31,240,31,91,31,97,31,133,31,57,31,57,30,19,31,19,30,105,31,39,31,69,31,69,30,69,29,109,31,109,30,118,31,118,30,44,31,89,31,49,31,69,31,238,31,238,30,238,29,238,28,192,31,61,31,114,31,103,31,217,31,39,31,105,31,105,30,105,31,105,30,119,31,21,31,65,31,136,31,108,31,108,30,59,31,59,30,80,31,241,31,68,31,39,31,247,31,33,31,200,31,191,31,191,30,241,31,19,31,241,31,241,30,215,31,215,30,230,31,230,30,230,29,87,31,136,31,153,31,25,31,216,31,144,31,60,31,166,31,79,31,229,31,252,31,146,31,120,31,216,31,177,31,165,31,165,30,65,31,246,31,225,31,167,31,73,31,110,31,110,30,105,31,105,30,105,29,120,31,120,30,114,31,129,31,105,31,60,31,83,31,1,31,139,31,55,31,55,30,171,31,24,31,224,31,121,31,121,30,131,31,131,30,218,31,37,31,178,31,21,31,150,31,136,31,136,30,2,31,223,31,144,31,144,30,192,31,170,31,11,31,70,31,163,31,54,31,54,30,34,31,165,31,58,31,190,31,190,30,190,29,175,31,67,31,67,30,240,31,245,31,100,31,54,31,80,31,152,31,229,31,224,31,228,31,67,31,67,30,183,31,48,31,93,31,93,30,231,31,10,31,196,31,35,31,138,31,231,31,42,31,28,31,123,31,6,31,75,31,218,31,146,31,152,31,24,31,155,31,64,31,225,31,177,31,171,31,26,31,157,31,157,30,213,31,213,30,59,31,55,31,196,31,3,31,63,31,223,31,220,31,71,31,125,31,48,31,80,31,17,31,214,31,214,30,214,29,214,28,147,31,147,30,43,31,95,31,14,31,14,30,120,31,12,31,214,31,214,30,213,31,233,31,233,30,35,31,35,30,156,31,51,31,119,31,113,31,113,30,113,29,59,31,186,31,53,31,59,31,3,31,247,31,92,31,92,30,139,31,139,30,8,31,169,31,169,30,28,31,182,31,182,30,232,31,178,31,157,31,109,31,28,31,28,30,53,31,53,30,53,29,138,31,138,30,66,31,164,31,195,31,34,31,140,31,34,31,32,31,133,31,205,31,205,30,205,29,217,31,217,30,67,31,23,31,53,31,232,31,232,30,232,29,232,28,16,31,16,30,16,29,16,31,16,30,32,31,83,31,84,31,59,31,209,31,209,30,228,31,148,31,178,31,239,31,90,31,59,31,90,31,108,31,105,31,129,31,181,31,214,31,21,31,101,31,112,31,227,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
