-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 804;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (223,0,111,0,106,0,62,0,0,0,0,0,30,0,234,0,0,0,229,0,29,0,84,0,221,0,62,0,0,0,10,0,84,0,17,0,204,0,178,0,115,0,122,0,0,0,159,0,90,0,0,0,83,0,129,0,80,0,197,0,180,0,0,0,175,0,160,0,0,0,55,0,104,0,61,0,144,0,76,0,0,0,81,0,0,0,0,0,47,0,180,0,20,0,192,0,211,0,154,0,74,0,246,0,188,0,10,0,0,0,246,0,128,0,58,0,72,0,0,0,47,0,255,0,186,0,54,0,0,0,0,0,191,0,166,0,138,0,247,0,36,0,189,0,0,0,56,0,35,0,106,0,126,0,0,0,208,0,199,0,0,0,32,0,151,0,0,0,243,0,156,0,0,0,36,0,2,0,194,0,229,0,0,0,254,0,12,0,73,0,86,0,233,0,10,0,235,0,239,0,39,0,238,0,0,0,163,0,2,0,188,0,0,0,76,0,0,0,255,0,42,0,239,0,228,0,0,0,210,0,0,0,131,0,107,0,222,0,250,0,34,0,206,0,0,0,147,0,174,0,18,0,0,0,0,0,18,0,131,0,115,0,235,0,220,0,30,0,100,0,180,0,26,0,238,0,156,0,173,0,203,0,2,0,111,0,177,0,6,0,238,0,127,0,149,0,145,0,11,0,214,0,207,0,159,0,27,0,0,0,238,0,92,0,23,0,0,0,72,0,223,0,0,0,182,0,48,0,198,0,0,0,0,0,33,0,140,0,0,0,16,0,241,0,151,0,248,0,22,0,47,0,247,0,42,0,76,0,246,0,0,0,62,0,161,0,67,0,135,0,164,0,180,0,106,0,240,0,84,0,0,0,151,0,97,0,235,0,121,0,117,0,4,0,0,0,48,0,210,0,234,0,232,0,6,0,167,0,83,0,110,0,89,0,224,0,0,0,1,0,135,0,100,0,146,0,193,0,12,0,130,0,39,0,217,0,6,0,209,0,126,0,0,0,125,0,163,0,169,0,69,0,165,0,49,0,167,0,33,0,54,0,43,0,121,0,156,0,16,0,94,0,0,0,99,0,0,0,88,0,116,0,209,0,204,0,229,0,173,0,0,0,200,0,0,0,116,0,203,0,0,0,0,0,0,0,0,0,63,0,191,0,80,0,237,0,0,0,110,0,6,0,0,0,1,0,0,0,0,0,0,0,123,0,30,0,154,0,200,0,106,0,215,0,0,0,9,0,182,0,225,0,235,0,89,0,27,0,0,0,0,0,210,0,130,0,233,0,92,0,0,0,253,0,86,0,164,0,255,0,242,0,60,0,231,0,0,0,232,0,164,0,71,0,13,0,166,0,0,0,54,0,105,0,132,0,222,0,185,0,132,0,242,0,0,0,5,0,149,0,0,0,165,0,0,0,22,0,227,0,105,0,0,0,23,0,111,0,70,0,215,0,0,0,239,0,161,0,109,0,29,0,235,0,214,0,44,0,231,0,227,0,213,0,241,0,0,0,215,0,136,0,249,0,42,0,234,0,195,0,22,0,31,0,0,0,35,0,119,0,0,0,29,0,207,0,11,0,186,0,0,0,4,0,0,0,177,0,248,0,49,0,0,0,210,0,94,0,241,0,0,0,0,0,0,0,250,0,0,0,31,0,115,0,186,0,208,0,58,0,244,0,109,0,41,0,89,0,113,0,69,0,0,0,180,0,69,0,160,0,82,0,145,0,88,0,102,0,157,0,129,0,203,0,120,0,111,0,230,0,151,0,135,0,216,0,0,0,43,0,53,0,0,0,199,0,156,0,209,0,134,0,170,0,31,0,255,0,79,0,118,0,250,0,137,0,206,0,53,0,30,0,0,0,89,0,0,0,79,0,0,0,216,0,0,0,51,0,0,0,126,0,48,0,216,0,0,0,200,0,30,0,46,0,255,0,118,0,240,0,6,0,175,0,0,0,207,0,154,0,48,0,242,0,103,0,30,0,135,0,191,0,195,0,4,0,0,0,72,0,193,0,87,0,1,0,44,0,36,0,253,0,124,0,0,0,4,0,69,0,29,0,29,0,192,0,68,0,150,0,173,0,0,0,0,0,23,0,50,0,224,0,83,0,208,0,66,0,6,0,147,0,75,0,233,0,0,0,0,0,59,0,155,0,73,0,236,0,44,0,0,0,0,0,159,0,0,0,0,0,25,0,0,0,48,0,15,0,50,0,157,0,213,0,163,0,165,0,34,0,0,0,230,0,221,0,187,0,106,0,181,0,0,0,252,0,216,0,52,0,3,0,142,0,97,0,69,0,108,0,216,0,157,0,234,0,0,0,0,0,82,0,173,0,187,0,67,0,234,0,94,0,180,0,232,0,151,0,194,0,207,0,208,0,0,0,158,0,0,0,206,0,94,0,195,0,208,0,0,0,204,0,214,0,236,0,0,0,0,0,199,0,0,0,178,0,18,0,152,0,178,0,169,0,51,0,0,0,221,0,152,0,93,0,243,0,131,0,53,0,1,0,91,0,0,0,135,0,0,0,17,0,0,0,0,0,43,0,0,0,55,0,133,0,0,0,0,0,150,0,0,0,208,0,98,0,219,0,187,0,131,0,48,0,26,0,169,0,28,0,193,0,213,0,81,0,123,0,0,0,183,0,180,0,218,0,65,0,43,0,201,0,18,0,3,0,254,0,118,0,0,0,235,0,66,0,150,0,9,0,232,0,163,0,10,0,129,0,115,0,64,0,23,0,0,0,27,0,227,0,55,0,178,0,71,0,86,0,0,0,135,0,91,0,144,0,104,0,155,0,7,0,207,0,137,0,180,0,0,0,0,0,0,0,161,0,0,0,52,0,74,0,137,0,21,0,27,0,193,0,198,0,131,0,120,0,166,0,213,0,0,0,170,0,207,0,0,0,164,0,195,0,252,0,0,0,9,0,187,0,247,0,247,0,0,0,89,0,96,0,160,0,37,0,0,0,167,0,189,0,38,0,162,0,0,0,231,0,26,0,0,0,252,0,91,0,95,0,203,0,166,0,32,0,148,0,4,0,135,0,183,0,28,0,54,0,161,0,127,0,0,0,7,0,141,0,41,0,178,0,0,0,0,0,165,0,12,0,0,0,1,0,75,0,196,0,0,0,0,0,61,0,216,0,155,0,165,0,183,0,59,0,0,0,0,0,76,0,0,0,127,0,21,0,0,0,64,0,224,0,129,0,223,0,107,0,248,0,16,0,46,0,43,0,208,0,244,0,132,0,217,0,34,0,98,0,151,0,208,0,62,0,65,0,6,0,168,0,155,0,37,0,183,0,128,0,232,0,45,0,19,0,25,0,201,0,49,0,76,0,0,0,64,0,84,0,68,0,32,0,80,0,202,0,162,0,86,0,41,0,0,0,92,0,172,0,39,0,0,0,246,0,247,0,113,0,0,0,0,0,150,0,60,0,229,0,0,0,158,0,123,0,215,0,163,0,203,0,236,0,108,0,6,0,186,0,15,0,53,0,21,0,0,0,0,0,177,0,56,0,7,0,37,0,93,0,175,0,137,0,132,0,209,0,249,0,76,0,0,0,119,0,72,0,105,0,131,0,15,0,115,0,0,0,229,0,202,0,92,0,107,0,136,0,252,0,145,0);
signal scenario_full  : scenario_type := (223,31,111,31,106,31,62,31,62,30,62,29,30,31,234,31,234,30,229,31,29,31,84,31,221,31,62,31,62,30,10,31,84,31,17,31,204,31,178,31,115,31,122,31,122,30,159,31,90,31,90,30,83,31,129,31,80,31,197,31,180,31,180,30,175,31,160,31,160,30,55,31,104,31,61,31,144,31,76,31,76,30,81,31,81,30,81,29,47,31,180,31,20,31,192,31,211,31,154,31,74,31,246,31,188,31,10,31,10,30,246,31,128,31,58,31,72,31,72,30,47,31,255,31,186,31,54,31,54,30,54,29,191,31,166,31,138,31,247,31,36,31,189,31,189,30,56,31,35,31,106,31,126,31,126,30,208,31,199,31,199,30,32,31,151,31,151,30,243,31,156,31,156,30,36,31,2,31,194,31,229,31,229,30,254,31,12,31,73,31,86,31,233,31,10,31,235,31,239,31,39,31,238,31,238,30,163,31,2,31,188,31,188,30,76,31,76,30,255,31,42,31,239,31,228,31,228,30,210,31,210,30,131,31,107,31,222,31,250,31,34,31,206,31,206,30,147,31,174,31,18,31,18,30,18,29,18,31,131,31,115,31,235,31,220,31,30,31,100,31,180,31,26,31,238,31,156,31,173,31,203,31,2,31,111,31,177,31,6,31,238,31,127,31,149,31,145,31,11,31,214,31,207,31,159,31,27,31,27,30,238,31,92,31,23,31,23,30,72,31,223,31,223,30,182,31,48,31,198,31,198,30,198,29,33,31,140,31,140,30,16,31,241,31,151,31,248,31,22,31,47,31,247,31,42,31,76,31,246,31,246,30,62,31,161,31,67,31,135,31,164,31,180,31,106,31,240,31,84,31,84,30,151,31,97,31,235,31,121,31,117,31,4,31,4,30,48,31,210,31,234,31,232,31,6,31,167,31,83,31,110,31,89,31,224,31,224,30,1,31,135,31,100,31,146,31,193,31,12,31,130,31,39,31,217,31,6,31,209,31,126,31,126,30,125,31,163,31,169,31,69,31,165,31,49,31,167,31,33,31,54,31,43,31,121,31,156,31,16,31,94,31,94,30,99,31,99,30,88,31,116,31,209,31,204,31,229,31,173,31,173,30,200,31,200,30,116,31,203,31,203,30,203,29,203,28,203,27,63,31,191,31,80,31,237,31,237,30,110,31,6,31,6,30,1,31,1,30,1,29,1,28,123,31,30,31,154,31,200,31,106,31,215,31,215,30,9,31,182,31,225,31,235,31,89,31,27,31,27,30,27,29,210,31,130,31,233,31,92,31,92,30,253,31,86,31,164,31,255,31,242,31,60,31,231,31,231,30,232,31,164,31,71,31,13,31,166,31,166,30,54,31,105,31,132,31,222,31,185,31,132,31,242,31,242,30,5,31,149,31,149,30,165,31,165,30,22,31,227,31,105,31,105,30,23,31,111,31,70,31,215,31,215,30,239,31,161,31,109,31,29,31,235,31,214,31,44,31,231,31,227,31,213,31,241,31,241,30,215,31,136,31,249,31,42,31,234,31,195,31,22,31,31,31,31,30,35,31,119,31,119,30,29,31,207,31,11,31,186,31,186,30,4,31,4,30,177,31,248,31,49,31,49,30,210,31,94,31,241,31,241,30,241,29,241,28,250,31,250,30,31,31,115,31,186,31,208,31,58,31,244,31,109,31,41,31,89,31,113,31,69,31,69,30,180,31,69,31,160,31,82,31,145,31,88,31,102,31,157,31,129,31,203,31,120,31,111,31,230,31,151,31,135,31,216,31,216,30,43,31,53,31,53,30,199,31,156,31,209,31,134,31,170,31,31,31,255,31,79,31,118,31,250,31,137,31,206,31,53,31,30,31,30,30,89,31,89,30,79,31,79,30,216,31,216,30,51,31,51,30,126,31,48,31,216,31,216,30,200,31,30,31,46,31,255,31,118,31,240,31,6,31,175,31,175,30,207,31,154,31,48,31,242,31,103,31,30,31,135,31,191,31,195,31,4,31,4,30,72,31,193,31,87,31,1,31,44,31,36,31,253,31,124,31,124,30,4,31,69,31,29,31,29,31,192,31,68,31,150,31,173,31,173,30,173,29,23,31,50,31,224,31,83,31,208,31,66,31,6,31,147,31,75,31,233,31,233,30,233,29,59,31,155,31,73,31,236,31,44,31,44,30,44,29,159,31,159,30,159,29,25,31,25,30,48,31,15,31,50,31,157,31,213,31,163,31,165,31,34,31,34,30,230,31,221,31,187,31,106,31,181,31,181,30,252,31,216,31,52,31,3,31,142,31,97,31,69,31,108,31,216,31,157,31,234,31,234,30,234,29,82,31,173,31,187,31,67,31,234,31,94,31,180,31,232,31,151,31,194,31,207,31,208,31,208,30,158,31,158,30,206,31,94,31,195,31,208,31,208,30,204,31,214,31,236,31,236,30,236,29,199,31,199,30,178,31,18,31,152,31,178,31,169,31,51,31,51,30,221,31,152,31,93,31,243,31,131,31,53,31,1,31,91,31,91,30,135,31,135,30,17,31,17,30,17,29,43,31,43,30,55,31,133,31,133,30,133,29,150,31,150,30,208,31,98,31,219,31,187,31,131,31,48,31,26,31,169,31,28,31,193,31,213,31,81,31,123,31,123,30,183,31,180,31,218,31,65,31,43,31,201,31,18,31,3,31,254,31,118,31,118,30,235,31,66,31,150,31,9,31,232,31,163,31,10,31,129,31,115,31,64,31,23,31,23,30,27,31,227,31,55,31,178,31,71,31,86,31,86,30,135,31,91,31,144,31,104,31,155,31,7,31,207,31,137,31,180,31,180,30,180,29,180,28,161,31,161,30,52,31,74,31,137,31,21,31,27,31,193,31,198,31,131,31,120,31,166,31,213,31,213,30,170,31,207,31,207,30,164,31,195,31,252,31,252,30,9,31,187,31,247,31,247,31,247,30,89,31,96,31,160,31,37,31,37,30,167,31,189,31,38,31,162,31,162,30,231,31,26,31,26,30,252,31,91,31,95,31,203,31,166,31,32,31,148,31,4,31,135,31,183,31,28,31,54,31,161,31,127,31,127,30,7,31,141,31,41,31,178,31,178,30,178,29,165,31,12,31,12,30,1,31,75,31,196,31,196,30,196,29,61,31,216,31,155,31,165,31,183,31,59,31,59,30,59,29,76,31,76,30,127,31,21,31,21,30,64,31,224,31,129,31,223,31,107,31,248,31,16,31,46,31,43,31,208,31,244,31,132,31,217,31,34,31,98,31,151,31,208,31,62,31,65,31,6,31,168,31,155,31,37,31,183,31,128,31,232,31,45,31,19,31,25,31,201,31,49,31,76,31,76,30,64,31,84,31,68,31,32,31,80,31,202,31,162,31,86,31,41,31,41,30,92,31,172,31,39,31,39,30,246,31,247,31,113,31,113,30,113,29,150,31,60,31,229,31,229,30,158,31,123,31,215,31,163,31,203,31,236,31,108,31,6,31,186,31,15,31,53,31,21,31,21,30,21,29,177,31,56,31,7,31,37,31,93,31,175,31,137,31,132,31,209,31,249,31,76,31,76,30,119,31,72,31,105,31,131,31,15,31,115,31,115,30,229,31,202,31,92,31,107,31,136,31,252,31,145,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
