-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 955;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (209,0,33,0,157,0,0,0,0,0,55,0,92,0,44,0,0,0,184,0,91,0,34,0,33,0,40,0,133,0,189,0,65,0,97,0,43,0,143,0,64,0,232,0,191,0,8,0,0,0,141,0,212,0,146,0,220,0,12,0,236,0,131,0,117,0,185,0,204,0,0,0,78,0,4,0,143,0,84,0,244,0,0,0,0,0,10,0,88,0,93,0,0,0,131,0,148,0,184,0,43,0,125,0,3,0,44,0,101,0,118,0,157,0,0,0,19,0,21,0,0,0,211,0,62,0,196,0,98,0,195,0,209,0,198,0,73,0,0,0,226,0,16,0,169,0,243,0,57,0,140,0,232,0,200,0,21,0,6,0,13,0,17,0,33,0,231,0,71,0,44,0,0,0,253,0,238,0,134,0,62,0,152,0,205,0,0,0,0,0,75,0,80,0,247,0,57,0,76,0,40,0,0,0,55,0,189,0,239,0,9,0,143,0,160,0,213,0,64,0,158,0,206,0,130,0,101,0,224,0,98,0,0,0,234,0,42,0,130,0,201,0,0,0,128,0,0,0,91,0,0,0,113,0,89,0,105,0,0,0,20,0,165,0,95,0,138,0,0,0,71,0,1,0,190,0,48,0,255,0,52,0,67,0,102,0,0,0,15,0,67,0,94,0,193,0,46,0,134,0,250,0,68,0,0,0,13,0,150,0,0,0,203,0,0,0,3,0,73,0,236,0,216,0,0,0,0,0,78,0,28,0,206,0,0,0,66,0,0,0,124,0,206,0,227,0,30,0,62,0,85,0,61,0,0,0,218,0,52,0,0,0,24,0,0,0,104,0,0,0,164,0,168,0,159,0,177,0,0,0,112,0,22,0,189,0,0,0,188,0,146,0,0,0,159,0,182,0,162,0,94,0,49,0,0,0,157,0,137,0,0,0,0,0,219,0,102,0,85,0,54,0,0,0,161,0,157,0,0,0,146,0,105,0,217,0,6,0,212,0,57,0,55,0,219,0,22,0,243,0,147,0,71,0,113,0,218,0,124,0,0,0,171,0,250,0,112,0,203,0,222,0,133,0,141,0,44,0,227,0,42,0,50,0,244,0,192,0,95,0,212,0,106,0,0,0,1,0,21,0,0,0,98,0,0,0,220,0,232,0,157,0,0,0,54,0,142,0,0,0,235,0,24,0,59,0,185,0,0,0,61,0,216,0,201,0,0,0,137,0,0,0,0,0,64,0,179,0,240,0,250,0,7,0,167,0,232,0,242,0,58,0,154,0,56,0,0,0,85,0,2,0,138,0,104,0,205,0,155,0,253,0,199,0,232,0,68,0,0,0,38,0,0,0,0,0,4,0,106,0,205,0,0,0,0,0,247,0,203,0,127,0,95,0,111,0,188,0,4,0,243,0,90,0,144,0,169,0,140,0,0,0,230,0,193,0,162,0,236,0,79,0,0,0,11,0,143,0,0,0,42,0,0,0,0,0,53,0,133,0,189,0,74,0,81,0,0,0,76,0,66,0,232,0,173,0,0,0,0,0,165,0,196,0,0,0,231,0,55,0,45,0,124,0,0,0,0,0,21,0,95,0,61,0,60,0,58,0,239,0,249,0,104,0,0,0,147,0,150,0,15,0,246,0,0,0,104,0,26,0,235,0,4,0,64,0,247,0,224,0,0,0,198,0,55,0,185,0,83,0,106,0,240,0,166,0,0,0,105,0,25,0,41,0,105,0,213,0,71,0,100,0,251,0,0,0,0,0,86,0,3,0,0,0,0,0,160,0,209,0,0,0,0,0,70,0,196,0,45,0,0,0,39,0,1,0,240,0,192,0,0,0,0,0,134,0,149,0,28,0,236,0,42,0,145,0,100,0,29,0,22,0,229,0,196,0,74,0,152,0,184,0,5,0,0,0,47,0,113,0,55,0,109,0,0,0,91,0,129,0,22,0,23,0,149,0,156,0,168,0,218,0,0,0,0,0,41,0,99,0,0,0,254,0,0,0,132,0,123,0,249,0,0,0,0,0,106,0,218,0,113,0,0,0,29,0,186,0,70,0,88,0,146,0,0,0,0,0,180,0,19,0,0,0,228,0,148,0,61,0,152,0,183,0,52,0,243,0,154,0,180,0,23,0,0,0,163,0,224,0,159,0,202,0,89,0,222,0,130,0,158,0,110,0,110,0,169,0,75,0,144,0,201,0,0,0,69,0,107,0,245,0,0,0,152,0,219,0,168,0,0,0,11,0,113,0,43,0,189,0,156,0,166,0,191,0,0,0,56,0,158,0,0,0,28,0,96,0,45,0,83,0,0,0,241,0,0,0,106,0,0,0,197,0,115,0,209,0,0,0,0,0,67,0,240,0,65,0,160,0,61,0,183,0,136,0,0,0,83,0,15,0,66,0,51,0,0,0,6,0,108,0,31,0,90,0,88,0,83,0,45,0,0,0,0,0,0,0,0,0,227,0,0,0,12,0,69,0,151,0,57,0,65,0,187,0,0,0,9,0,72,0,172,0,48,0,0,0,195,0,150,0,52,0,245,0,37,0,19,0,156,0,241,0,204,0,107,0,95,0,27,0,80,0,0,0,36,0,191,0,160,0,224,0,37,0,235,0,112,0,104,0,107,0,39,0,86,0,0,0,204,0,121,0,124,0,52,0,189,0,104,0,0,0,25,0,78,0,170,0,0,0,0,0,113,0,170,0,0,0,124,0,167,0,210,0,195,0,247,0,95,0,14,0,231,0,120,0,141,0,61,0,2,0,237,0,154,0,89,0,0,0,8,0,243,0,4,0,0,0,23,0,19,0,0,0,0,0,192,0,29,0,228,0,234,0,25,0,209,0,35,0,56,0,7,0,160,0,126,0,186,0,47,0,93,0,93,0,255,0,187,0,210,0,21,0,119,0,5,0,129,0,0,0,98,0,16,0,215,0,177,0,157,0,0,0,0,0,59,0,0,0,21,0,90,0,164,0,61,0,231,0,120,0,229,0,233,0,54,0,116,0,0,0,208,0,6,0,250,0,94,0,22,0,190,0,0,0,92,0,0,0,17,0,176,0,146,0,240,0,53,0,37,0,110,0,205,0,222,0,242,0,173,0,15,0,168,0,137,0,0,0,227,0,34,0,107,0,230,0,0,0,85,0,0,0,91,0,78,0,136,0,207,0,69,0,116,0,28,0,107,0,0,0,191,0,78,0,62,0,108,0,47,0,120,0,101,0,42,0,205,0,111,0,0,0,0,0,177,0,79,0,0,0,38,0,215,0,0,0,205,0,22,0,0,0,89,0,209,0,153,0,0,0,142,0,97,0,220,0,205,0,167,0,247,0,43,0,78,0,32,0,154,0,46,0,191,0,0,0,0,0,228,0,0,0,0,0,54,0,119,0,141,0,103,0,193,0,0,0,199,0,120,0,250,0,7,0,0,0,80,0,49,0,24,0,0,0,36,0,61,0,0,0,53,0,180,0,0,0,202,0,85,0,172,0,63,0,117,0,8,0,122,0,182,0,118,0,0,0,171,0,0,0,192,0,253,0,147,0,147,0,70,0,99,0,36,0,6,0,228,0,97,0,215,0,0,0,43,0,94,0,148,0,134,0,152,0,225,0,8,0,10,0,110,0,65,0,151,0,145,0,77,0,251,0,83,0,218,0,92,0,62,0,206,0,62,0,255,0,127,0,124,0,0,0,225,0,17,0,196,0,166,0,88,0,201,0,251,0,39,0,222,0,205,0,142,0,0,0,80,0,74,0,55,0,92,0,34,0,31,0,165,0,0,0,133,0,0,0,100,0,68,0,11,0,0,0,80,0,0,0,88,0,207,0,134,0,204,0,61,0,92,0,98,0,163,0,252,0,36,0,0,0,0,0,42,0,124,0,0,0,196,0,50,0,29,0,195,0,245,0,228,0,0,0,216,0,10,0,186,0,0,0,111,0,49,0,37,0,200,0,242,0,58,0,0,0,0,0,0,0,6,0,151,0,0,0,141,0,141,0,45,0,33,0,200,0,143,0,0,0,49,0,166,0,170,0,237,0,211,0,184,0,7,0,0,0,255,0,114,0,155,0,90,0,151,0,131,0,131,0,151,0,0,0,96,0,159,0,248,0,219,0,0,0,129,0,168,0,220,0,138,0,166,0,187,0,108,0,51,0,176,0,22,0,180,0,75,0,82,0,0,0,221,0,251,0,181,0,26,0,104,0,0,0,0,0,216,0,103,0,234,0,82,0,159,0,31,0,133,0,50,0,230,0,91,0,46,0,38,0,65,0,0,0,207,0,0,0,106,0,0,0,120,0,0,0,88,0);
signal scenario_full  : scenario_type := (209,31,33,31,157,31,157,30,157,29,55,31,92,31,44,31,44,30,184,31,91,31,34,31,33,31,40,31,133,31,189,31,65,31,97,31,43,31,143,31,64,31,232,31,191,31,8,31,8,30,141,31,212,31,146,31,220,31,12,31,236,31,131,31,117,31,185,31,204,31,204,30,78,31,4,31,143,31,84,31,244,31,244,30,244,29,10,31,88,31,93,31,93,30,131,31,148,31,184,31,43,31,125,31,3,31,44,31,101,31,118,31,157,31,157,30,19,31,21,31,21,30,211,31,62,31,196,31,98,31,195,31,209,31,198,31,73,31,73,30,226,31,16,31,169,31,243,31,57,31,140,31,232,31,200,31,21,31,6,31,13,31,17,31,33,31,231,31,71,31,44,31,44,30,253,31,238,31,134,31,62,31,152,31,205,31,205,30,205,29,75,31,80,31,247,31,57,31,76,31,40,31,40,30,55,31,189,31,239,31,9,31,143,31,160,31,213,31,64,31,158,31,206,31,130,31,101,31,224,31,98,31,98,30,234,31,42,31,130,31,201,31,201,30,128,31,128,30,91,31,91,30,113,31,89,31,105,31,105,30,20,31,165,31,95,31,138,31,138,30,71,31,1,31,190,31,48,31,255,31,52,31,67,31,102,31,102,30,15,31,67,31,94,31,193,31,46,31,134,31,250,31,68,31,68,30,13,31,150,31,150,30,203,31,203,30,3,31,73,31,236,31,216,31,216,30,216,29,78,31,28,31,206,31,206,30,66,31,66,30,124,31,206,31,227,31,30,31,62,31,85,31,61,31,61,30,218,31,52,31,52,30,24,31,24,30,104,31,104,30,164,31,168,31,159,31,177,31,177,30,112,31,22,31,189,31,189,30,188,31,146,31,146,30,159,31,182,31,162,31,94,31,49,31,49,30,157,31,137,31,137,30,137,29,219,31,102,31,85,31,54,31,54,30,161,31,157,31,157,30,146,31,105,31,217,31,6,31,212,31,57,31,55,31,219,31,22,31,243,31,147,31,71,31,113,31,218,31,124,31,124,30,171,31,250,31,112,31,203,31,222,31,133,31,141,31,44,31,227,31,42,31,50,31,244,31,192,31,95,31,212,31,106,31,106,30,1,31,21,31,21,30,98,31,98,30,220,31,232,31,157,31,157,30,54,31,142,31,142,30,235,31,24,31,59,31,185,31,185,30,61,31,216,31,201,31,201,30,137,31,137,30,137,29,64,31,179,31,240,31,250,31,7,31,167,31,232,31,242,31,58,31,154,31,56,31,56,30,85,31,2,31,138,31,104,31,205,31,155,31,253,31,199,31,232,31,68,31,68,30,38,31,38,30,38,29,4,31,106,31,205,31,205,30,205,29,247,31,203,31,127,31,95,31,111,31,188,31,4,31,243,31,90,31,144,31,169,31,140,31,140,30,230,31,193,31,162,31,236,31,79,31,79,30,11,31,143,31,143,30,42,31,42,30,42,29,53,31,133,31,189,31,74,31,81,31,81,30,76,31,66,31,232,31,173,31,173,30,173,29,165,31,196,31,196,30,231,31,55,31,45,31,124,31,124,30,124,29,21,31,95,31,61,31,60,31,58,31,239,31,249,31,104,31,104,30,147,31,150,31,15,31,246,31,246,30,104,31,26,31,235,31,4,31,64,31,247,31,224,31,224,30,198,31,55,31,185,31,83,31,106,31,240,31,166,31,166,30,105,31,25,31,41,31,105,31,213,31,71,31,100,31,251,31,251,30,251,29,86,31,3,31,3,30,3,29,160,31,209,31,209,30,209,29,70,31,196,31,45,31,45,30,39,31,1,31,240,31,192,31,192,30,192,29,134,31,149,31,28,31,236,31,42,31,145,31,100,31,29,31,22,31,229,31,196,31,74,31,152,31,184,31,5,31,5,30,47,31,113,31,55,31,109,31,109,30,91,31,129,31,22,31,23,31,149,31,156,31,168,31,218,31,218,30,218,29,41,31,99,31,99,30,254,31,254,30,132,31,123,31,249,31,249,30,249,29,106,31,218,31,113,31,113,30,29,31,186,31,70,31,88,31,146,31,146,30,146,29,180,31,19,31,19,30,228,31,148,31,61,31,152,31,183,31,52,31,243,31,154,31,180,31,23,31,23,30,163,31,224,31,159,31,202,31,89,31,222,31,130,31,158,31,110,31,110,31,169,31,75,31,144,31,201,31,201,30,69,31,107,31,245,31,245,30,152,31,219,31,168,31,168,30,11,31,113,31,43,31,189,31,156,31,166,31,191,31,191,30,56,31,158,31,158,30,28,31,96,31,45,31,83,31,83,30,241,31,241,30,106,31,106,30,197,31,115,31,209,31,209,30,209,29,67,31,240,31,65,31,160,31,61,31,183,31,136,31,136,30,83,31,15,31,66,31,51,31,51,30,6,31,108,31,31,31,90,31,88,31,83,31,45,31,45,30,45,29,45,28,45,27,227,31,227,30,12,31,69,31,151,31,57,31,65,31,187,31,187,30,9,31,72,31,172,31,48,31,48,30,195,31,150,31,52,31,245,31,37,31,19,31,156,31,241,31,204,31,107,31,95,31,27,31,80,31,80,30,36,31,191,31,160,31,224,31,37,31,235,31,112,31,104,31,107,31,39,31,86,31,86,30,204,31,121,31,124,31,52,31,189,31,104,31,104,30,25,31,78,31,170,31,170,30,170,29,113,31,170,31,170,30,124,31,167,31,210,31,195,31,247,31,95,31,14,31,231,31,120,31,141,31,61,31,2,31,237,31,154,31,89,31,89,30,8,31,243,31,4,31,4,30,23,31,19,31,19,30,19,29,192,31,29,31,228,31,234,31,25,31,209,31,35,31,56,31,7,31,160,31,126,31,186,31,47,31,93,31,93,31,255,31,187,31,210,31,21,31,119,31,5,31,129,31,129,30,98,31,16,31,215,31,177,31,157,31,157,30,157,29,59,31,59,30,21,31,90,31,164,31,61,31,231,31,120,31,229,31,233,31,54,31,116,31,116,30,208,31,6,31,250,31,94,31,22,31,190,31,190,30,92,31,92,30,17,31,176,31,146,31,240,31,53,31,37,31,110,31,205,31,222,31,242,31,173,31,15,31,168,31,137,31,137,30,227,31,34,31,107,31,230,31,230,30,85,31,85,30,91,31,78,31,136,31,207,31,69,31,116,31,28,31,107,31,107,30,191,31,78,31,62,31,108,31,47,31,120,31,101,31,42,31,205,31,111,31,111,30,111,29,177,31,79,31,79,30,38,31,215,31,215,30,205,31,22,31,22,30,89,31,209,31,153,31,153,30,142,31,97,31,220,31,205,31,167,31,247,31,43,31,78,31,32,31,154,31,46,31,191,31,191,30,191,29,228,31,228,30,228,29,54,31,119,31,141,31,103,31,193,31,193,30,199,31,120,31,250,31,7,31,7,30,80,31,49,31,24,31,24,30,36,31,61,31,61,30,53,31,180,31,180,30,202,31,85,31,172,31,63,31,117,31,8,31,122,31,182,31,118,31,118,30,171,31,171,30,192,31,253,31,147,31,147,31,70,31,99,31,36,31,6,31,228,31,97,31,215,31,215,30,43,31,94,31,148,31,134,31,152,31,225,31,8,31,10,31,110,31,65,31,151,31,145,31,77,31,251,31,83,31,218,31,92,31,62,31,206,31,62,31,255,31,127,31,124,31,124,30,225,31,17,31,196,31,166,31,88,31,201,31,251,31,39,31,222,31,205,31,142,31,142,30,80,31,74,31,55,31,92,31,34,31,31,31,165,31,165,30,133,31,133,30,100,31,68,31,11,31,11,30,80,31,80,30,88,31,207,31,134,31,204,31,61,31,92,31,98,31,163,31,252,31,36,31,36,30,36,29,42,31,124,31,124,30,196,31,50,31,29,31,195,31,245,31,228,31,228,30,216,31,10,31,186,31,186,30,111,31,49,31,37,31,200,31,242,31,58,31,58,30,58,29,58,28,6,31,151,31,151,30,141,31,141,31,45,31,33,31,200,31,143,31,143,30,49,31,166,31,170,31,237,31,211,31,184,31,7,31,7,30,255,31,114,31,155,31,90,31,151,31,131,31,131,31,151,31,151,30,96,31,159,31,248,31,219,31,219,30,129,31,168,31,220,31,138,31,166,31,187,31,108,31,51,31,176,31,22,31,180,31,75,31,82,31,82,30,221,31,251,31,181,31,26,31,104,31,104,30,104,29,216,31,103,31,234,31,82,31,159,31,31,31,133,31,50,31,230,31,91,31,46,31,38,31,65,31,65,30,207,31,207,30,106,31,106,30,120,31,120,30,88,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
