-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_775 is
end project_tb_775;

architecture project_tb_arch_775 of project_tb_775 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 199;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,180,0,131,0,86,0,105,0,0,0,154,0,0,0,235,0,95,0,168,0,164,0,90,0,0,0,43,0,167,0,0,0,152,0,219,0,157,0,121,0,234,0,132,0,0,0,0,0,0,0,235,0,16,0,160,0,110,0,0,0,62,0,210,0,35,0,34,0,0,0,0,0,0,0,145,0,142,0,135,0,0,0,45,0,90,0,29,0,106,0,0,0,33,0,0,0,0,0,110,0,0,0,133,0,0,0,202,0,193,0,150,0,0,0,45,0,0,0,0,0,0,0,93,0,133,0,176,0,90,0,108,0,19,0,176,0,106,0,0,0,235,0,12,0,152,0,82,0,25,0,0,0,158,0,126,0,122,0,215,0,231,0,167,0,0,0,84,0,51,0,225,0,221,0,239,0,102,0,0,0,142,0,55,0,213,0,120,0,105,0,230,0,0,0,0,0,182,0,0,0,169,0,119,0,42,0,0,0,19,0,91,0,47,0,242,0,57,0,215,0,0,0,9,0,0,0,118,0,192,0,173,0,13,0,5,0,126,0,172,0,138,0,106,0,0,0,0,0,96,0,115,0,20,0,0,0,56,0,153,0,120,0,0,0,193,0,82,0,151,0,196,0,194,0,21,0,76,0,26,0,252,0,200,0,241,0,213,0,0,0,0,0,0,0,0,0,0,0,196,0,91,0,140,0,21,0,162,0,0,0,33,0,0,0,88,0,90,0,0,0,110,0,48,0,103,0,6,0,238,0,101,0,172,0,59,0,0,0,112,0,0,0,96,0,118,0,94,0,0,0,136,0,155,0,9,0,146,0,246,0,177,0,253,0,0,0,176,0,253,0,240,0,245,0,220,0,148,0,32,0,139,0,185,0,161,0,2,0,228,0,98,0,176,0,226,0);
signal scenario_full  : scenario_type := (0,0,180,31,131,31,86,31,105,31,105,30,154,31,154,30,235,31,95,31,168,31,164,31,90,31,90,30,43,31,167,31,167,30,152,31,219,31,157,31,121,31,234,31,132,31,132,30,132,29,132,28,235,31,16,31,160,31,110,31,110,30,62,31,210,31,35,31,34,31,34,30,34,29,34,28,145,31,142,31,135,31,135,30,45,31,90,31,29,31,106,31,106,30,33,31,33,30,33,29,110,31,110,30,133,31,133,30,202,31,193,31,150,31,150,30,45,31,45,30,45,29,45,28,93,31,133,31,176,31,90,31,108,31,19,31,176,31,106,31,106,30,235,31,12,31,152,31,82,31,25,31,25,30,158,31,126,31,122,31,215,31,231,31,167,31,167,30,84,31,51,31,225,31,221,31,239,31,102,31,102,30,142,31,55,31,213,31,120,31,105,31,230,31,230,30,230,29,182,31,182,30,169,31,119,31,42,31,42,30,19,31,91,31,47,31,242,31,57,31,215,31,215,30,9,31,9,30,118,31,192,31,173,31,13,31,5,31,126,31,172,31,138,31,106,31,106,30,106,29,96,31,115,31,20,31,20,30,56,31,153,31,120,31,120,30,193,31,82,31,151,31,196,31,194,31,21,31,76,31,26,31,252,31,200,31,241,31,213,31,213,30,213,29,213,28,213,27,213,26,196,31,91,31,140,31,21,31,162,31,162,30,33,31,33,30,88,31,90,31,90,30,110,31,48,31,103,31,6,31,238,31,101,31,172,31,59,31,59,30,112,31,112,30,96,31,118,31,94,31,94,30,136,31,155,31,9,31,146,31,246,31,177,31,253,31,253,30,176,31,253,31,240,31,245,31,220,31,148,31,32,31,139,31,185,31,161,31,2,31,228,31,98,31,176,31,226,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
