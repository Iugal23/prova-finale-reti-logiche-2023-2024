-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 678;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (67,0,218,0,0,0,252,0,253,0,167,0,0,0,0,0,28,0,16,0,114,0,173,0,0,0,17,0,0,0,58,0,194,0,207,0,171,0,22,0,138,0,230,0,198,0,30,0,0,0,13,0,0,0,14,0,67,0,0,0,60,0,0,0,87,0,0,0,205,0,0,0,0,0,221,0,0,0,17,0,152,0,252,0,244,0,133,0,17,0,92,0,170,0,109,0,185,0,0,0,67,0,227,0,239,0,0,0,50,0,0,0,158,0,251,0,0,0,34,0,91,0,0,0,164,0,72,0,140,0,235,0,213,0,0,0,79,0,132,0,196,0,199,0,239,0,186,0,109,0,190,0,69,0,146,0,46,0,250,0,156,0,129,0,113,0,203,0,0,0,201,0,0,0,0,0,246,0,241,0,0,0,37,0,60,0,70,0,70,0,60,0,0,0,0,0,0,0,164,0,103,0,247,0,163,0,209,0,25,0,3,0,217,0,36,0,87,0,185,0,0,0,145,0,68,0,79,0,132,0,234,0,0,0,32,0,55,0,93,0,0,0,91,0,113,0,249,0,87,0,0,0,170,0,0,0,243,0,20,0,92,0,197,0,125,0,229,0,160,0,115,0,84,0,0,0,65,0,80,0,234,0,74,0,0,0,0,0,105,0,0,0,0,0,87,0,180,0,138,0,18,0,106,0,0,0,13,0,22,0,110,0,108,0,214,0,61,0,134,0,0,0,66,0,161,0,91,0,0,0,126,0,102,0,163,0,149,0,62,0,0,0,0,0,122,0,0,0,0,0,20,0,99,0,46,0,17,0,13,0,0,0,100,0,114,0,237,0,0,0,48,0,59,0,136,0,198,0,0,0,0,0,196,0,126,0,0,0,197,0,89,0,164,0,113,0,253,0,230,0,104,0,255,0,149,0,196,0,156,0,86,0,123,0,22,0,233,0,48,0,24,0,181,0,24,0,90,0,197,0,215,0,0,0,102,0,66,0,248,0,193,0,129,0,58,0,79,0,82,0,193,0,150,0,246,0,83,0,140,0,0,0,211,0,55,0,46,0,230,0,196,0,0,0,109,0,221,0,0,0,0,0,0,0,15,0,140,0,230,0,111,0,240,0,133,0,26,0,191,0,4,0,122,0,152,0,205,0,76,0,162,0,239,0,193,0,198,0,207,0,250,0,0,0,0,0,46,0,248,0,43,0,241,0,34,0,164,0,0,0,11,0,32,0,129,0,30,0,168,0,1,0,71,0,3,0,0,0,16,0,103,0,167,0,126,0,208,0,56,0,0,0,61,0,0,0,49,0,41,0,106,0,197,0,64,0,245,0,192,0,107,0,118,0,0,0,105,0,0,0,155,0,0,0,0,0,202,0,130,0,176,0,180,0,0,0,137,0,24,0,2,0,142,0,138,0,225,0,168,0,0,0,162,0,14,0,219,0,0,0,26,0,150,0,208,0,0,0,0,0,150,0,158,0,0,0,26,0,0,0,0,0,91,0,60,0,129,0,0,0,0,0,57,0,122,0,155,0,227,0,170,0,7,0,100,0,238,0,231,0,56,0,61,0,249,0,0,0,217,0,175,0,97,0,0,0,238,0,236,0,17,0,168,0,61,0,45,0,255,0,23,0,86,0,30,0,115,0,0,0,96,0,40,0,211,0,0,0,16,0,58,0,16,0,191,0,33,0,0,0,202,0,169,0,62,0,180,0,233,0,233,0,60,0,208,0,106,0,68,0,0,0,198,0,193,0,53,0,86,0,228,0,0,0,221,0,0,0,12,0,0,0,200,0,209,0,196,0,104,0,252,0,0,0,0,0,214,0,246,0,242,0,231,0,28,0,81,0,239,0,118,0,74,0,110,0,125,0,219,0,0,0,0,0,147,0,0,0,0,0,237,0,0,0,5,0,146,0,138,0,14,0,122,0,29,0,235,0,138,0,71,0,175,0,67,0,170,0,245,0,0,0,198,0,138,0,243,0,0,0,92,0,109,0,134,0,0,0,227,0,48,0,190,0,51,0,0,0,111,0,6,0,189,0,61,0,0,0,141,0,227,0,130,0,179,0,8,0,97,0,139,0,0,0,0,0,213,0,95,0,177,0,177,0,84,0,0,0,0,0,0,0,135,0,25,0,251,0,211,0,156,0,62,0,173,0,217,0,83,0,56,0,71,0,74,0,0,0,148,0,99,0,218,0,29,0,225,0,244,0,243,0,123,0,27,0,134,0,84,0,233,0,49,0,179,0,228,0,0,0,214,0,160,0,5,0,0,0,6,0,0,0,0,0,0,0,0,0,23,0,234,0,72,0,248,0,0,0,0,0,0,0,141,0,216,0,81,0,169,0,248,0,7,0,169,0,34,0,188,0,0,0,147,0,181,0,236,0,31,0,32,0,0,0,19,0,80,0,0,0,22,0,152,0,230,0,29,0,192,0,123,0,224,0,163,0,43,0,6,0,233,0,0,0,205,0,16,0,0,0,166,0,0,0,110,0,82,0,155,0,226,0,224,0,111,0,75,0,242,0,165,0,70,0,44,0,0,0,100,0,175,0,83,0,5,0,0,0,72,0,123,0,203,0,134,0,230,0,44,0,77,0,0,0,0,0,206,0,23,0,93,0,0,0,41,0,47,0,92,0,47,0,152,0,202,0,0,0,98,0,0,0,0,0,215,0,51,0,0,0,56,0,0,0,137,0,60,0,247,0,210,0,0,0,59,0,29,0,178,0,209,0,83,0,38,0,0,0,66,0,120,0,15,0,0,0,67,0,0,0,0,0,0,0,220,0,30,0,105,0,152,0,188,0,108,0,30,0,0,0,0,0,144,0,77,0,0,0,167,0,0,0,237,0,62,0,11,0,246,0,156,0,90,0,3,0,0,0,150,0,0,0,88,0,0,0,172,0,67,0,214,0,249,0,0,0,0,0,7,0,165,0,221,0,22,0,188,0,54,0,0,0,40,0,131,0,202,0,168,0,112,0,0,0,168,0,0,0,254,0,115,0,168,0,192,0,26,0,152,0,214,0,223,0,16,0,62,0,0,0,160,0,211,0,73,0);
signal scenario_full  : scenario_type := (67,31,218,31,218,30,252,31,253,31,167,31,167,30,167,29,28,31,16,31,114,31,173,31,173,30,17,31,17,30,58,31,194,31,207,31,171,31,22,31,138,31,230,31,198,31,30,31,30,30,13,31,13,30,14,31,67,31,67,30,60,31,60,30,87,31,87,30,205,31,205,30,205,29,221,31,221,30,17,31,152,31,252,31,244,31,133,31,17,31,92,31,170,31,109,31,185,31,185,30,67,31,227,31,239,31,239,30,50,31,50,30,158,31,251,31,251,30,34,31,91,31,91,30,164,31,72,31,140,31,235,31,213,31,213,30,79,31,132,31,196,31,199,31,239,31,186,31,109,31,190,31,69,31,146,31,46,31,250,31,156,31,129,31,113,31,203,31,203,30,201,31,201,30,201,29,246,31,241,31,241,30,37,31,60,31,70,31,70,31,60,31,60,30,60,29,60,28,164,31,103,31,247,31,163,31,209,31,25,31,3,31,217,31,36,31,87,31,185,31,185,30,145,31,68,31,79,31,132,31,234,31,234,30,32,31,55,31,93,31,93,30,91,31,113,31,249,31,87,31,87,30,170,31,170,30,243,31,20,31,92,31,197,31,125,31,229,31,160,31,115,31,84,31,84,30,65,31,80,31,234,31,74,31,74,30,74,29,105,31,105,30,105,29,87,31,180,31,138,31,18,31,106,31,106,30,13,31,22,31,110,31,108,31,214,31,61,31,134,31,134,30,66,31,161,31,91,31,91,30,126,31,102,31,163,31,149,31,62,31,62,30,62,29,122,31,122,30,122,29,20,31,99,31,46,31,17,31,13,31,13,30,100,31,114,31,237,31,237,30,48,31,59,31,136,31,198,31,198,30,198,29,196,31,126,31,126,30,197,31,89,31,164,31,113,31,253,31,230,31,104,31,255,31,149,31,196,31,156,31,86,31,123,31,22,31,233,31,48,31,24,31,181,31,24,31,90,31,197,31,215,31,215,30,102,31,66,31,248,31,193,31,129,31,58,31,79,31,82,31,193,31,150,31,246,31,83,31,140,31,140,30,211,31,55,31,46,31,230,31,196,31,196,30,109,31,221,31,221,30,221,29,221,28,15,31,140,31,230,31,111,31,240,31,133,31,26,31,191,31,4,31,122,31,152,31,205,31,76,31,162,31,239,31,193,31,198,31,207,31,250,31,250,30,250,29,46,31,248,31,43,31,241,31,34,31,164,31,164,30,11,31,32,31,129,31,30,31,168,31,1,31,71,31,3,31,3,30,16,31,103,31,167,31,126,31,208,31,56,31,56,30,61,31,61,30,49,31,41,31,106,31,197,31,64,31,245,31,192,31,107,31,118,31,118,30,105,31,105,30,155,31,155,30,155,29,202,31,130,31,176,31,180,31,180,30,137,31,24,31,2,31,142,31,138,31,225,31,168,31,168,30,162,31,14,31,219,31,219,30,26,31,150,31,208,31,208,30,208,29,150,31,158,31,158,30,26,31,26,30,26,29,91,31,60,31,129,31,129,30,129,29,57,31,122,31,155,31,227,31,170,31,7,31,100,31,238,31,231,31,56,31,61,31,249,31,249,30,217,31,175,31,97,31,97,30,238,31,236,31,17,31,168,31,61,31,45,31,255,31,23,31,86,31,30,31,115,31,115,30,96,31,40,31,211,31,211,30,16,31,58,31,16,31,191,31,33,31,33,30,202,31,169,31,62,31,180,31,233,31,233,31,60,31,208,31,106,31,68,31,68,30,198,31,193,31,53,31,86,31,228,31,228,30,221,31,221,30,12,31,12,30,200,31,209,31,196,31,104,31,252,31,252,30,252,29,214,31,246,31,242,31,231,31,28,31,81,31,239,31,118,31,74,31,110,31,125,31,219,31,219,30,219,29,147,31,147,30,147,29,237,31,237,30,5,31,146,31,138,31,14,31,122,31,29,31,235,31,138,31,71,31,175,31,67,31,170,31,245,31,245,30,198,31,138,31,243,31,243,30,92,31,109,31,134,31,134,30,227,31,48,31,190,31,51,31,51,30,111,31,6,31,189,31,61,31,61,30,141,31,227,31,130,31,179,31,8,31,97,31,139,31,139,30,139,29,213,31,95,31,177,31,177,31,84,31,84,30,84,29,84,28,135,31,25,31,251,31,211,31,156,31,62,31,173,31,217,31,83,31,56,31,71,31,74,31,74,30,148,31,99,31,218,31,29,31,225,31,244,31,243,31,123,31,27,31,134,31,84,31,233,31,49,31,179,31,228,31,228,30,214,31,160,31,5,31,5,30,6,31,6,30,6,29,6,28,6,27,23,31,234,31,72,31,248,31,248,30,248,29,248,28,141,31,216,31,81,31,169,31,248,31,7,31,169,31,34,31,188,31,188,30,147,31,181,31,236,31,31,31,32,31,32,30,19,31,80,31,80,30,22,31,152,31,230,31,29,31,192,31,123,31,224,31,163,31,43,31,6,31,233,31,233,30,205,31,16,31,16,30,166,31,166,30,110,31,82,31,155,31,226,31,224,31,111,31,75,31,242,31,165,31,70,31,44,31,44,30,100,31,175,31,83,31,5,31,5,30,72,31,123,31,203,31,134,31,230,31,44,31,77,31,77,30,77,29,206,31,23,31,93,31,93,30,41,31,47,31,92,31,47,31,152,31,202,31,202,30,98,31,98,30,98,29,215,31,51,31,51,30,56,31,56,30,137,31,60,31,247,31,210,31,210,30,59,31,29,31,178,31,209,31,83,31,38,31,38,30,66,31,120,31,15,31,15,30,67,31,67,30,67,29,67,28,220,31,30,31,105,31,152,31,188,31,108,31,30,31,30,30,30,29,144,31,77,31,77,30,167,31,167,30,237,31,62,31,11,31,246,31,156,31,90,31,3,31,3,30,150,31,150,30,88,31,88,30,172,31,67,31,214,31,249,31,249,30,249,29,7,31,165,31,221,31,22,31,188,31,54,31,54,30,40,31,131,31,202,31,168,31,112,31,112,30,168,31,168,30,254,31,115,31,168,31,192,31,26,31,152,31,214,31,223,31,16,31,62,31,62,30,160,31,211,31,73,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
