-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 683;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (147,0,186,0,234,0,197,0,241,0,163,0,33,0,182,0,61,0,74,0,254,0,237,0,10,0,34,0,0,0,68,0,242,0,141,0,3,0,225,0,124,0,180,0,221,0,0,0,227,0,30,0,0,0,109,0,231,0,148,0,81,0,120,0,31,0,227,0,74,0,194,0,43,0,0,0,176,0,130,0,30,0,234,0,241,0,94,0,169,0,95,0,219,0,206,0,49,0,0,0,0,0,94,0,129,0,129,0,0,0,142,0,58,0,0,0,2,0,0,0,113,0,30,0,191,0,0,0,57,0,213,0,131,0,74,0,120,0,0,0,22,0,0,0,158,0,176,0,0,0,0,0,181,0,247,0,0,0,0,0,0,0,0,0,108,0,179,0,0,0,40,0,19,0,67,0,70,0,141,0,235,0,87,0,124,0,109,0,160,0,134,0,67,0,206,0,246,0,247,0,227,0,246,0,237,0,217,0,62,0,0,0,240,0,101,0,98,0,152,0,120,0,245,0,155,0,203,0,254,0,206,0,112,0,0,0,232,0,159,0,193,0,60,0,127,0,9,0,31,0,232,0,55,0,0,0,37,0,0,0,105,0,0,0,129,0,76,0,0,0,0,0,195,0,32,0,0,0,121,0,217,0,46,0,178,0,170,0,6,0,23,0,233,0,248,0,160,0,247,0,199,0,0,0,66,0,94,0,0,0,0,0,40,0,61,0,0,0,121,0,38,0,0,0,39,0,0,0,125,0,71,0,65,0,101,0,87,0,217,0,26,0,183,0,0,0,0,0,228,0,138,0,0,0,250,0,126,0,161,0,158,0,246,0,64,0,138,0,201,0,0,0,126,0,0,0,148,0,74,0,83,0,223,0,0,0,0,0,0,0,167,0,0,0,0,0,207,0,172,0,1,0,132,0,164,0,180,0,0,0,205,0,210,0,20,0,123,0,56,0,243,0,198,0,22,0,52,0,105,0,238,0,250,0,0,0,47,0,0,0,57,0,195,0,27,0,120,0,0,0,180,0,17,0,18,0,84,0,0,0,0,0,0,0,0,0,40,0,1,0,227,0,108,0,98,0,128,0,116,0,50,0,17,0,162,0,0,0,241,0,70,0,76,0,0,0,162,0,9,0,22,0,182,0,0,0,188,0,192,0,0,0,152,0,92,0,197,0,0,0,21,0,102,0,208,0,0,0,249,0,141,0,122,0,109,0,0,0,0,0,77,0,22,0,0,0,0,0,53,0,0,0,0,0,55,0,52,0,231,0,83,0,0,0,0,0,0,0,174,0,133,0,125,0,211,0,77,0,170,0,38,0,167,0,0,0,0,0,137,0,144,0,205,0,94,0,235,0,169,0,0,0,26,0,0,0,0,0,0,0,0,0,119,0,37,0,0,0,0,0,131,0,51,0,0,0,17,0,0,0,61,0,0,0,156,0,179,0,227,0,155,0,0,0,150,0,240,0,218,0,238,0,215,0,172,0,143,0,63,0,0,0,198,0,220,0,241,0,38,0,177,0,236,0,117,0,146,0,211,0,0,0,0,0,184,0,148,0,0,0,0,0,241,0,77,0,0,0,114,0,111,0,39,0,0,0,182,0,124,0,247,0,214,0,85,0,0,0,117,0,0,0,0,0,0,0,171,0,47,0,188,0,97,0,233,0,125,0,3,0,60,0,0,0,213,0,101,0,10,0,105,0,171,0,0,0,107,0,247,0,0,0,175,0,0,0,0,0,62,0,134,0,78,0,222,0,200,0,107,0,204,0,135,0,248,0,217,0,219,0,5,0,0,0,135,0,0,0,0,0,116,0,0,0,0,0,78,0,192,0,147,0,38,0,189,0,0,0,28,0,0,0,0,0,174,0,100,0,174,0,36,0,63,0,101,0,22,0,0,0,207,0,211,0,0,0,0,0,111,0,47,0,69,0,0,0,245,0,98,0,53,0,55,0,192,0,87,0,64,0,105,0,41,0,253,0,57,0,81,0,85,0,0,0,0,0,226,0,208,0,68,0,27,0,20,0,253,0,184,0,221,0,63,0,78,0,140,0,240,0,141,0,229,0,0,0,209,0,164,0,131,0,116,0,0,0,84,0,93,0,152,0,34,0,61,0,255,0,63,0,35,0,26,0,140,0,152,0,60,0,26,0,255,0,105,0,254,0,211,0,10,0,169,0,30,0,105,0,82,0,178,0,202,0,80,0,0,0,0,0,250,0,72,0,192,0,69,0,242,0,163,0,0,0,79,0,0,0,169,0,49,0,143,0,0,0,0,0,0,0,35,0,0,0,158,0,153,0,0,0,93,0,60,0,200,0,86,0,167,0,100,0,43,0,109,0,83,0,184,0,0,0,0,0,220,0,159,0,27,0,105,0,88,0,189,0,94,0,14,0,153,0,19,0,0,0,6,0,0,0,0,0,162,0,201,0,137,0,0,0,83,0,72,0,191,0,50,0,229,0,251,0,206,0,160,0,81,0,132,0,209,0,0,0,218,0,0,0,185,0,5,0,144,0,0,0,121,0,172,0,51,0,9,0,27,0,211,0,128,0,28,0,141,0,220,0,0,0,0,0,158,0,188,0,8,0,10,0,225,0,7,0,125,0,93,0,81,0,86,0,250,0,243,0,34,0,11,0,59,0,0,0,0,0,68,0,175,0,160,0,236,0,0,0,213,0,179,0,106,0,180,0,93,0,52,0,39,0,130,0,17,0,0,0,104,0,0,0,250,0,79,0,213,0,0,0,228,0,0,0,56,0,80,0,51,0,0,0,121,0,0,0,251,0,214,0,42,0,0,0,166,0,108,0,224,0,113,0,0,0,157,0,0,0,0,0,0,0,54,0,235,0,0,0,45,0,201,0,221,0,116,0,0,0,107,0,128,0,26,0,238,0,0,0,88,0,117,0,250,0,249,0,96,0,0,0,213,0,202,0,0,0,130,0,143,0,0,0,191,0,45,0,38,0,164,0,59,0,104,0,150,0,215,0,28,0,31,0,100,0,200,0,83,0,0,0,59,0,209,0,66,0,238,0,141,0,52,0,0,0,0,0,186,0,198,0,204,0,237,0,0,0,0,0,197,0);
signal scenario_full  : scenario_type := (147,31,186,31,234,31,197,31,241,31,163,31,33,31,182,31,61,31,74,31,254,31,237,31,10,31,34,31,34,30,68,31,242,31,141,31,3,31,225,31,124,31,180,31,221,31,221,30,227,31,30,31,30,30,109,31,231,31,148,31,81,31,120,31,31,31,227,31,74,31,194,31,43,31,43,30,176,31,130,31,30,31,234,31,241,31,94,31,169,31,95,31,219,31,206,31,49,31,49,30,49,29,94,31,129,31,129,31,129,30,142,31,58,31,58,30,2,31,2,30,113,31,30,31,191,31,191,30,57,31,213,31,131,31,74,31,120,31,120,30,22,31,22,30,158,31,176,31,176,30,176,29,181,31,247,31,247,30,247,29,247,28,247,27,108,31,179,31,179,30,40,31,19,31,67,31,70,31,141,31,235,31,87,31,124,31,109,31,160,31,134,31,67,31,206,31,246,31,247,31,227,31,246,31,237,31,217,31,62,31,62,30,240,31,101,31,98,31,152,31,120,31,245,31,155,31,203,31,254,31,206,31,112,31,112,30,232,31,159,31,193,31,60,31,127,31,9,31,31,31,232,31,55,31,55,30,37,31,37,30,105,31,105,30,129,31,76,31,76,30,76,29,195,31,32,31,32,30,121,31,217,31,46,31,178,31,170,31,6,31,23,31,233,31,248,31,160,31,247,31,199,31,199,30,66,31,94,31,94,30,94,29,40,31,61,31,61,30,121,31,38,31,38,30,39,31,39,30,125,31,71,31,65,31,101,31,87,31,217,31,26,31,183,31,183,30,183,29,228,31,138,31,138,30,250,31,126,31,161,31,158,31,246,31,64,31,138,31,201,31,201,30,126,31,126,30,148,31,74,31,83,31,223,31,223,30,223,29,223,28,167,31,167,30,167,29,207,31,172,31,1,31,132,31,164,31,180,31,180,30,205,31,210,31,20,31,123,31,56,31,243,31,198,31,22,31,52,31,105,31,238,31,250,31,250,30,47,31,47,30,57,31,195,31,27,31,120,31,120,30,180,31,17,31,18,31,84,31,84,30,84,29,84,28,84,27,40,31,1,31,227,31,108,31,98,31,128,31,116,31,50,31,17,31,162,31,162,30,241,31,70,31,76,31,76,30,162,31,9,31,22,31,182,31,182,30,188,31,192,31,192,30,152,31,92,31,197,31,197,30,21,31,102,31,208,31,208,30,249,31,141,31,122,31,109,31,109,30,109,29,77,31,22,31,22,30,22,29,53,31,53,30,53,29,55,31,52,31,231,31,83,31,83,30,83,29,83,28,174,31,133,31,125,31,211,31,77,31,170,31,38,31,167,31,167,30,167,29,137,31,144,31,205,31,94,31,235,31,169,31,169,30,26,31,26,30,26,29,26,28,26,27,119,31,37,31,37,30,37,29,131,31,51,31,51,30,17,31,17,30,61,31,61,30,156,31,179,31,227,31,155,31,155,30,150,31,240,31,218,31,238,31,215,31,172,31,143,31,63,31,63,30,198,31,220,31,241,31,38,31,177,31,236,31,117,31,146,31,211,31,211,30,211,29,184,31,148,31,148,30,148,29,241,31,77,31,77,30,114,31,111,31,39,31,39,30,182,31,124,31,247,31,214,31,85,31,85,30,117,31,117,30,117,29,117,28,171,31,47,31,188,31,97,31,233,31,125,31,3,31,60,31,60,30,213,31,101,31,10,31,105,31,171,31,171,30,107,31,247,31,247,30,175,31,175,30,175,29,62,31,134,31,78,31,222,31,200,31,107,31,204,31,135,31,248,31,217,31,219,31,5,31,5,30,135,31,135,30,135,29,116,31,116,30,116,29,78,31,192,31,147,31,38,31,189,31,189,30,28,31,28,30,28,29,174,31,100,31,174,31,36,31,63,31,101,31,22,31,22,30,207,31,211,31,211,30,211,29,111,31,47,31,69,31,69,30,245,31,98,31,53,31,55,31,192,31,87,31,64,31,105,31,41,31,253,31,57,31,81,31,85,31,85,30,85,29,226,31,208,31,68,31,27,31,20,31,253,31,184,31,221,31,63,31,78,31,140,31,240,31,141,31,229,31,229,30,209,31,164,31,131,31,116,31,116,30,84,31,93,31,152,31,34,31,61,31,255,31,63,31,35,31,26,31,140,31,152,31,60,31,26,31,255,31,105,31,254,31,211,31,10,31,169,31,30,31,105,31,82,31,178,31,202,31,80,31,80,30,80,29,250,31,72,31,192,31,69,31,242,31,163,31,163,30,79,31,79,30,169,31,49,31,143,31,143,30,143,29,143,28,35,31,35,30,158,31,153,31,153,30,93,31,60,31,200,31,86,31,167,31,100,31,43,31,109,31,83,31,184,31,184,30,184,29,220,31,159,31,27,31,105,31,88,31,189,31,94,31,14,31,153,31,19,31,19,30,6,31,6,30,6,29,162,31,201,31,137,31,137,30,83,31,72,31,191,31,50,31,229,31,251,31,206,31,160,31,81,31,132,31,209,31,209,30,218,31,218,30,185,31,5,31,144,31,144,30,121,31,172,31,51,31,9,31,27,31,211,31,128,31,28,31,141,31,220,31,220,30,220,29,158,31,188,31,8,31,10,31,225,31,7,31,125,31,93,31,81,31,86,31,250,31,243,31,34,31,11,31,59,31,59,30,59,29,68,31,175,31,160,31,236,31,236,30,213,31,179,31,106,31,180,31,93,31,52,31,39,31,130,31,17,31,17,30,104,31,104,30,250,31,79,31,213,31,213,30,228,31,228,30,56,31,80,31,51,31,51,30,121,31,121,30,251,31,214,31,42,31,42,30,166,31,108,31,224,31,113,31,113,30,157,31,157,30,157,29,157,28,54,31,235,31,235,30,45,31,201,31,221,31,116,31,116,30,107,31,128,31,26,31,238,31,238,30,88,31,117,31,250,31,249,31,96,31,96,30,213,31,202,31,202,30,130,31,143,31,143,30,191,31,45,31,38,31,164,31,59,31,104,31,150,31,215,31,28,31,31,31,100,31,200,31,83,31,83,30,59,31,209,31,66,31,238,31,141,31,52,31,52,30,52,29,186,31,198,31,204,31,237,31,237,30,237,29,197,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
