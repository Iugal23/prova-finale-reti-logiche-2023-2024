-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 601;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,87,0,117,0,197,0,35,0,252,0,239,0,177,0,59,0,237,0,220,0,37,0,107,0,215,0,0,0,193,0,0,0,128,0,13,0,252,0,1,0,178,0,157,0,0,0,36,0,139,0,201,0,209,0,22,0,118,0,24,0,205,0,187,0,64,0,47,0,139,0,244,0,212,0,216,0,0,0,184,0,206,0,136,0,173,0,66,0,168,0,139,0,0,0,156,0,101,0,191,0,40,0,103,0,12,0,104,0,195,0,0,0,111,0,27,0,29,0,0,0,89,0,240,0,159,0,14,0,127,0,238,0,201,0,0,0,95,0,218,0,41,0,91,0,0,0,243,0,37,0,68,0,32,0,186,0,0,0,116,0,129,0,144,0,0,0,224,0,0,0,181,0,31,0,220,0,38,0,0,0,252,0,194,0,123,0,0,0,0,0,198,0,11,0,253,0,120,0,249,0,197,0,0,0,0,0,165,0,9,0,155,0,0,0,187,0,97,0,0,0,0,0,148,0,0,0,249,0,48,0,145,0,0,0,116,0,139,0,0,0,197,0,0,0,2,0,10,0,0,0,186,0,98,0,57,0,195,0,230,0,222,0,166,0,144,0,32,0,183,0,0,0,0,0,0,0,92,0,235,0,193,0,243,0,255,0,252,0,0,0,7,0,129,0,198,0,57,0,19,0,0,0,0,0,202,0,110,0,222,0,220,0,50,0,0,0,136,0,0,0,34,0,253,0,221,0,0,0,44,0,23,0,137,0,44,0,12,0,16,0,0,0,90,0,204,0,12,0,74,0,0,0,67,0,226,0,244,0,23,0,197,0,215,0,45,0,147,0,94,0,100,0,163,0,238,0,28,0,0,0,0,0,48,0,192,0,242,0,73,0,175,0,176,0,0,0,0,0,0,0,41,0,98,0,84,0,251,0,43,0,181,0,148,0,0,0,134,0,26,0,234,0,183,0,159,0,42,0,0,0,44,0,223,0,221,0,243,0,252,0,203,0,0,0,113,0,0,0,50,0,0,0,228,0,0,0,202,0,0,0,240,0,2,0,196,0,70,0,1,0,0,0,0,0,209,0,0,0,0,0,134,0,247,0,54,0,153,0,41,0,35,0,156,0,51,0,252,0,121,0,1,0,98,0,16,0,210,0,126,0,107,0,0,0,4,0,0,0,144,0,2,0,35,0,185,0,0,0,0,0,0,0,237,0,121,0,205,0,0,0,14,0,0,0,0,0,95,0,101,0,62,0,155,0,138,0,106,0,165,0,181,0,53,0,128,0,84,0,211,0,11,0,199,0,239,0,166,0,23,0,35,0,23,0,38,0,0,0,213,0,49,0,0,0,156,0,6,0,0,0,242,0,98,0,0,0,70,0,224,0,0,0,123,0,15,0,60,0,58,0,252,0,0,0,84,0,23,0,209,0,3,0,71,0,175,0,0,0,104,0,146,0,15,0,175,0,234,0,0,0,134,0,116,0,35,0,14,0,241,0,106,0,160,0,16,0,151,0,22,0,59,0,190,0,115,0,0,0,0,0,105,0,42,0,196,0,183,0,0,0,46,0,108,0,159,0,0,0,167,0,141,0,247,0,186,0,248,0,0,0,0,0,0,0,207,0,78,0,31,0,0,0,36,0,7,0,204,0,0,0,157,0,90,0,137,0,135,0,35,0,255,0,18,0,198,0,114,0,226,0,78,0,180,0,1,0,182,0,228,0,79,0,35,0,242,0,0,0,2,0,0,0,110,0,0,0,76,0,204,0,131,0,0,0,0,0,89,0,219,0,133,0,127,0,112,0,11,0,108,0,246,0,253,0,162,0,155,0,119,0,0,0,214,0,102,0,0,0,222,0,251,0,0,0,0,0,44,0,0,0,0,0,158,0,78,0,40,0,164,0,0,0,45,0,146,0,128,0,110,0,187,0,12,0,236,0,56,0,135,0,15,0,0,0,133,0,0,0,92,0,0,0,0,0,224,0,93,0,149,0,220,0,80,0,37,0,196,0,202,0,0,0,163,0,102,0,25,0,0,0,198,0,150,0,88,0,0,0,154,0,61,0,86,0,184,0,179,0,173,0,110,0,13,0,172,0,27,0,118,0,96,0,0,0,203,0,160,0,0,0,205,0,229,0,254,0,47,0,131,0,0,0,130,0,241,0,79,0,6,0,85,0,152,0,86,0,0,0,255,0,102,0,220,0,29,0,49,0,226,0,216,0,5,0,226,0,223,0,174,0,0,0,0,0,228,0,9,0,154,0,18,0,224,0,78,0,0,0,0,0,25,0,182,0,138,0,0,0,206,0,0,0,233,0,15,0,212,0,193,0,237,0,137,0,69,0,82,0,191,0,0,0,178,0,142,0,152,0,15,0,102,0,0,0,137,0,243,0,250,0,148,0,220,0,144,0,15,0,0,0,229,0,238,0,132,0,0,0,0,0,64,0,225,0,89,0,167,0,133,0,0,0,188,0,0,0,159,0,170,0,121,0,135,0,126,0,37,0,8,0,178,0,144,0,60,0,179,0,186,0,84,0,0,0,44,0,0,0,0,0,84,0,0,0,53,0,103,0,15,0,25,0,0,0,0,0,78,0,238,0,11,0,61,0,0,0,0,0,0,0,0,0,57,0,117,0,244,0,0,0,189,0,63,0,0,0,56,0,253,0,14,0,148,0,0,0,6,0,187,0,248,0,228,0,6,0,74,0,200,0);
signal scenario_full  : scenario_type := (0,0,87,31,117,31,197,31,35,31,252,31,239,31,177,31,59,31,237,31,220,31,37,31,107,31,215,31,215,30,193,31,193,30,128,31,13,31,252,31,1,31,178,31,157,31,157,30,36,31,139,31,201,31,209,31,22,31,118,31,24,31,205,31,187,31,64,31,47,31,139,31,244,31,212,31,216,31,216,30,184,31,206,31,136,31,173,31,66,31,168,31,139,31,139,30,156,31,101,31,191,31,40,31,103,31,12,31,104,31,195,31,195,30,111,31,27,31,29,31,29,30,89,31,240,31,159,31,14,31,127,31,238,31,201,31,201,30,95,31,218,31,41,31,91,31,91,30,243,31,37,31,68,31,32,31,186,31,186,30,116,31,129,31,144,31,144,30,224,31,224,30,181,31,31,31,220,31,38,31,38,30,252,31,194,31,123,31,123,30,123,29,198,31,11,31,253,31,120,31,249,31,197,31,197,30,197,29,165,31,9,31,155,31,155,30,187,31,97,31,97,30,97,29,148,31,148,30,249,31,48,31,145,31,145,30,116,31,139,31,139,30,197,31,197,30,2,31,10,31,10,30,186,31,98,31,57,31,195,31,230,31,222,31,166,31,144,31,32,31,183,31,183,30,183,29,183,28,92,31,235,31,193,31,243,31,255,31,252,31,252,30,7,31,129,31,198,31,57,31,19,31,19,30,19,29,202,31,110,31,222,31,220,31,50,31,50,30,136,31,136,30,34,31,253,31,221,31,221,30,44,31,23,31,137,31,44,31,12,31,16,31,16,30,90,31,204,31,12,31,74,31,74,30,67,31,226,31,244,31,23,31,197,31,215,31,45,31,147,31,94,31,100,31,163,31,238,31,28,31,28,30,28,29,48,31,192,31,242,31,73,31,175,31,176,31,176,30,176,29,176,28,41,31,98,31,84,31,251,31,43,31,181,31,148,31,148,30,134,31,26,31,234,31,183,31,159,31,42,31,42,30,44,31,223,31,221,31,243,31,252,31,203,31,203,30,113,31,113,30,50,31,50,30,228,31,228,30,202,31,202,30,240,31,2,31,196,31,70,31,1,31,1,30,1,29,209,31,209,30,209,29,134,31,247,31,54,31,153,31,41,31,35,31,156,31,51,31,252,31,121,31,1,31,98,31,16,31,210,31,126,31,107,31,107,30,4,31,4,30,144,31,2,31,35,31,185,31,185,30,185,29,185,28,237,31,121,31,205,31,205,30,14,31,14,30,14,29,95,31,101,31,62,31,155,31,138,31,106,31,165,31,181,31,53,31,128,31,84,31,211,31,11,31,199,31,239,31,166,31,23,31,35,31,23,31,38,31,38,30,213,31,49,31,49,30,156,31,6,31,6,30,242,31,98,31,98,30,70,31,224,31,224,30,123,31,15,31,60,31,58,31,252,31,252,30,84,31,23,31,209,31,3,31,71,31,175,31,175,30,104,31,146,31,15,31,175,31,234,31,234,30,134,31,116,31,35,31,14,31,241,31,106,31,160,31,16,31,151,31,22,31,59,31,190,31,115,31,115,30,115,29,105,31,42,31,196,31,183,31,183,30,46,31,108,31,159,31,159,30,167,31,141,31,247,31,186,31,248,31,248,30,248,29,248,28,207,31,78,31,31,31,31,30,36,31,7,31,204,31,204,30,157,31,90,31,137,31,135,31,35,31,255,31,18,31,198,31,114,31,226,31,78,31,180,31,1,31,182,31,228,31,79,31,35,31,242,31,242,30,2,31,2,30,110,31,110,30,76,31,204,31,131,31,131,30,131,29,89,31,219,31,133,31,127,31,112,31,11,31,108,31,246,31,253,31,162,31,155,31,119,31,119,30,214,31,102,31,102,30,222,31,251,31,251,30,251,29,44,31,44,30,44,29,158,31,78,31,40,31,164,31,164,30,45,31,146,31,128,31,110,31,187,31,12,31,236,31,56,31,135,31,15,31,15,30,133,31,133,30,92,31,92,30,92,29,224,31,93,31,149,31,220,31,80,31,37,31,196,31,202,31,202,30,163,31,102,31,25,31,25,30,198,31,150,31,88,31,88,30,154,31,61,31,86,31,184,31,179,31,173,31,110,31,13,31,172,31,27,31,118,31,96,31,96,30,203,31,160,31,160,30,205,31,229,31,254,31,47,31,131,31,131,30,130,31,241,31,79,31,6,31,85,31,152,31,86,31,86,30,255,31,102,31,220,31,29,31,49,31,226,31,216,31,5,31,226,31,223,31,174,31,174,30,174,29,228,31,9,31,154,31,18,31,224,31,78,31,78,30,78,29,25,31,182,31,138,31,138,30,206,31,206,30,233,31,15,31,212,31,193,31,237,31,137,31,69,31,82,31,191,31,191,30,178,31,142,31,152,31,15,31,102,31,102,30,137,31,243,31,250,31,148,31,220,31,144,31,15,31,15,30,229,31,238,31,132,31,132,30,132,29,64,31,225,31,89,31,167,31,133,31,133,30,188,31,188,30,159,31,170,31,121,31,135,31,126,31,37,31,8,31,178,31,144,31,60,31,179,31,186,31,84,31,84,30,44,31,44,30,44,29,84,31,84,30,53,31,103,31,15,31,25,31,25,30,25,29,78,31,238,31,11,31,61,31,61,30,61,29,61,28,61,27,57,31,117,31,244,31,244,30,189,31,63,31,63,30,56,31,253,31,14,31,148,31,148,30,6,31,187,31,248,31,228,31,6,31,74,31,200,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
