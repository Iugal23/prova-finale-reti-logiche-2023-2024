-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_105 is
end project_tb_105;

architecture project_tb_arch_105 of project_tb_105 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 771;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (62,0,118,0,37,0,43,0,49,0,184,0,125,0,126,0,210,0,108,0,148,0,79,0,110,0,189,0,158,0,237,0,191,0,190,0,50,0,141,0,26,0,83,0,121,0,108,0,116,0,0,0,35,0,255,0,213,0,167,0,0,0,229,0,215,0,0,0,240,0,98,0,0,0,200,0,117,0,217,0,118,0,89,0,147,0,192,0,174,0,221,0,139,0,108,0,98,0,182,0,179,0,134,0,91,0,188,0,0,0,179,0,27,0,164,0,85,0,0,0,174,0,97,0,9,0,83,0,187,0,218,0,11,0,167,0,223,0,0,0,32,0,0,0,0,0,16,0,7,0,0,0,0,0,0,0,206,0,0,0,0,0,201,0,38,0,183,0,43,0,249,0,0,0,94,0,0,0,0,0,0,0,159,0,19,0,113,0,154,0,0,0,173,0,0,0,214,0,89,0,1,0,68,0,65,0,0,0,141,0,205,0,211,0,136,0,180,0,143,0,232,0,138,0,0,0,0,0,65,0,39,0,183,0,39,0,209,0,0,0,246,0,0,0,84,0,224,0,53,0,127,0,121,0,0,0,220,0,0,0,0,0,114,0,186,0,247,0,207,0,254,0,0,0,184,0,109,0,136,0,0,0,0,0,0,0,0,0,62,0,9,0,9,0,0,0,0,0,70,0,57,0,97,0,11,0,211,0,0,0,208,0,91,0,0,0,119,0,203,0,202,0,237,0,253,0,132,0,57,0,94,0,156,0,181,0,91,0,224,0,12,0,245,0,0,0,19,0,9,0,253,0,4,0,195,0,117,0,114,0,102,0,0,0,182,0,0,0,223,0,5,0,115,0,0,0,27,0,194,0,236,0,0,0,0,0,218,0,77,0,168,0,237,0,195,0,60,0,92,0,156,0,0,0,151,0,0,0,129,0,192,0,0,0,0,0,20,0,28,0,0,0,0,0,212,0,188,0,28,0,0,0,34,0,139,0,246,0,71,0,43,0,24,0,0,0,23,0,214,0,143,0,243,0,76,0,252,0,10,0,132,0,209,0,101,0,228,0,176,0,0,0,182,0,175,0,80,0,118,0,104,0,1,0,246,0,0,0,228,0,146,0,16,0,0,0,103,0,36,0,238,0,0,0,227,0,81,0,0,0,21,0,152,0,170,0,0,0,246,0,73,0,178,0,229,0,250,0,91,0,230,0,1,0,193,0,188,0,0,0,0,0,7,0,46,0,116,0,151,0,171,0,115,0,0,0,171,0,255,0,234,0,10,0,17,0,70,0,252,0,247,0,57,0,0,0,0,0,218,0,246,0,239,0,62,0,223,0,144,0,103,0,56,0,250,0,79,0,203,0,238,0,134,0,0,0,181,0,65,0,0,0,248,0,190,0,167,0,246,0,68,0,0,0,0,0,0,0,0,0,0,0,0,0,87,0,105,0,186,0,215,0,191,0,2,0,149,0,65,0,207,0,105,0,252,0,75,0,67,0,0,0,218,0,132,0,86,0,0,0,0,0,42,0,0,0,0,0,199,0,81,0,182,0,64,0,93,0,52,0,38,0,140,0,161,0,31,0,147,0,168,0,0,0,45,0,0,0,0,0,241,0,138,0,247,0,0,0,123,0,46,0,77,0,0,0,0,0,155,0,162,0,245,0,0,0,253,0,142,0,181,0,121,0,0,0,0,0,187,0,98,0,0,0,251,0,114,0,167,0,53,0,62,0,63,0,123,0,0,0,58,0,15,0,0,0,168,0,48,0,0,0,210,0,0,0,0,0,0,0,3,0,73,0,127,0,254,0,211,0,205,0,173,0,222,0,0,0,172,0,211,0,160,0,132,0,139,0,0,0,0,0,99,0,255,0,138,0,5,0,254,0,250,0,158,0,3,0,1,0,98,0,62,0,0,0,201,0,50,0,20,0,2,0,168,0,0,0,99,0,198,0,250,0,181,0,150,0,218,0,22,0,197,0,36,0,50,0,199,0,121,0,235,0,129,0,16,0,242,0,91,0,164,0,133,0,76,0,81,0,204,0,31,0,0,0,120,0,124,0,114,0,89,0,157,0,193,0,118,0,255,0,45,0,235,0,22,0,182,0,115,0,191,0,239,0,210,0,209,0,0,0,207,0,45,0,0,0,57,0,232,0,73,0,144,0,241,0,0,0,0,0,205,0,0,0,46,0,0,0,246,0,243,0,252,0,0,0,145,0,0,0,216,0,228,0,40,0,124,0,253,0,115,0,8,0,121,0,193,0,73,0,254,0,11,0,119,0,59,0,15,0,171,0,28,0,131,0,191,0,96,0,115,0,10,0,0,0,228,0,0,0,0,0,0,0,84,0,128,0,0,0,196,0,78,0,91,0,175,0,206,0,253,0,46,0,23,0,68,0,0,0,228,0,0,0,158,0,104,0,183,0,72,0,222,0,125,0,244,0,62,0,198,0,161,0,30,0,0,0,209,0,17,0,188,0,0,0,35,0,142,0,5,0,245,0,45,0,0,0,0,0,98,0,19,0,161,0,216,0,240,0,65,0,107,0,224,0,176,0,92,0,139,0,96,0,169,0,12,0,109,0,126,0,196,0,81,0,156,0,0,0,186,0,0,0,41,0,26,0,120,0,135,0,116,0,230,0,0,0,30,0,0,0,58,0,202,0,233,0,209,0,50,0,59,0,0,0,40,0,0,0,66,0,184,0,0,0,0,0,191,0,114,0,0,0,0,0,0,0,99,0,0,0,209,0,37,0,0,0,171,0,88,0,228,0,206,0,162,0,224,0,241,0,196,0,0,0,93,0,72,0,150,0,209,0,99,0,104,0,0,0,237,0,33,0,138,0,52,0,69,0,0,0,0,0,0,0,230,0,246,0,90,0,142,0,207,0,249,0,84,0,28,0,0,0,0,0,91,0,114,0,83,0,124,0,0,0,32,0,88,0,157,0,161,0,0,0,0,0,237,0,182,0,43,0,0,0,85,0,230,0,101,0,136,0,0,0,0,0,67,0,106,0,194,0,65,0,19,0,79,0,219,0,133,0,23,0,123,0,87,0,91,0,0,0,222,0,138,0,0,0,93,0,66,0,66,0,221,0,167,0,73,0,208,0,137,0,0,0,0,0,77,0,20,0,148,0,0,0,47,0,0,0,23,0,225,0,0,0,53,0,240,0,52,0,196,0,71,0,0,0,124,0,238,0,178,0,238,0,28,0,63,0,235,0,116,0,229,0,17,0,0,0,50,0,63,0,235,0,249,0,253,0,219,0,10,0,150,0,222,0,192,0,209,0,116,0,86,0,69,0,118,0,0,0,0,0,117,0,120,0,99,0,111,0,79,0,0,0,25,0,145,0,75,0,81,0,1,0,120,0,112,0,0,0,88,0,0,0,37,0,0,0,124,0,86,0,0,0,81,0,96,0,138,0,3,0,159,0,180,0,5,0,187,0,72,0,0,0,47,0,172,0,235,0,0,0,0,0,70,0);
signal scenario_full  : scenario_type := (62,31,118,31,37,31,43,31,49,31,184,31,125,31,126,31,210,31,108,31,148,31,79,31,110,31,189,31,158,31,237,31,191,31,190,31,50,31,141,31,26,31,83,31,121,31,108,31,116,31,116,30,35,31,255,31,213,31,167,31,167,30,229,31,215,31,215,30,240,31,98,31,98,30,200,31,117,31,217,31,118,31,89,31,147,31,192,31,174,31,221,31,139,31,108,31,98,31,182,31,179,31,134,31,91,31,188,31,188,30,179,31,27,31,164,31,85,31,85,30,174,31,97,31,9,31,83,31,187,31,218,31,11,31,167,31,223,31,223,30,32,31,32,30,32,29,16,31,7,31,7,30,7,29,7,28,206,31,206,30,206,29,201,31,38,31,183,31,43,31,249,31,249,30,94,31,94,30,94,29,94,28,159,31,19,31,113,31,154,31,154,30,173,31,173,30,214,31,89,31,1,31,68,31,65,31,65,30,141,31,205,31,211,31,136,31,180,31,143,31,232,31,138,31,138,30,138,29,65,31,39,31,183,31,39,31,209,31,209,30,246,31,246,30,84,31,224,31,53,31,127,31,121,31,121,30,220,31,220,30,220,29,114,31,186,31,247,31,207,31,254,31,254,30,184,31,109,31,136,31,136,30,136,29,136,28,136,27,62,31,9,31,9,31,9,30,9,29,70,31,57,31,97,31,11,31,211,31,211,30,208,31,91,31,91,30,119,31,203,31,202,31,237,31,253,31,132,31,57,31,94,31,156,31,181,31,91,31,224,31,12,31,245,31,245,30,19,31,9,31,253,31,4,31,195,31,117,31,114,31,102,31,102,30,182,31,182,30,223,31,5,31,115,31,115,30,27,31,194,31,236,31,236,30,236,29,218,31,77,31,168,31,237,31,195,31,60,31,92,31,156,31,156,30,151,31,151,30,129,31,192,31,192,30,192,29,20,31,28,31,28,30,28,29,212,31,188,31,28,31,28,30,34,31,139,31,246,31,71,31,43,31,24,31,24,30,23,31,214,31,143,31,243,31,76,31,252,31,10,31,132,31,209,31,101,31,228,31,176,31,176,30,182,31,175,31,80,31,118,31,104,31,1,31,246,31,246,30,228,31,146,31,16,31,16,30,103,31,36,31,238,31,238,30,227,31,81,31,81,30,21,31,152,31,170,31,170,30,246,31,73,31,178,31,229,31,250,31,91,31,230,31,1,31,193,31,188,31,188,30,188,29,7,31,46,31,116,31,151,31,171,31,115,31,115,30,171,31,255,31,234,31,10,31,17,31,70,31,252,31,247,31,57,31,57,30,57,29,218,31,246,31,239,31,62,31,223,31,144,31,103,31,56,31,250,31,79,31,203,31,238,31,134,31,134,30,181,31,65,31,65,30,248,31,190,31,167,31,246,31,68,31,68,30,68,29,68,28,68,27,68,26,68,25,87,31,105,31,186,31,215,31,191,31,2,31,149,31,65,31,207,31,105,31,252,31,75,31,67,31,67,30,218,31,132,31,86,31,86,30,86,29,42,31,42,30,42,29,199,31,81,31,182,31,64,31,93,31,52,31,38,31,140,31,161,31,31,31,147,31,168,31,168,30,45,31,45,30,45,29,241,31,138,31,247,31,247,30,123,31,46,31,77,31,77,30,77,29,155,31,162,31,245,31,245,30,253,31,142,31,181,31,121,31,121,30,121,29,187,31,98,31,98,30,251,31,114,31,167,31,53,31,62,31,63,31,123,31,123,30,58,31,15,31,15,30,168,31,48,31,48,30,210,31,210,30,210,29,210,28,3,31,73,31,127,31,254,31,211,31,205,31,173,31,222,31,222,30,172,31,211,31,160,31,132,31,139,31,139,30,139,29,99,31,255,31,138,31,5,31,254,31,250,31,158,31,3,31,1,31,98,31,62,31,62,30,201,31,50,31,20,31,2,31,168,31,168,30,99,31,198,31,250,31,181,31,150,31,218,31,22,31,197,31,36,31,50,31,199,31,121,31,235,31,129,31,16,31,242,31,91,31,164,31,133,31,76,31,81,31,204,31,31,31,31,30,120,31,124,31,114,31,89,31,157,31,193,31,118,31,255,31,45,31,235,31,22,31,182,31,115,31,191,31,239,31,210,31,209,31,209,30,207,31,45,31,45,30,57,31,232,31,73,31,144,31,241,31,241,30,241,29,205,31,205,30,46,31,46,30,246,31,243,31,252,31,252,30,145,31,145,30,216,31,228,31,40,31,124,31,253,31,115,31,8,31,121,31,193,31,73,31,254,31,11,31,119,31,59,31,15,31,171,31,28,31,131,31,191,31,96,31,115,31,10,31,10,30,228,31,228,30,228,29,228,28,84,31,128,31,128,30,196,31,78,31,91,31,175,31,206,31,253,31,46,31,23,31,68,31,68,30,228,31,228,30,158,31,104,31,183,31,72,31,222,31,125,31,244,31,62,31,198,31,161,31,30,31,30,30,209,31,17,31,188,31,188,30,35,31,142,31,5,31,245,31,45,31,45,30,45,29,98,31,19,31,161,31,216,31,240,31,65,31,107,31,224,31,176,31,92,31,139,31,96,31,169,31,12,31,109,31,126,31,196,31,81,31,156,31,156,30,186,31,186,30,41,31,26,31,120,31,135,31,116,31,230,31,230,30,30,31,30,30,58,31,202,31,233,31,209,31,50,31,59,31,59,30,40,31,40,30,66,31,184,31,184,30,184,29,191,31,114,31,114,30,114,29,114,28,99,31,99,30,209,31,37,31,37,30,171,31,88,31,228,31,206,31,162,31,224,31,241,31,196,31,196,30,93,31,72,31,150,31,209,31,99,31,104,31,104,30,237,31,33,31,138,31,52,31,69,31,69,30,69,29,69,28,230,31,246,31,90,31,142,31,207,31,249,31,84,31,28,31,28,30,28,29,91,31,114,31,83,31,124,31,124,30,32,31,88,31,157,31,161,31,161,30,161,29,237,31,182,31,43,31,43,30,85,31,230,31,101,31,136,31,136,30,136,29,67,31,106,31,194,31,65,31,19,31,79,31,219,31,133,31,23,31,123,31,87,31,91,31,91,30,222,31,138,31,138,30,93,31,66,31,66,31,221,31,167,31,73,31,208,31,137,31,137,30,137,29,77,31,20,31,148,31,148,30,47,31,47,30,23,31,225,31,225,30,53,31,240,31,52,31,196,31,71,31,71,30,124,31,238,31,178,31,238,31,28,31,63,31,235,31,116,31,229,31,17,31,17,30,50,31,63,31,235,31,249,31,253,31,219,31,10,31,150,31,222,31,192,31,209,31,116,31,86,31,69,31,118,31,118,30,118,29,117,31,120,31,99,31,111,31,79,31,79,30,25,31,145,31,75,31,81,31,1,31,120,31,112,31,112,30,88,31,88,30,37,31,37,30,124,31,86,31,86,30,81,31,96,31,138,31,3,31,159,31,180,31,5,31,187,31,72,31,72,30,47,31,172,31,235,31,235,30,235,29,70,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
