-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_875 is
end project_tb_875;

architecture project_tb_arch_875 of project_tb_875 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 461;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (98,0,0,0,225,0,251,0,182,0,0,0,129,0,147,0,225,0,158,0,33,0,134,0,0,0,201,0,0,0,0,0,0,0,152,0,0,0,236,0,73,0,0,0,32,0,246,0,0,0,15,0,113,0,0,0,205,0,81,0,132,0,139,0,221,0,96,0,11,0,0,0,13,0,43,0,114,0,243,0,143,0,253,0,237,0,183,0,200,0,42,0,132,0,0,0,0,0,221,0,219,0,125,0,84,0,212,0,235,0,254,0,255,0,0,0,0,0,234,0,223,0,145,0,58,0,225,0,86,0,41,0,48,0,242,0,249,0,65,0,248,0,185,0,97,0,182,0,0,0,67,0,10,0,52,0,124,0,22,0,116,0,190,0,209,0,0,0,11,0,163,0,32,0,0,0,1,0,0,0,221,0,90,0,204,0,0,0,180,0,20,0,23,0,2,0,0,0,110,0,183,0,50,0,123,0,254,0,7,0,146,0,68,0,125,0,80,0,218,0,6,0,0,0,169,0,0,0,0,0,147,0,5,0,0,0,247,0,182,0,179,0,0,0,217,0,76,0,75,0,239,0,0,0,133,0,43,0,242,0,143,0,215,0,234,0,83,0,118,0,26,0,191,0,190,0,0,0,42,0,60,0,53,0,204,0,91,0,146,0,0,0,186,0,204,0,0,0,160,0,97,0,28,0,57,0,0,0,0,0,140,0,87,0,54,0,216,0,151,0,146,0,0,0,102,0,131,0,189,0,192,0,69,0,0,0,69,0,47,0,250,0,77,0,132,0,188,0,6,0,104,0,174,0,25,0,71,0,0,0,34,0,247,0,17,0,229,0,0,0,142,0,227,0,167,0,13,0,140,0,236,0,126,0,116,0,126,0,0,0,0,0,105,0,248,0,57,0,172,0,208,0,206,0,85,0,13,0,121,0,160,0,166,0,188,0,175,0,0,0,110,0,103,0,166,0,0,0,47,0,64,0,33,0,182,0,188,0,0,0,152,0,189,0,105,0,229,0,214,0,41,0,197,0,246,0,0,0,20,0,227,0,29,0,48,0,190,0,127,0,208,0,22,0,98,0,93,0,195,0,40,0,160,0,0,0,62,0,183,0,179,0,132,0,165,0,3,0,85,0,246,0,181,0,178,0,0,0,162,0,73,0,0,0,0,0,245,0,0,0,149,0,219,0,154,0,147,0,0,0,0,0,208,0,125,0,45,0,247,0,59,0,20,0,246,0,0,0,115,0,0,0,0,0,0,0,0,0,5,0,0,0,29,0,138,0,0,0,32,0,0,0,134,0,78,0,232,0,245,0,19,0,254,0,233,0,183,0,170,0,0,0,0,0,66,0,20,0,0,0,207,0,0,0,104,0,227,0,0,0,0,0,233,0,158,0,22,0,240,0,0,0,232,0,0,0,96,0,0,0,0,0,56,0,201,0,158,0,54,0,64,0,253,0,149,0,146,0,39,0,7,0,20,0,0,0,126,0,94,0,214,0,127,0,107,0,205,0,76,0,162,0,60,0,130,0,0,0,22,0,0,0,39,0,0,0,68,0,234,0,81,0,35,0,83,0,224,0,0,0,8,0,229,0,78,0,0,0,127,0,0,0,58,0,133,0,48,0,217,0,171,0,38,0,197,0,19,0,229,0,194,0,122,0,247,0,44,0,188,0,253,0,0,0,97,0,52,0,21,0,46,0,211,0,0,0,0,0,145,0,155,0,48,0,137,0,123,0,0,0,20,0,0,0,106,0,147,0,36,0,0,0,34,0,0,0,32,0,0,0,93,0,57,0,74,0,2,0,236,0,0,0,170,0,58,0,0,0,76,0,142,0,0,0,48,0,247,0,215,0,94,0,59,0,162,0,128,0,132,0,154,0,18,0,4,0,90,0,23,0,153,0,132,0,0,0,0,0,50,0,0,0,25,0,245,0,225,0,95,0,104,0,46,0,100,0,0,0,95,0,114,0,74,0,215,0,17,0,40,0,26,0,164,0,78,0,55,0,3,0,200,0,0,0,244,0,51,0,0,0,9,0,102,0,0,0,18,0,223,0,90,0,125,0,15,0,58,0,20,0,217,0);
signal scenario_full  : scenario_type := (98,31,98,30,225,31,251,31,182,31,182,30,129,31,147,31,225,31,158,31,33,31,134,31,134,30,201,31,201,30,201,29,201,28,152,31,152,30,236,31,73,31,73,30,32,31,246,31,246,30,15,31,113,31,113,30,205,31,81,31,132,31,139,31,221,31,96,31,11,31,11,30,13,31,43,31,114,31,243,31,143,31,253,31,237,31,183,31,200,31,42,31,132,31,132,30,132,29,221,31,219,31,125,31,84,31,212,31,235,31,254,31,255,31,255,30,255,29,234,31,223,31,145,31,58,31,225,31,86,31,41,31,48,31,242,31,249,31,65,31,248,31,185,31,97,31,182,31,182,30,67,31,10,31,52,31,124,31,22,31,116,31,190,31,209,31,209,30,11,31,163,31,32,31,32,30,1,31,1,30,221,31,90,31,204,31,204,30,180,31,20,31,23,31,2,31,2,30,110,31,183,31,50,31,123,31,254,31,7,31,146,31,68,31,125,31,80,31,218,31,6,31,6,30,169,31,169,30,169,29,147,31,5,31,5,30,247,31,182,31,179,31,179,30,217,31,76,31,75,31,239,31,239,30,133,31,43,31,242,31,143,31,215,31,234,31,83,31,118,31,26,31,191,31,190,31,190,30,42,31,60,31,53,31,204,31,91,31,146,31,146,30,186,31,204,31,204,30,160,31,97,31,28,31,57,31,57,30,57,29,140,31,87,31,54,31,216,31,151,31,146,31,146,30,102,31,131,31,189,31,192,31,69,31,69,30,69,31,47,31,250,31,77,31,132,31,188,31,6,31,104,31,174,31,25,31,71,31,71,30,34,31,247,31,17,31,229,31,229,30,142,31,227,31,167,31,13,31,140,31,236,31,126,31,116,31,126,31,126,30,126,29,105,31,248,31,57,31,172,31,208,31,206,31,85,31,13,31,121,31,160,31,166,31,188,31,175,31,175,30,110,31,103,31,166,31,166,30,47,31,64,31,33,31,182,31,188,31,188,30,152,31,189,31,105,31,229,31,214,31,41,31,197,31,246,31,246,30,20,31,227,31,29,31,48,31,190,31,127,31,208,31,22,31,98,31,93,31,195,31,40,31,160,31,160,30,62,31,183,31,179,31,132,31,165,31,3,31,85,31,246,31,181,31,178,31,178,30,162,31,73,31,73,30,73,29,245,31,245,30,149,31,219,31,154,31,147,31,147,30,147,29,208,31,125,31,45,31,247,31,59,31,20,31,246,31,246,30,115,31,115,30,115,29,115,28,115,27,5,31,5,30,29,31,138,31,138,30,32,31,32,30,134,31,78,31,232,31,245,31,19,31,254,31,233,31,183,31,170,31,170,30,170,29,66,31,20,31,20,30,207,31,207,30,104,31,227,31,227,30,227,29,233,31,158,31,22,31,240,31,240,30,232,31,232,30,96,31,96,30,96,29,56,31,201,31,158,31,54,31,64,31,253,31,149,31,146,31,39,31,7,31,20,31,20,30,126,31,94,31,214,31,127,31,107,31,205,31,76,31,162,31,60,31,130,31,130,30,22,31,22,30,39,31,39,30,68,31,234,31,81,31,35,31,83,31,224,31,224,30,8,31,229,31,78,31,78,30,127,31,127,30,58,31,133,31,48,31,217,31,171,31,38,31,197,31,19,31,229,31,194,31,122,31,247,31,44,31,188,31,253,31,253,30,97,31,52,31,21,31,46,31,211,31,211,30,211,29,145,31,155,31,48,31,137,31,123,31,123,30,20,31,20,30,106,31,147,31,36,31,36,30,34,31,34,30,32,31,32,30,93,31,57,31,74,31,2,31,236,31,236,30,170,31,58,31,58,30,76,31,142,31,142,30,48,31,247,31,215,31,94,31,59,31,162,31,128,31,132,31,154,31,18,31,4,31,90,31,23,31,153,31,132,31,132,30,132,29,50,31,50,30,25,31,245,31,225,31,95,31,104,31,46,31,100,31,100,30,95,31,114,31,74,31,215,31,17,31,40,31,26,31,164,31,78,31,55,31,3,31,200,31,200,30,244,31,51,31,51,30,9,31,102,31,102,30,18,31,223,31,90,31,125,31,15,31,58,31,20,31,217,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
