-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 298;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (230,0,38,0,173,0,134,0,133,0,20,0,95,0,0,0,24,0,116,0,155,0,158,0,247,0,0,0,35,0,6,0,142,0,197,0,84,0,0,0,104,0,164,0,40,0,92,0,19,0,199,0,0,0,148,0,128,0,44,0,229,0,246,0,222,0,235,0,101,0,185,0,75,0,148,0,0,0,0,0,240,0,198,0,167,0,167,0,126,0,131,0,183,0,48,0,204,0,115,0,111,0,42,0,135,0,212,0,101,0,178,0,0,0,0,0,63,0,16,0,207,0,157,0,120,0,47,0,165,0,98,0,237,0,200,0,64,0,186,0,0,0,191,0,44,0,26,0,15,0,237,0,16,0,179,0,36,0,26,0,169,0,47,0,0,0,1,0,27,0,139,0,0,0,164,0,130,0,209,0,29,0,12,0,221,0,156,0,0,0,0,0,61,0,239,0,237,0,199,0,252,0,131,0,40,0,176,0,64,0,200,0,69,0,181,0,0,0,202,0,121,0,88,0,0,0,0,0,227,0,92,0,67,0,0,0,0,0,0,0,180,0,146,0,181,0,34,0,0,0,62,0,42,0,217,0,233,0,133,0,17,0,59,0,94,0,247,0,196,0,0,0,62,0,0,0,0,0,69,0,8,0,164,0,28,0,102,0,0,0,121,0,40,0,118,0,247,0,204,0,43,0,99,0,108,0,157,0,0,0,17,0,25,0,44,0,176,0,231,0,104,0,0,0,137,0,0,0,188,0,129,0,53,0,250,0,3,0,179,0,44,0,0,0,72,0,232,0,5,0,29,0,64,0,0,0,188,0,83,0,35,0,8,0,0,0,132,0,148,0,154,0,0,0,4,0,158,0,0,0,146,0,84,0,86,0,217,0,131,0,100,0,77,0,199,0,140,0,0,0,15,0,151,0,181,0,58,0,177,0,119,0,160,0,58,0,0,0,194,0,236,0,157,0,236,0,128,0,181,0,238,0,225,0,173,0,178,0,162,0,63,0,26,0,58,0,198,0,243,0,223,0,46,0,168,0,176,0,0,0,218,0,101,0,0,0,0,0,88,0,32,0,132,0,0,0,49,0,47,0,100,0,241,0,0,0,181,0,110,0,40,0,163,0,0,0,0,0,0,0,140,0,172,0,0,0,0,0,0,0,127,0,255,0,204,0,20,0,0,0,109,0,186,0,33,0,250,0,219,0,78,0,60,0,99,0,50,0,142,0,0,0,0,0,56,0,190,0,206,0,0,0,14,0,231,0,34,0,111,0,47,0,130,0,124,0,226,0,0,0,122,0,0,0,0,0,114,0,0,0,211,0,46,0,46,0,181,0,31,0,197,0,179,0,175,0);
signal scenario_full  : scenario_type := (230,31,38,31,173,31,134,31,133,31,20,31,95,31,95,30,24,31,116,31,155,31,158,31,247,31,247,30,35,31,6,31,142,31,197,31,84,31,84,30,104,31,164,31,40,31,92,31,19,31,199,31,199,30,148,31,128,31,44,31,229,31,246,31,222,31,235,31,101,31,185,31,75,31,148,31,148,30,148,29,240,31,198,31,167,31,167,31,126,31,131,31,183,31,48,31,204,31,115,31,111,31,42,31,135,31,212,31,101,31,178,31,178,30,178,29,63,31,16,31,207,31,157,31,120,31,47,31,165,31,98,31,237,31,200,31,64,31,186,31,186,30,191,31,44,31,26,31,15,31,237,31,16,31,179,31,36,31,26,31,169,31,47,31,47,30,1,31,27,31,139,31,139,30,164,31,130,31,209,31,29,31,12,31,221,31,156,31,156,30,156,29,61,31,239,31,237,31,199,31,252,31,131,31,40,31,176,31,64,31,200,31,69,31,181,31,181,30,202,31,121,31,88,31,88,30,88,29,227,31,92,31,67,31,67,30,67,29,67,28,180,31,146,31,181,31,34,31,34,30,62,31,42,31,217,31,233,31,133,31,17,31,59,31,94,31,247,31,196,31,196,30,62,31,62,30,62,29,69,31,8,31,164,31,28,31,102,31,102,30,121,31,40,31,118,31,247,31,204,31,43,31,99,31,108,31,157,31,157,30,17,31,25,31,44,31,176,31,231,31,104,31,104,30,137,31,137,30,188,31,129,31,53,31,250,31,3,31,179,31,44,31,44,30,72,31,232,31,5,31,29,31,64,31,64,30,188,31,83,31,35,31,8,31,8,30,132,31,148,31,154,31,154,30,4,31,158,31,158,30,146,31,84,31,86,31,217,31,131,31,100,31,77,31,199,31,140,31,140,30,15,31,151,31,181,31,58,31,177,31,119,31,160,31,58,31,58,30,194,31,236,31,157,31,236,31,128,31,181,31,238,31,225,31,173,31,178,31,162,31,63,31,26,31,58,31,198,31,243,31,223,31,46,31,168,31,176,31,176,30,218,31,101,31,101,30,101,29,88,31,32,31,132,31,132,30,49,31,47,31,100,31,241,31,241,30,181,31,110,31,40,31,163,31,163,30,163,29,163,28,140,31,172,31,172,30,172,29,172,28,127,31,255,31,204,31,20,31,20,30,109,31,186,31,33,31,250,31,219,31,78,31,60,31,99,31,50,31,142,31,142,30,142,29,56,31,190,31,206,31,206,30,14,31,231,31,34,31,111,31,47,31,130,31,124,31,226,31,226,30,122,31,122,30,122,29,114,31,114,30,211,31,46,31,46,31,181,31,31,31,197,31,179,31,175,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
