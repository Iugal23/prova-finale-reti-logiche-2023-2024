-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 728;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (209,0,149,0,0,0,0,0,225,0,254,0,178,0,29,0,113,0,0,0,135,0,0,0,248,0,73,0,0,0,84,0,89,0,138,0,60,0,0,0,52,0,0,0,0,0,69,0,0,0,82,0,35,0,195,0,0,0,90,0,167,0,213,0,54,0,16,0,162,0,0,0,0,0,0,0,0,0,219,0,248,0,23,0,243,0,125,0,93,0,87,0,159,0,1,0,138,0,0,0,143,0,0,0,102,0,101,0,0,0,0,0,0,0,10,0,230,0,69,0,101,0,44,0,25,0,115,0,233,0,155,0,0,0,85,0,0,0,200,0,0,0,1,0,0,0,169,0,111,0,0,0,157,0,0,0,232,0,116,0,249,0,0,0,49,0,172,0,20,0,244,0,201,0,227,0,166,0,0,0,137,0,0,0,99,0,210,0,143,0,194,0,229,0,0,0,153,0,0,0,0,0,225,0,0,0,100,0,21,0,0,0,128,0,108,0,9,0,138,0,237,0,0,0,0,0,0,0,136,0,0,0,249,0,9,0,236,0,203,0,28,0,34,0,111,0,0,0,62,0,13,0,6,0,69,0,123,0,91,0,94,0,0,0,0,0,43,0,29,0,145,0,182,0,133,0,221,0,142,0,102,0,0,0,241,0,74,0,38,0,0,0,184,0,228,0,79,0,212,0,0,0,207,0,42,0,14,0,1,0,105,0,5,0,0,0,103,0,74,0,49,0,0,0,130,0,0,0,66,0,192,0,0,0,156,0,0,0,215,0,88,0,29,0,89,0,84,0,0,0,86,0,36,0,85,0,115,0,46,0,160,0,0,0,249,0,196,0,0,0,173,0,0,0,0,0,121,0,41,0,231,0,0,0,62,0,43,0,150,0,215,0,132,0,19,0,94,0,193,0,33,0,0,0,0,0,225,0,120,0,77,0,198,0,118,0,98,0,213,0,238,0,112,0,0,0,234,0,93,0,175,0,39,0,33,0,28,0,248,0,224,0,35,0,159,0,119,0,93,0,0,0,115,0,220,0,83,0,0,0,95,0,158,0,231,0,32,0,135,0,201,0,0,0,196,0,71,0,0,0,0,0,0,0,127,0,143,0,0,0,34,0,113,0,0,0,0,0,58,0,121,0,0,0,223,0,0,0,181,0,253,0,78,0,104,0,34,0,162,0,163,0,91,0,75,0,52,0,218,0,0,0,164,0,89,0,213,0,252,0,117,0,0,0,46,0,102,0,246,0,0,0,97,0,28,0,116,0,252,0,81,0,0,0,122,0,105,0,156,0,90,0,0,0,61,0,71,0,229,0,0,0,119,0,21,0,77,0,75,0,72,0,111,0,137,0,0,0,135,0,126,0,84,0,187,0,211,0,26,0,0,0,127,0,15,0,0,0,238,0,26,0,0,0,64,0,0,0,201,0,57,0,124,0,0,0,125,0,10,0,222,0,230,0,206,0,136,0,3,0,137,0,179,0,14,0,65,0,93,0,213,0,0,0,116,0,93,0,201,0,70,0,120,0,209,0,16,0,173,0,248,0,96,0,74,0,118,0,74,0,143,0,0,0,144,0,207,0,0,0,0,0,153,0,95,0,29,0,47,0,50,0,114,0,51,0,140,0,0,0,0,0,42,0,155,0,254,0,0,0,251,0,176,0,237,0,136,0,184,0,0,0,107,0,79,0,16,0,104,0,0,0,197,0,0,0,0,0,0,0,82,0,71,0,110,0,193,0,34,0,154,0,246,0,38,0,0,0,245,0,120,0,0,0,14,0,38,0,9,0,81,0,218,0,12,0,0,0,170,0,76,0,71,0,84,0,70,0,99,0,241,0,34,0,51,0,10,0,0,0,107,0,0,0,0,0,0,0,159,0,0,0,0,0,210,0,89,0,33,0,144,0,171,0,0,0,0,0,42,0,102,0,12,0,0,0,190,0,72,0,76,0,19,0,99,0,42,0,0,0,18,0,146,0,55,0,151,0,0,0,189,0,0,0,203,0,216,0,28,0,244,0,240,0,0,0,38,0,2,0,0,0,0,0,148,0,225,0,60,0,241,0,26,0,0,0,0,0,10,0,53,0,113,0,169,0,102,0,208,0,46,0,17,0,0,0,226,0,0,0,0,0,0,0,106,0,39,0,0,0,0,0,0,0,222,0,41,0,52,0,0,0,238,0,232,0,43,0,245,0,154,0,200,0,65,0,82,0,56,0,193,0,192,0,239,0,130,0,164,0,0,0,34,0,141,0,0,0,179,0,0,0,124,0,143,0,169,0,227,0,58,0,0,0,110,0,20,0,201,0,202,0,17,0,116,0,181,0,226,0,0,0,127,0,0,0,52,0,215,0,139,0,180,0,0,0,0,0,248,0,31,0,22,0,195,0,107,0,53,0,106,0,194,0,131,0,235,0,0,0,76,0,126,0,148,0,148,0,218,0,116,0,48,0,0,0,161,0,151,0,71,0,0,0,198,0,106,0,78,0,152,0,211,0,0,0,64,0,0,0,184,0,129,0,242,0,28,0,160,0,0,0,0,0,0,0,167,0,63,0,198,0,76,0,192,0,0,0,0,0,0,0,0,0,0,0,214,0,249,0,225,0,187,0,0,0,49,0,207,0,182,0,115,0,199,0,132,0,0,0,45,0,41,0,124,0,187,0,85,0,193,0,0,0,103,0,122,0,0,0,224,0,87,0,51,0,6,0,214,0,41,0,168,0,143,0,182,0,180,0,25,0,146,0,147,0,125,0,230,0,14,0,117,0,58,0,143,0,119,0,0,0,0,0,157,0,195,0,161,0,55,0,101,0,0,0,0,0,243,0,16,0,247,0,85,0,0,0,12,0,154,0,21,0,57,0,0,0,235,0,0,0,252,0,115,0,118,0,41,0,127,0,219,0,0,0,90,0,102,0,83,0,132,0,0,0,127,0,205,0,0,0,200,0,0,0,82,0,0,0,156,0,101,0,242,0,240,0,103,0,187,0,0,0,106,0,0,0,195,0,98,0,52,0,0,0,19,0,74,0,234,0,229,0,0,0,68,0,208,0,23,0,0,0,0,0,75,0,217,0,29,0,208,0,0,0,0,0,133,0,246,0,0,0,89,0,81,0,205,0,218,0,193,0,91,0,243,0,155,0,226,0,117,0,85,0,132,0,128,0,0,0,179,0,26,0,88,0,136,0,113,0,0,0,240,0,0,0,43,0,88,0,106,0,145,0,0,0,98,0,236,0,0,0,94,0,47,0,45,0,55,0,0,0,94,0,118,0,122,0,0,0,135,0,125,0);
signal scenario_full  : scenario_type := (209,31,149,31,149,30,149,29,225,31,254,31,178,31,29,31,113,31,113,30,135,31,135,30,248,31,73,31,73,30,84,31,89,31,138,31,60,31,60,30,52,31,52,30,52,29,69,31,69,30,82,31,35,31,195,31,195,30,90,31,167,31,213,31,54,31,16,31,162,31,162,30,162,29,162,28,162,27,219,31,248,31,23,31,243,31,125,31,93,31,87,31,159,31,1,31,138,31,138,30,143,31,143,30,102,31,101,31,101,30,101,29,101,28,10,31,230,31,69,31,101,31,44,31,25,31,115,31,233,31,155,31,155,30,85,31,85,30,200,31,200,30,1,31,1,30,169,31,111,31,111,30,157,31,157,30,232,31,116,31,249,31,249,30,49,31,172,31,20,31,244,31,201,31,227,31,166,31,166,30,137,31,137,30,99,31,210,31,143,31,194,31,229,31,229,30,153,31,153,30,153,29,225,31,225,30,100,31,21,31,21,30,128,31,108,31,9,31,138,31,237,31,237,30,237,29,237,28,136,31,136,30,249,31,9,31,236,31,203,31,28,31,34,31,111,31,111,30,62,31,13,31,6,31,69,31,123,31,91,31,94,31,94,30,94,29,43,31,29,31,145,31,182,31,133,31,221,31,142,31,102,31,102,30,241,31,74,31,38,31,38,30,184,31,228,31,79,31,212,31,212,30,207,31,42,31,14,31,1,31,105,31,5,31,5,30,103,31,74,31,49,31,49,30,130,31,130,30,66,31,192,31,192,30,156,31,156,30,215,31,88,31,29,31,89,31,84,31,84,30,86,31,36,31,85,31,115,31,46,31,160,31,160,30,249,31,196,31,196,30,173,31,173,30,173,29,121,31,41,31,231,31,231,30,62,31,43,31,150,31,215,31,132,31,19,31,94,31,193,31,33,31,33,30,33,29,225,31,120,31,77,31,198,31,118,31,98,31,213,31,238,31,112,31,112,30,234,31,93,31,175,31,39,31,33,31,28,31,248,31,224,31,35,31,159,31,119,31,93,31,93,30,115,31,220,31,83,31,83,30,95,31,158,31,231,31,32,31,135,31,201,31,201,30,196,31,71,31,71,30,71,29,71,28,127,31,143,31,143,30,34,31,113,31,113,30,113,29,58,31,121,31,121,30,223,31,223,30,181,31,253,31,78,31,104,31,34,31,162,31,163,31,91,31,75,31,52,31,218,31,218,30,164,31,89,31,213,31,252,31,117,31,117,30,46,31,102,31,246,31,246,30,97,31,28,31,116,31,252,31,81,31,81,30,122,31,105,31,156,31,90,31,90,30,61,31,71,31,229,31,229,30,119,31,21,31,77,31,75,31,72,31,111,31,137,31,137,30,135,31,126,31,84,31,187,31,211,31,26,31,26,30,127,31,15,31,15,30,238,31,26,31,26,30,64,31,64,30,201,31,57,31,124,31,124,30,125,31,10,31,222,31,230,31,206,31,136,31,3,31,137,31,179,31,14,31,65,31,93,31,213,31,213,30,116,31,93,31,201,31,70,31,120,31,209,31,16,31,173,31,248,31,96,31,74,31,118,31,74,31,143,31,143,30,144,31,207,31,207,30,207,29,153,31,95,31,29,31,47,31,50,31,114,31,51,31,140,31,140,30,140,29,42,31,155,31,254,31,254,30,251,31,176,31,237,31,136,31,184,31,184,30,107,31,79,31,16,31,104,31,104,30,197,31,197,30,197,29,197,28,82,31,71,31,110,31,193,31,34,31,154,31,246,31,38,31,38,30,245,31,120,31,120,30,14,31,38,31,9,31,81,31,218,31,12,31,12,30,170,31,76,31,71,31,84,31,70,31,99,31,241,31,34,31,51,31,10,31,10,30,107,31,107,30,107,29,107,28,159,31,159,30,159,29,210,31,89,31,33,31,144,31,171,31,171,30,171,29,42,31,102,31,12,31,12,30,190,31,72,31,76,31,19,31,99,31,42,31,42,30,18,31,146,31,55,31,151,31,151,30,189,31,189,30,203,31,216,31,28,31,244,31,240,31,240,30,38,31,2,31,2,30,2,29,148,31,225,31,60,31,241,31,26,31,26,30,26,29,10,31,53,31,113,31,169,31,102,31,208,31,46,31,17,31,17,30,226,31,226,30,226,29,226,28,106,31,39,31,39,30,39,29,39,28,222,31,41,31,52,31,52,30,238,31,232,31,43,31,245,31,154,31,200,31,65,31,82,31,56,31,193,31,192,31,239,31,130,31,164,31,164,30,34,31,141,31,141,30,179,31,179,30,124,31,143,31,169,31,227,31,58,31,58,30,110,31,20,31,201,31,202,31,17,31,116,31,181,31,226,31,226,30,127,31,127,30,52,31,215,31,139,31,180,31,180,30,180,29,248,31,31,31,22,31,195,31,107,31,53,31,106,31,194,31,131,31,235,31,235,30,76,31,126,31,148,31,148,31,218,31,116,31,48,31,48,30,161,31,151,31,71,31,71,30,198,31,106,31,78,31,152,31,211,31,211,30,64,31,64,30,184,31,129,31,242,31,28,31,160,31,160,30,160,29,160,28,167,31,63,31,198,31,76,31,192,31,192,30,192,29,192,28,192,27,192,26,214,31,249,31,225,31,187,31,187,30,49,31,207,31,182,31,115,31,199,31,132,31,132,30,45,31,41,31,124,31,187,31,85,31,193,31,193,30,103,31,122,31,122,30,224,31,87,31,51,31,6,31,214,31,41,31,168,31,143,31,182,31,180,31,25,31,146,31,147,31,125,31,230,31,14,31,117,31,58,31,143,31,119,31,119,30,119,29,157,31,195,31,161,31,55,31,101,31,101,30,101,29,243,31,16,31,247,31,85,31,85,30,12,31,154,31,21,31,57,31,57,30,235,31,235,30,252,31,115,31,118,31,41,31,127,31,219,31,219,30,90,31,102,31,83,31,132,31,132,30,127,31,205,31,205,30,200,31,200,30,82,31,82,30,156,31,101,31,242,31,240,31,103,31,187,31,187,30,106,31,106,30,195,31,98,31,52,31,52,30,19,31,74,31,234,31,229,31,229,30,68,31,208,31,23,31,23,30,23,29,75,31,217,31,29,31,208,31,208,30,208,29,133,31,246,31,246,30,89,31,81,31,205,31,218,31,193,31,91,31,243,31,155,31,226,31,117,31,85,31,132,31,128,31,128,30,179,31,26,31,88,31,136,31,113,31,113,30,240,31,240,30,43,31,88,31,106,31,145,31,145,30,98,31,236,31,236,30,94,31,47,31,45,31,55,31,55,30,94,31,118,31,122,31,122,30,135,31,125,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
