-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 168;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (12,0,178,0,0,0,116,0,233,0,81,0,49,0,0,0,195,0,159,0,227,0,201,0,215,0,90,0,0,0,6,0,135,0,64,0,0,0,139,0,51,0,68,0,0,0,0,0,157,0,0,0,233,0,57,0,184,0,92,0,47,0,207,0,110,0,4,0,144,0,213,0,195,0,0,0,0,0,26,0,181,0,0,0,0,0,41,0,249,0,0,0,233,0,45,0,3,0,0,0,77,0,176,0,96,0,0,0,198,0,74,0,48,0,99,0,60,0,92,0,0,0,162,0,199,0,11,0,192,0,1,0,242,0,54,0,0,0,200,0,190,0,72,0,124,0,50,0,69,0,0,0,114,0,36,0,181,0,199,0,1,0,237,0,0,0,123,0,223,0,26,0,0,0,30,0,6,0,5,0,97,0,55,0,27,0,0,0,194,0,173,0,0,0,0,0,247,0,76,0,221,0,129,0,130,0,34,0,0,0,51,0,158,0,177,0,135,0,252,0,113,0,137,0,120,0,108,0,109,0,209,0,180,0,171,0,0,0,6,0,0,0,171,0,176,0,236,0,0,0,1,0,236,0,0,0,142,0,103,0,116,0,75,0,198,0,114,0,183,0,91,0,0,0,210,0,0,0,141,0,0,0,0,0,240,0,131,0,175,0,84,0,145,0,0,0,120,0,0,0,75,0,0,0,217,0,245,0,64,0,19,0,228,0,40,0,164,0,0,0,242,0,83,0,0,0,121,0,242,0,223,0,197,0,59,0);
signal scenario_full  : scenario_type := (12,31,178,31,178,30,116,31,233,31,81,31,49,31,49,30,195,31,159,31,227,31,201,31,215,31,90,31,90,30,6,31,135,31,64,31,64,30,139,31,51,31,68,31,68,30,68,29,157,31,157,30,233,31,57,31,184,31,92,31,47,31,207,31,110,31,4,31,144,31,213,31,195,31,195,30,195,29,26,31,181,31,181,30,181,29,41,31,249,31,249,30,233,31,45,31,3,31,3,30,77,31,176,31,96,31,96,30,198,31,74,31,48,31,99,31,60,31,92,31,92,30,162,31,199,31,11,31,192,31,1,31,242,31,54,31,54,30,200,31,190,31,72,31,124,31,50,31,69,31,69,30,114,31,36,31,181,31,199,31,1,31,237,31,237,30,123,31,223,31,26,31,26,30,30,31,6,31,5,31,97,31,55,31,27,31,27,30,194,31,173,31,173,30,173,29,247,31,76,31,221,31,129,31,130,31,34,31,34,30,51,31,158,31,177,31,135,31,252,31,113,31,137,31,120,31,108,31,109,31,209,31,180,31,171,31,171,30,6,31,6,30,171,31,176,31,236,31,236,30,1,31,236,31,236,30,142,31,103,31,116,31,75,31,198,31,114,31,183,31,91,31,91,30,210,31,210,30,141,31,141,30,141,29,240,31,131,31,175,31,84,31,145,31,145,30,120,31,120,30,75,31,75,30,217,31,245,31,64,31,19,31,228,31,40,31,164,31,164,30,242,31,83,31,83,30,121,31,242,31,223,31,197,31,59,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
