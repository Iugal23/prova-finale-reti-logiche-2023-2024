-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_761 is
end project_tb_761;

architecture project_tb_arch_761 of project_tb_761 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 801;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (195,0,73,0,37,0,140,0,157,0,42,0,240,0,161,0,71,0,87,0,209,0,0,0,110,0,90,0,15,0,80,0,102,0,202,0,127,0,170,0,3,0,4,0,193,0,0,0,116,0,147,0,0,0,40,0,27,0,0,0,169,0,0,0,64,0,103,0,231,0,0,0,182,0,50,0,175,0,107,0,197,0,167,0,182,0,159,0,165,0,0,0,254,0,116,0,204,0,103,0,13,0,65,0,76,0,167,0,179,0,229,0,229,0,147,0,83,0,4,0,162,0,136,0,179,0,94,0,92,0,0,0,0,0,200,0,5,0,0,0,44,0,0,0,181,0,0,0,123,0,0,0,95,0,191,0,220,0,0,0,107,0,18,0,24,0,0,0,0,0,255,0,93,0,159,0,227,0,129,0,33,0,223,0,79,0,250,0,2,0,50,0,77,0,27,0,133,0,209,0,134,0,169,0,255,0,11,0,13,0,118,0,200,0,215,0,0,0,0,0,154,0,125,0,0,0,166,0,0,0,73,0,0,0,38,0,225,0,157,0,148,0,39,0,149,0,70,0,22,0,54,0,82,0,254,0,62,0,181,0,163,0,174,0,145,0,201,0,0,0,112,0,44,0,1,0,95,0,125,0,185,0,4,0,194,0,223,0,87,0,164,0,76,0,21,0,195,0,0,0,133,0,113,0,254,0,199,0,36,0,26,0,45,0,152,0,62,0,207,0,142,0,129,0,11,0,224,0,198,0,240,0,0,0,102,0,0,0,131,0,78,0,131,0,12,0,98,0,93,0,160,0,32,0,3,0,99,0,1,0,109,0,144,0,0,0,198,0,89,0,134,0,19,0,40,0,5,0,0,0,0,0,116,0,0,0,0,0,169,0,63,0,122,0,150,0,170,0,0,0,140,0,146,0,244,0,115,0,127,0,63,0,0,0,250,0,0,0,0,0,63,0,157,0,61,0,0,0,145,0,157,0,194,0,0,0,0,0,90,0,68,0,0,0,113,0,226,0,171,0,0,0,0,0,199,0,0,0,175,0,0,0,40,0,0,0,203,0,236,0,123,0,0,0,125,0,91,0,96,0,0,0,124,0,121,0,222,0,183,0,136,0,142,0,236,0,21,0,0,0,48,0,89,0,181,0,241,0,88,0,37,0,201,0,106,0,0,0,121,0,0,0,246,0,86,0,189,0,151,0,212,0,25,0,0,0,219,0,0,0,117,0,236,0,211,0,167,0,233,0,89,0,196,0,25,0,78,0,79,0,144,0,13,0,246,0,178,0,196,0,111,0,0,0,0,0,252,0,227,0,59,0,7,0,215,0,135,0,3,0,0,0,157,0,0,0,132,0,12,0,165,0,151,0,56,0,0,0,240,0,7,0,165,0,191,0,202,0,33,0,164,0,105,0,0,0,177,0,223,0,0,0,212,0,12,0,0,0,55,0,1,0,134,0,0,0,219,0,47,0,249,0,71,0,166,0,247,0,99,0,207,0,196,0,0,0,0,0,0,0,49,0,166,0,251,0,147,0,28,0,195,0,14,0,116,0,148,0,0,0,0,0,114,0,0,0,48,0,135,0,45,0,88,0,10,0,0,0,44,0,7,0,169,0,108,0,205,0,130,0,193,0,181,0,117,0,218,0,238,0,208,0,248,0,175,0,60,0,36,0,223,0,108,0,16,0,255,0,11,0,76,0,165,0,133,0,0,0,216,0,130,0,80,0,1,0,37,0,0,0,147,0,24,0,0,0,81,0,41,0,22,0,201,0,44,0,166,0,206,0,0,0,204,0,125,0,42,0,20,0,199,0,0,0,255,0,50,0,230,0,196,0,0,0,63,0,155,0,180,0,0,0,28,0,147,0,176,0,0,0,0,0,206,0,10,0,227,0,182,0,145,0,106,0,0,0,171,0,14,0,0,0,0,0,0,0,78,0,0,0,185,0,29,0,69,0,94,0,226,0,0,0,85,0,231,0,0,0,177,0,121,0,217,0,25,0,207,0,0,0,69,0,190,0,74,0,160,0,179,0,18,0,0,0,117,0,142,0,97,0,148,0,83,0,22,0,0,0,238,0,250,0,42,0,48,0,0,0,79,0,194,0,187,0,0,0,110,0,68,0,118,0,230,0,134,0,186,0,37,0,0,0,253,0,125,0,0,0,219,0,175,0,0,0,189,0,137,0,21,0,0,0,101,0,57,0,0,0,159,0,0,0,127,0,126,0,11,0,0,0,6,0,242,0,128,0,201,0,0,0,0,0,0,0,233,0,174,0,0,0,238,0,205,0,239,0,73,0,125,0,155,0,8,0,167,0,2,0,0,0,85,0,95,0,114,0,0,0,135,0,26,0,186,0,94,0,51,0,0,0,154,0,112,0,0,0,43,0,137,0,192,0,168,0,0,0,0,0,0,0,161,0,172,0,0,0,127,0,249,0,60,0,142,0,0,0,0,0,64,0,11,0,10,0,171,0,0,0,87,0,22,0,151,0,0,0,86,0,0,0,221,0,86,0,154,0,0,0,151,0,0,0,142,0,188,0,18,0,223,0,45,0,113,0,157,0,187,0,58,0,158,0,238,0,0,0,0,0,47,0,152,0,219,0,92,0,224,0,0,0,0,0,132,0,0,0,213,0,226,0,29,0,51,0,141,0,14,0,0,0,0,0,69,0,159,0,142,0,101,0,211,0,76,0,0,0,0,0,175,0,180,0,3,0,0,0,157,0,160,0,8,0,0,0,229,0,224,0,208,0,133,0,82,0,115,0,170,0,44,0,87,0,0,0,19,0,0,0,0,0,98,0,14,0,149,0,65,0,0,0,248,0,37,0,155,0,163,0,0,0,245,0,81,0,0,0,3,0,0,0,208,0,78,0,0,0,40,0,99,0,0,0,7,0,216,0,57,0,64,0,131,0,51,0,143,0,163,0,183,0,71,0,88,0,136,0,0,0,191,0,0,0,68,0,229,0,60,0,251,0,34,0,162,0,0,0,21,0,149,0,0,0,51,0,201,0,74,0,196,0,232,0,140,0,0,0,19,0,151,0,142,0,216,0,0,0,78,0,79,0,82,0,0,0,248,0,223,0,0,0,0,0,252,0,0,0,91,0,139,0,182,0,0,0,24,0,61,0,176,0,251,0,219,0,143,0,184,0,0,0,155,0,167,0,224,0,220,0,0,0,76,0,165,0,122,0,101,0,125,0,139,0,0,0,39,0,144,0,0,0,26,0,27,0,0,0,73,0,179,0,89,0,148,0,207,0,12,0,150,0,184,0,29,0,234,0,173,0,223,0,127,0,192,0,210,0,18,0,0,0,48,0,151,0,166,0,0,0,0,0,0,0,28,0,146,0,212,0,39,0,83,0,85,0,68,0,34,0,63,0,176,0,0,0,0,0,163,0,76,0,223,0,0,0,238,0,0,0,159,0,0,0,0,0,205,0,225,0,213,0,174,0,136,0,40,0,58,0,244,0,251,0,0,0,0,0,62,0,67,0,123,0,247,0,25,0,252,0,212,0,0,0,179,0,55,0,67,0,232,0,98,0,61,0,0,0,119,0,197,0,128,0,240,0,174,0,2,0,129,0,50,0,135,0,0,0,59,0,54,0,195,0);
signal scenario_full  : scenario_type := (195,31,73,31,37,31,140,31,157,31,42,31,240,31,161,31,71,31,87,31,209,31,209,30,110,31,90,31,15,31,80,31,102,31,202,31,127,31,170,31,3,31,4,31,193,31,193,30,116,31,147,31,147,30,40,31,27,31,27,30,169,31,169,30,64,31,103,31,231,31,231,30,182,31,50,31,175,31,107,31,197,31,167,31,182,31,159,31,165,31,165,30,254,31,116,31,204,31,103,31,13,31,65,31,76,31,167,31,179,31,229,31,229,31,147,31,83,31,4,31,162,31,136,31,179,31,94,31,92,31,92,30,92,29,200,31,5,31,5,30,44,31,44,30,181,31,181,30,123,31,123,30,95,31,191,31,220,31,220,30,107,31,18,31,24,31,24,30,24,29,255,31,93,31,159,31,227,31,129,31,33,31,223,31,79,31,250,31,2,31,50,31,77,31,27,31,133,31,209,31,134,31,169,31,255,31,11,31,13,31,118,31,200,31,215,31,215,30,215,29,154,31,125,31,125,30,166,31,166,30,73,31,73,30,38,31,225,31,157,31,148,31,39,31,149,31,70,31,22,31,54,31,82,31,254,31,62,31,181,31,163,31,174,31,145,31,201,31,201,30,112,31,44,31,1,31,95,31,125,31,185,31,4,31,194,31,223,31,87,31,164,31,76,31,21,31,195,31,195,30,133,31,113,31,254,31,199,31,36,31,26,31,45,31,152,31,62,31,207,31,142,31,129,31,11,31,224,31,198,31,240,31,240,30,102,31,102,30,131,31,78,31,131,31,12,31,98,31,93,31,160,31,32,31,3,31,99,31,1,31,109,31,144,31,144,30,198,31,89,31,134,31,19,31,40,31,5,31,5,30,5,29,116,31,116,30,116,29,169,31,63,31,122,31,150,31,170,31,170,30,140,31,146,31,244,31,115,31,127,31,63,31,63,30,250,31,250,30,250,29,63,31,157,31,61,31,61,30,145,31,157,31,194,31,194,30,194,29,90,31,68,31,68,30,113,31,226,31,171,31,171,30,171,29,199,31,199,30,175,31,175,30,40,31,40,30,203,31,236,31,123,31,123,30,125,31,91,31,96,31,96,30,124,31,121,31,222,31,183,31,136,31,142,31,236,31,21,31,21,30,48,31,89,31,181,31,241,31,88,31,37,31,201,31,106,31,106,30,121,31,121,30,246,31,86,31,189,31,151,31,212,31,25,31,25,30,219,31,219,30,117,31,236,31,211,31,167,31,233,31,89,31,196,31,25,31,78,31,79,31,144,31,13,31,246,31,178,31,196,31,111,31,111,30,111,29,252,31,227,31,59,31,7,31,215,31,135,31,3,31,3,30,157,31,157,30,132,31,12,31,165,31,151,31,56,31,56,30,240,31,7,31,165,31,191,31,202,31,33,31,164,31,105,31,105,30,177,31,223,31,223,30,212,31,12,31,12,30,55,31,1,31,134,31,134,30,219,31,47,31,249,31,71,31,166,31,247,31,99,31,207,31,196,31,196,30,196,29,196,28,49,31,166,31,251,31,147,31,28,31,195,31,14,31,116,31,148,31,148,30,148,29,114,31,114,30,48,31,135,31,45,31,88,31,10,31,10,30,44,31,7,31,169,31,108,31,205,31,130,31,193,31,181,31,117,31,218,31,238,31,208,31,248,31,175,31,60,31,36,31,223,31,108,31,16,31,255,31,11,31,76,31,165,31,133,31,133,30,216,31,130,31,80,31,1,31,37,31,37,30,147,31,24,31,24,30,81,31,41,31,22,31,201,31,44,31,166,31,206,31,206,30,204,31,125,31,42,31,20,31,199,31,199,30,255,31,50,31,230,31,196,31,196,30,63,31,155,31,180,31,180,30,28,31,147,31,176,31,176,30,176,29,206,31,10,31,227,31,182,31,145,31,106,31,106,30,171,31,14,31,14,30,14,29,14,28,78,31,78,30,185,31,29,31,69,31,94,31,226,31,226,30,85,31,231,31,231,30,177,31,121,31,217,31,25,31,207,31,207,30,69,31,190,31,74,31,160,31,179,31,18,31,18,30,117,31,142,31,97,31,148,31,83,31,22,31,22,30,238,31,250,31,42,31,48,31,48,30,79,31,194,31,187,31,187,30,110,31,68,31,118,31,230,31,134,31,186,31,37,31,37,30,253,31,125,31,125,30,219,31,175,31,175,30,189,31,137,31,21,31,21,30,101,31,57,31,57,30,159,31,159,30,127,31,126,31,11,31,11,30,6,31,242,31,128,31,201,31,201,30,201,29,201,28,233,31,174,31,174,30,238,31,205,31,239,31,73,31,125,31,155,31,8,31,167,31,2,31,2,30,85,31,95,31,114,31,114,30,135,31,26,31,186,31,94,31,51,31,51,30,154,31,112,31,112,30,43,31,137,31,192,31,168,31,168,30,168,29,168,28,161,31,172,31,172,30,127,31,249,31,60,31,142,31,142,30,142,29,64,31,11,31,10,31,171,31,171,30,87,31,22,31,151,31,151,30,86,31,86,30,221,31,86,31,154,31,154,30,151,31,151,30,142,31,188,31,18,31,223,31,45,31,113,31,157,31,187,31,58,31,158,31,238,31,238,30,238,29,47,31,152,31,219,31,92,31,224,31,224,30,224,29,132,31,132,30,213,31,226,31,29,31,51,31,141,31,14,31,14,30,14,29,69,31,159,31,142,31,101,31,211,31,76,31,76,30,76,29,175,31,180,31,3,31,3,30,157,31,160,31,8,31,8,30,229,31,224,31,208,31,133,31,82,31,115,31,170,31,44,31,87,31,87,30,19,31,19,30,19,29,98,31,14,31,149,31,65,31,65,30,248,31,37,31,155,31,163,31,163,30,245,31,81,31,81,30,3,31,3,30,208,31,78,31,78,30,40,31,99,31,99,30,7,31,216,31,57,31,64,31,131,31,51,31,143,31,163,31,183,31,71,31,88,31,136,31,136,30,191,31,191,30,68,31,229,31,60,31,251,31,34,31,162,31,162,30,21,31,149,31,149,30,51,31,201,31,74,31,196,31,232,31,140,31,140,30,19,31,151,31,142,31,216,31,216,30,78,31,79,31,82,31,82,30,248,31,223,31,223,30,223,29,252,31,252,30,91,31,139,31,182,31,182,30,24,31,61,31,176,31,251,31,219,31,143,31,184,31,184,30,155,31,167,31,224,31,220,31,220,30,76,31,165,31,122,31,101,31,125,31,139,31,139,30,39,31,144,31,144,30,26,31,27,31,27,30,73,31,179,31,89,31,148,31,207,31,12,31,150,31,184,31,29,31,234,31,173,31,223,31,127,31,192,31,210,31,18,31,18,30,48,31,151,31,166,31,166,30,166,29,166,28,28,31,146,31,212,31,39,31,83,31,85,31,68,31,34,31,63,31,176,31,176,30,176,29,163,31,76,31,223,31,223,30,238,31,238,30,159,31,159,30,159,29,205,31,225,31,213,31,174,31,136,31,40,31,58,31,244,31,251,31,251,30,251,29,62,31,67,31,123,31,247,31,25,31,252,31,212,31,212,30,179,31,55,31,67,31,232,31,98,31,61,31,61,30,119,31,197,31,128,31,240,31,174,31,2,31,129,31,50,31,135,31,135,30,59,31,54,31,195,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
