-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_418 is
end project_tb_418;

architecture project_tb_arch_418 of project_tb_418 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 628;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,58,0,50,0,19,0,0,0,150,0,49,0,72,0,137,0,67,0,78,0,226,0,124,0,86,0,126,0,169,0,130,0,44,0,237,0,0,0,61,0,0,0,24,0,216,0,135,0,122,0,205,0,57,0,178,0,159,0,138,0,236,0,166,0,191,0,0,0,50,0,236,0,0,0,0,0,71,0,104,0,0,0,9,0,25,0,128,0,28,0,77,0,45,0,0,0,163,0,94,0,0,0,116,0,181,0,0,0,165,0,67,0,0,0,101,0,0,0,139,0,224,0,0,0,208,0,95,0,31,0,29,0,127,0,4,0,251,0,0,0,164,0,233,0,91,0,55,0,128,0,111,0,77,0,184,0,89,0,83,0,0,0,0,0,36,0,7,0,0,0,142,0,0,0,0,0,101,0,0,0,113,0,207,0,133,0,83,0,153,0,154,0,109,0,163,0,2,0,140,0,190,0,29,0,4,0,40,0,9,0,180,0,24,0,133,0,0,0,253,0,131,0,162,0,118,0,0,0,101,0,146,0,253,0,21,0,0,0,144,0,48,0,119,0,0,0,62,0,142,0,0,0,118,0,132,0,61,0,242,0,210,0,253,0,60,0,48,0,0,0,178,0,0,0,128,0,221,0,179,0,154,0,128,0,21,0,0,0,94,0,50,0,137,0,0,0,4,0,241,0,96,0,80,0,99,0,130,0,137,0,145,0,53,0,71,0,0,0,236,0,163,0,0,0,239,0,149,0,0,0,211,0,77,0,134,0,0,0,140,0,54,0,0,0,65,0,177,0,87,0,201,0,51,0,138,0,0,0,224,0,0,0,179,0,0,0,16,0,102,0,235,0,133,0,9,0,0,0,58,0,134,0,18,0,183,0,0,0,18,0,226,0,250,0,0,0,18,0,220,0,120,0,180,0,0,0,0,0,0,0,16,0,115,0,0,0,151,0,0,0,18,0,246,0,0,0,0,0,0,0,250,0,36,0,243,0,16,0,202,0,42,0,232,0,251,0,1,0,0,0,177,0,97,0,30,0,132,0,0,0,207,0,255,0,74,0,204,0,148,0,0,0,121,0,103,0,154,0,155,0,216,0,242,0,250,0,119,0,197,0,0,0,223,0,95,0,193,0,137,0,71,0,213,0,92,0,187,0,41,0,66,0,119,0,0,0,104,0,0,0,195,0,24,0,166,0,0,0,0,0,0,0,215,0,232,0,0,0,107,0,26,0,165,0,154,0,0,0,0,0,65,0,147,0,228,0,168,0,48,0,191,0,2,0,92,0,72,0,155,0,0,0,112,0,190,0,66,0,206,0,228,0,90,0,194,0,0,0,219,0,176,0,241,0,179,0,0,0,76,0,0,0,117,0,109,0,120,0,0,0,186,0,213,0,0,0,224,0,134,0,126,0,78,0,38,0,0,0,195,0,0,0,8,0,199,0,0,0,116,0,0,0,0,0,0,0,210,0,0,0,148,0,128,0,153,0,0,0,19,0,190,0,6,0,66,0,29,0,147,0,193,0,0,0,49,0,177,0,100,0,217,0,27,0,224,0,170,0,31,0,182,0,152,0,147,0,112,0,96,0,106,0,0,0,254,0,190,0,73,0,0,0,231,0,176,0,60,0,152,0,40,0,187,0,0,0,0,0,91,0,72,0,93,0,136,0,97,0,97,0,152,0,57,0,159,0,0,0,84,0,45,0,180,0,225,0,98,0,0,0,0,0,144,0,119,0,38,0,187,0,138,0,85,0,130,0,164,0,0,0,194,0,173,0,234,0,0,0,110,0,193,0,115,0,224,0,242,0,126,0,0,0,225,0,72,0,0,0,40,0,143,0,185,0,27,0,0,0,158,0,0,0,8,0,6,0,29,0,223,0,40,0,4,0,0,0,173,0,76,0,99,0,39,0,113,0,154,0,184,0,97,0,0,0,18,0,247,0,35,0,16,0,121,0,0,0,167,0,9,0,150,0,171,0,188,0,140,0,62,0,21,0,105,0,95,0,0,0,121,0,23,0,162,0,96,0,214,0,134,0,1,0,81,0,63,0,126,0,125,0,66,0,218,0,75,0,202,0,182,0,93,0,178,0,0,0,224,0,76,0,241,0,56,0,242,0,171,0,44,0,80,0,223,0,135,0,51,0,119,0,0,0,145,0,0,0,247,0,189,0,250,0,26,0,39,0,196,0,186,0,205,0,210,0,235,0,40,0,201,0,186,0,0,0,9,0,134,0,189,0,137,0,252,0,220,0,139,0,0,0,0,0,176,0,0,0,122,0,36,0,205,0,123,0,172,0,51,0,0,0,246,0,115,0,0,0,199,0,134,0,125,0,0,0,5,0,100,0,181,0,142,0,137,0,0,0,47,0,0,0,148,0,86,0,104,0,168,0,81,0,79,0,75,0,106,0,234,0,6,0,0,0,175,0,51,0,151,0,211,0,48,0,42,0,90,0,224,0,140,0,0,0,0,0,253,0,221,0,180,0,0,0,80,0,30,0,194,0,110,0,77,0,114,0,0,0,132,0,94,0,140,0,91,0,153,0,238,0,128,0,187,0,62,0,26,0,0,0,150,0,22,0,250,0,77,0,35,0,169,0,19,0,85,0,252,0,66,0,149,0,0,0,0,0,0,0,214,0,203,0,24,0,220,0,0,0,52,0,243,0,0,0,19,0,115,0,91,0,248,0,27,0,218,0,0,0,240,0,43,0,42,0,70,0,121,0,0,0,226,0,146,0,153,0,199,0,137,0,199,0,124,0,147,0,84,0,13,0,128,0,245,0,0,0,131,0,0,0,194,0,0,0,244,0,56,0,6,0,200,0,0,0,55,0);
signal scenario_full  : scenario_type := (0,0,58,31,50,31,19,31,19,30,150,31,49,31,72,31,137,31,67,31,78,31,226,31,124,31,86,31,126,31,169,31,130,31,44,31,237,31,237,30,61,31,61,30,24,31,216,31,135,31,122,31,205,31,57,31,178,31,159,31,138,31,236,31,166,31,191,31,191,30,50,31,236,31,236,30,236,29,71,31,104,31,104,30,9,31,25,31,128,31,28,31,77,31,45,31,45,30,163,31,94,31,94,30,116,31,181,31,181,30,165,31,67,31,67,30,101,31,101,30,139,31,224,31,224,30,208,31,95,31,31,31,29,31,127,31,4,31,251,31,251,30,164,31,233,31,91,31,55,31,128,31,111,31,77,31,184,31,89,31,83,31,83,30,83,29,36,31,7,31,7,30,142,31,142,30,142,29,101,31,101,30,113,31,207,31,133,31,83,31,153,31,154,31,109,31,163,31,2,31,140,31,190,31,29,31,4,31,40,31,9,31,180,31,24,31,133,31,133,30,253,31,131,31,162,31,118,31,118,30,101,31,146,31,253,31,21,31,21,30,144,31,48,31,119,31,119,30,62,31,142,31,142,30,118,31,132,31,61,31,242,31,210,31,253,31,60,31,48,31,48,30,178,31,178,30,128,31,221,31,179,31,154,31,128,31,21,31,21,30,94,31,50,31,137,31,137,30,4,31,241,31,96,31,80,31,99,31,130,31,137,31,145,31,53,31,71,31,71,30,236,31,163,31,163,30,239,31,149,31,149,30,211,31,77,31,134,31,134,30,140,31,54,31,54,30,65,31,177,31,87,31,201,31,51,31,138,31,138,30,224,31,224,30,179,31,179,30,16,31,102,31,235,31,133,31,9,31,9,30,58,31,134,31,18,31,183,31,183,30,18,31,226,31,250,31,250,30,18,31,220,31,120,31,180,31,180,30,180,29,180,28,16,31,115,31,115,30,151,31,151,30,18,31,246,31,246,30,246,29,246,28,250,31,36,31,243,31,16,31,202,31,42,31,232,31,251,31,1,31,1,30,177,31,97,31,30,31,132,31,132,30,207,31,255,31,74,31,204,31,148,31,148,30,121,31,103,31,154,31,155,31,216,31,242,31,250,31,119,31,197,31,197,30,223,31,95,31,193,31,137,31,71,31,213,31,92,31,187,31,41,31,66,31,119,31,119,30,104,31,104,30,195,31,24,31,166,31,166,30,166,29,166,28,215,31,232,31,232,30,107,31,26,31,165,31,154,31,154,30,154,29,65,31,147,31,228,31,168,31,48,31,191,31,2,31,92,31,72,31,155,31,155,30,112,31,190,31,66,31,206,31,228,31,90,31,194,31,194,30,219,31,176,31,241,31,179,31,179,30,76,31,76,30,117,31,109,31,120,31,120,30,186,31,213,31,213,30,224,31,134,31,126,31,78,31,38,31,38,30,195,31,195,30,8,31,199,31,199,30,116,31,116,30,116,29,116,28,210,31,210,30,148,31,128,31,153,31,153,30,19,31,190,31,6,31,66,31,29,31,147,31,193,31,193,30,49,31,177,31,100,31,217,31,27,31,224,31,170,31,31,31,182,31,152,31,147,31,112,31,96,31,106,31,106,30,254,31,190,31,73,31,73,30,231,31,176,31,60,31,152,31,40,31,187,31,187,30,187,29,91,31,72,31,93,31,136,31,97,31,97,31,152,31,57,31,159,31,159,30,84,31,45,31,180,31,225,31,98,31,98,30,98,29,144,31,119,31,38,31,187,31,138,31,85,31,130,31,164,31,164,30,194,31,173,31,234,31,234,30,110,31,193,31,115,31,224,31,242,31,126,31,126,30,225,31,72,31,72,30,40,31,143,31,185,31,27,31,27,30,158,31,158,30,8,31,6,31,29,31,223,31,40,31,4,31,4,30,173,31,76,31,99,31,39,31,113,31,154,31,184,31,97,31,97,30,18,31,247,31,35,31,16,31,121,31,121,30,167,31,9,31,150,31,171,31,188,31,140,31,62,31,21,31,105,31,95,31,95,30,121,31,23,31,162,31,96,31,214,31,134,31,1,31,81,31,63,31,126,31,125,31,66,31,218,31,75,31,202,31,182,31,93,31,178,31,178,30,224,31,76,31,241,31,56,31,242,31,171,31,44,31,80,31,223,31,135,31,51,31,119,31,119,30,145,31,145,30,247,31,189,31,250,31,26,31,39,31,196,31,186,31,205,31,210,31,235,31,40,31,201,31,186,31,186,30,9,31,134,31,189,31,137,31,252,31,220,31,139,31,139,30,139,29,176,31,176,30,122,31,36,31,205,31,123,31,172,31,51,31,51,30,246,31,115,31,115,30,199,31,134,31,125,31,125,30,5,31,100,31,181,31,142,31,137,31,137,30,47,31,47,30,148,31,86,31,104,31,168,31,81,31,79,31,75,31,106,31,234,31,6,31,6,30,175,31,51,31,151,31,211,31,48,31,42,31,90,31,224,31,140,31,140,30,140,29,253,31,221,31,180,31,180,30,80,31,30,31,194,31,110,31,77,31,114,31,114,30,132,31,94,31,140,31,91,31,153,31,238,31,128,31,187,31,62,31,26,31,26,30,150,31,22,31,250,31,77,31,35,31,169,31,19,31,85,31,252,31,66,31,149,31,149,30,149,29,149,28,214,31,203,31,24,31,220,31,220,30,52,31,243,31,243,30,19,31,115,31,91,31,248,31,27,31,218,31,218,30,240,31,43,31,42,31,70,31,121,31,121,30,226,31,146,31,153,31,199,31,137,31,199,31,124,31,147,31,84,31,13,31,128,31,245,31,245,30,131,31,131,30,194,31,194,30,244,31,56,31,6,31,200,31,200,30,55,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
