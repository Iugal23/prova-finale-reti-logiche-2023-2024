-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_497 is
end project_tb_497;

architecture project_tb_arch_497 of project_tb_497 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 975;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (207,0,220,0,0,0,0,0,61,0,27,0,26,0,125,0,56,0,0,0,101,0,175,0,194,0,191,0,32,0,51,0,165,0,142,0,0,0,47,0,143,0,147,0,5,0,139,0,239,0,43,0,113,0,253,0,0,0,177,0,25,0,0,0,0,0,55,0,216,0,122,0,152,0,142,0,149,0,136,0,24,0,158,0,0,0,117,0,253,0,0,0,0,0,23,0,219,0,56,0,41,0,0,0,132,0,42,0,85,0,151,0,145,0,5,0,30,0,45,0,0,0,180,0,210,0,129,0,135,0,44,0,76,0,151,0,23,0,108,0,104,0,40,0,218,0,193,0,0,0,0,0,72,0,63,0,79,0,209,0,136,0,0,0,213,0,114,0,254,0,0,0,162,0,128,0,177,0,133,0,215,0,23,0,190,0,239,0,14,0,160,0,86,0,214,0,33,0,124,0,61,0,0,0,214,0,0,0,155,0,0,0,16,0,20,0,20,0,20,0,191,0,0,0,0,0,80,0,29,0,214,0,54,0,129,0,207,0,79,0,132,0,205,0,241,0,211,0,0,0,13,0,212,0,152,0,210,0,0,0,104,0,0,0,0,0,0,0,0,0,201,0,235,0,19,0,208,0,109,0,0,0,12,0,32,0,74,0,91,0,178,0,164,0,24,0,0,0,213,0,66,0,194,0,0,0,147,0,34,0,33,0,0,0,141,0,31,0,89,0,24,0,141,0,129,0,73,0,179,0,0,0,80,0,132,0,208,0,125,0,18,0,237,0,148,0,187,0,22,0,217,0,186,0,114,0,144,0,88,0,81,0,95,0,86,0,215,0,222,0,0,0,156,0,0,0,58,0,77,0,106,0,62,0,146,0,21,0,144,0,5,0,124,0,146,0,121,0,190,0,152,0,0,0,64,0,193,0,90,0,203,0,233,0,0,0,185,0,56,0,141,0,120,0,164,0,247,0,8,0,112,0,150,0,216,0,102,0,170,0,135,0,0,0,0,0,0,0,187,0,246,0,61,0,169,0,163,0,72,0,8,0,100,0,129,0,218,0,188,0,22,0,35,0,46,0,205,0,134,0,115,0,209,0,198,0,57,0,123,0,249,0,0,0,155,0,0,0,0,0,110,0,0,0,91,0,239,0,44,0,41,0,230,0,183,0,73,0,53,0,132,0,158,0,219,0,69,0,125,0,24,0,207,0,185,0,212,0,218,0,186,0,152,0,0,0,201,0,196,0,59,0,0,0,0,0,18,0,0,0,172,0,5,0,100,0,217,0,4,0,252,0,0,0,145,0,146,0,48,0,35,0,223,0,168,0,250,0,0,0,162,0,181,0,154,0,174,0,0,0,192,0,195,0,0,0,206,0,0,0,0,0,187,0,239,0,226,0,0,0,100,0,0,0,195,0,167,0,69,0,22,0,232,0,0,0,210,0,137,0,227,0,84,0,174,0,68,0,148,0,0,0,136,0,236,0,82,0,162,0,57,0,125,0,0,0,54,0,82,0,0,0,245,0,83,0,96,0,234,0,36,0,149,0,92,0,135,0,129,0,137,0,153,0,248,0,0,0,56,0,193,0,119,0,102,0,0,0,207,0,180,0,0,0,52,0,106,0,110,0,56,0,190,0,240,0,108,0,0,0,198,0,90,0,130,0,0,0,122,0,135,0,0,0,0,0,85,0,0,0,0,0,17,0,253,0,77,0,53,0,150,0,91,0,0,0,65,0,175,0,223,0,0,0,248,0,198,0,206,0,33,0,0,0,54,0,101,0,139,0,51,0,2,0,26,0,229,0,136,0,200,0,0,0,109,0,200,0,0,0,237,0,179,0,202,0,2,0,0,0,224,0,230,0,65,0,98,0,110,0,100,0,0,0,0,0,0,0,235,0,8,0,0,0,7,0,61,0,98,0,77,0,66,0,157,0,0,0,6,0,0,0,93,0,86,0,158,0,201,0,15,0,31,0,155,0,98,0,114,0,170,0,0,0,196,0,92,0,193,0,120,0,126,0,24,0,12,0,0,0,42,0,163,0,104,0,120,0,27,0,0,0,29,0,177,0,0,0,255,0,0,0,176,0,173,0,189,0,175,0,8,0,226,0,0,0,239,0,0,0,112,0,80,0,222,0,4,0,0,0,90,0,70,0,179,0,0,0,87,0,1,0,73,0,184,0,35,0,58,0,0,0,159,0,234,0,61,0,241,0,137,0,119,0,38,0,0,0,125,0,0,0,27,0,142,0,5,0,87,0,133,0,184,0,17,0,111,0,32,0,99,0,227,0,233,0,90,0,134,0,0,0,0,0,0,0,5,0,190,0,86,0,86,0,106,0,159,0,18,0,21,0,0,0,141,0,0,0,195,0,249,0,70,0,127,0,197,0,17,0,0,0,160,0,140,0,33,0,0,0,26,0,107,0,70,0,22,0,147,0,185,0,29,0,253,0,21,0,156,0,32,0,143,0,235,0,0,0,240,0,168,0,8,0,212,0,212,0,0,0,59,0,131,0,0,0,91,0,235,0,0,0,36,0,25,0,94,0,155,0,157,0,0,0,133,0,213,0,140,0,0,0,10,0,229,0,1,0,0,0,71,0,200,0,46,0,179,0,179,0,115,0,7,0,240,0,147,0,196,0,94,0,55,0,182,0,6,0,0,0,43,0,53,0,155,0,98,0,218,0,27,0,230,0,49,0,119,0,66,0,0,0,0,0,0,0,116,0,113,0,97,0,21,0,245,0,253,0,94,0,116,0,125,0,16,0,206,0,171,0,177,0,250,0,30,0,214,0,154,0,114,0,66,0,0,0,76,0,134,0,0,0,197,0,40,0,233,0,0,0,21,0,0,0,16,0,202,0,95,0,245,0,209,0,0,0,0,0,20,0,52,0,62,0,51,0,89,0,169,0,0,0,153,0,39,0,1,0,179,0,0,0,50,0,119,0,195,0,57,0,131,0,44,0,237,0,222,0,116,0,0,0,0,0,0,0,0,0,240,0,104,0,8,0,101,0,168,0,0,0,36,0,0,0,60,0,20,0,40,0,35,0,125,0,90,0,0,0,105,0,112,0,156,0,109,0,225,0,84,0,179,0,0,0,59,0,0,0,0,0,6,0,198,0,122,0,183,0,53,0,230,0,23,0,247,0,32,0,0,0,53,0,240,0,0,0,230,0,227,0,164,0,197,0,179,0,0,0,97,0,171,0,173,0,23,0,219,0,137,0,116,0,13,0,236,0,251,0,184,0,73,0,0,0,36,0,224,0,108,0,155,0,67,0,44,0,126,0,211,0,41,0,169,0,128,0,175,0,238,0,154,0,148,0,0,0,231,0,235,0,0,0,15,0,0,0,10,0,171,0,0,0,170,0,68,0,74,0,37,0,185,0,181,0,0,0,0,0,145,0,196,0,189,0,163,0,107,0,77,0,153,0,112,0,0,0,110,0,38,0,154,0,0,0,204,0,155,0,114,0,19,0,46,0,79,0,0,0,92,0,41,0,91,0,0,0,234,0,56,0,227,0,0,0,0,0,155,0,105,0,118,0,142,0,163,0,39,0,134,0,43,0,95,0,0,0,17,0,0,0,70,0,116,0,61,0,0,0,177,0,230,0,48,0,245,0,201,0,202,0,42,0,0,0,227,0,0,0,0,0,0,0,157,0,129,0,244,0,0,0,209,0,153,0,195,0,248,0,149,0,200,0,101,0,67,0,46,0,101,0,31,0,60,0,171,0,0,0,119,0,126,0,21,0,0,0,28,0,43,0,66,0,0,0,24,0,189,0,178,0,137,0,72,0,0,0,71,0,66,0,157,0,4,0,46,0,0,0,221,0,238,0,225,0,169,0,130,0,232,0,26,0,164,0,0,0,132,0,195,0,199,0,0,0,73,0,68,0,246,0,162,0,126,0,0,0,197,0,45,0,0,0,0,0,0,0,191,0,0,0,168,0,0,0,234,0,80,0,235,0,36,0,186,0,0,0,0,0,127,0,60,0,82,0,8,0,222,0,0,0,0,0,52,0,0,0,60,0,131,0,72,0,66,0,118,0,32,0,208,0,0,0,0,0,213,0,113,0,229,0,254,0,60,0,200,0,232,0,212,0,216,0,0,0,37,0,59,0,0,0,164,0,0,0,0,0,94,0,163,0,223,0,205,0,196,0,0,0,0,0,0,0,0,0,110,0,4,0,14,0,166,0,178,0,5,0,0,0,199,0,0,0,79,0,80,0,56,0,191,0,15,0,0,0,184,0,187,0,126,0,121,0,31,0,70,0,148,0,0,0,194,0,149,0,218,0,150,0,118,0,240,0,218,0,189,0,42,0,45,0,126,0,11,0,175,0,206,0,246,0,35,0,73,0,1,0,155,0,202,0,195,0,136,0,0,0,44,0,232,0);
signal scenario_full  : scenario_type := (207,31,220,31,220,30,220,29,61,31,27,31,26,31,125,31,56,31,56,30,101,31,175,31,194,31,191,31,32,31,51,31,165,31,142,31,142,30,47,31,143,31,147,31,5,31,139,31,239,31,43,31,113,31,253,31,253,30,177,31,25,31,25,30,25,29,55,31,216,31,122,31,152,31,142,31,149,31,136,31,24,31,158,31,158,30,117,31,253,31,253,30,253,29,23,31,219,31,56,31,41,31,41,30,132,31,42,31,85,31,151,31,145,31,5,31,30,31,45,31,45,30,180,31,210,31,129,31,135,31,44,31,76,31,151,31,23,31,108,31,104,31,40,31,218,31,193,31,193,30,193,29,72,31,63,31,79,31,209,31,136,31,136,30,213,31,114,31,254,31,254,30,162,31,128,31,177,31,133,31,215,31,23,31,190,31,239,31,14,31,160,31,86,31,214,31,33,31,124,31,61,31,61,30,214,31,214,30,155,31,155,30,16,31,20,31,20,31,20,31,191,31,191,30,191,29,80,31,29,31,214,31,54,31,129,31,207,31,79,31,132,31,205,31,241,31,211,31,211,30,13,31,212,31,152,31,210,31,210,30,104,31,104,30,104,29,104,28,104,27,201,31,235,31,19,31,208,31,109,31,109,30,12,31,32,31,74,31,91,31,178,31,164,31,24,31,24,30,213,31,66,31,194,31,194,30,147,31,34,31,33,31,33,30,141,31,31,31,89,31,24,31,141,31,129,31,73,31,179,31,179,30,80,31,132,31,208,31,125,31,18,31,237,31,148,31,187,31,22,31,217,31,186,31,114,31,144,31,88,31,81,31,95,31,86,31,215,31,222,31,222,30,156,31,156,30,58,31,77,31,106,31,62,31,146,31,21,31,144,31,5,31,124,31,146,31,121,31,190,31,152,31,152,30,64,31,193,31,90,31,203,31,233,31,233,30,185,31,56,31,141,31,120,31,164,31,247,31,8,31,112,31,150,31,216,31,102,31,170,31,135,31,135,30,135,29,135,28,187,31,246,31,61,31,169,31,163,31,72,31,8,31,100,31,129,31,218,31,188,31,22,31,35,31,46,31,205,31,134,31,115,31,209,31,198,31,57,31,123,31,249,31,249,30,155,31,155,30,155,29,110,31,110,30,91,31,239,31,44,31,41,31,230,31,183,31,73,31,53,31,132,31,158,31,219,31,69,31,125,31,24,31,207,31,185,31,212,31,218,31,186,31,152,31,152,30,201,31,196,31,59,31,59,30,59,29,18,31,18,30,172,31,5,31,100,31,217,31,4,31,252,31,252,30,145,31,146,31,48,31,35,31,223,31,168,31,250,31,250,30,162,31,181,31,154,31,174,31,174,30,192,31,195,31,195,30,206,31,206,30,206,29,187,31,239,31,226,31,226,30,100,31,100,30,195,31,167,31,69,31,22,31,232,31,232,30,210,31,137,31,227,31,84,31,174,31,68,31,148,31,148,30,136,31,236,31,82,31,162,31,57,31,125,31,125,30,54,31,82,31,82,30,245,31,83,31,96,31,234,31,36,31,149,31,92,31,135,31,129,31,137,31,153,31,248,31,248,30,56,31,193,31,119,31,102,31,102,30,207,31,180,31,180,30,52,31,106,31,110,31,56,31,190,31,240,31,108,31,108,30,198,31,90,31,130,31,130,30,122,31,135,31,135,30,135,29,85,31,85,30,85,29,17,31,253,31,77,31,53,31,150,31,91,31,91,30,65,31,175,31,223,31,223,30,248,31,198,31,206,31,33,31,33,30,54,31,101,31,139,31,51,31,2,31,26,31,229,31,136,31,200,31,200,30,109,31,200,31,200,30,237,31,179,31,202,31,2,31,2,30,224,31,230,31,65,31,98,31,110,31,100,31,100,30,100,29,100,28,235,31,8,31,8,30,7,31,61,31,98,31,77,31,66,31,157,31,157,30,6,31,6,30,93,31,86,31,158,31,201,31,15,31,31,31,155,31,98,31,114,31,170,31,170,30,196,31,92,31,193,31,120,31,126,31,24,31,12,31,12,30,42,31,163,31,104,31,120,31,27,31,27,30,29,31,177,31,177,30,255,31,255,30,176,31,173,31,189,31,175,31,8,31,226,31,226,30,239,31,239,30,112,31,80,31,222,31,4,31,4,30,90,31,70,31,179,31,179,30,87,31,1,31,73,31,184,31,35,31,58,31,58,30,159,31,234,31,61,31,241,31,137,31,119,31,38,31,38,30,125,31,125,30,27,31,142,31,5,31,87,31,133,31,184,31,17,31,111,31,32,31,99,31,227,31,233,31,90,31,134,31,134,30,134,29,134,28,5,31,190,31,86,31,86,31,106,31,159,31,18,31,21,31,21,30,141,31,141,30,195,31,249,31,70,31,127,31,197,31,17,31,17,30,160,31,140,31,33,31,33,30,26,31,107,31,70,31,22,31,147,31,185,31,29,31,253,31,21,31,156,31,32,31,143,31,235,31,235,30,240,31,168,31,8,31,212,31,212,31,212,30,59,31,131,31,131,30,91,31,235,31,235,30,36,31,25,31,94,31,155,31,157,31,157,30,133,31,213,31,140,31,140,30,10,31,229,31,1,31,1,30,71,31,200,31,46,31,179,31,179,31,115,31,7,31,240,31,147,31,196,31,94,31,55,31,182,31,6,31,6,30,43,31,53,31,155,31,98,31,218,31,27,31,230,31,49,31,119,31,66,31,66,30,66,29,66,28,116,31,113,31,97,31,21,31,245,31,253,31,94,31,116,31,125,31,16,31,206,31,171,31,177,31,250,31,30,31,214,31,154,31,114,31,66,31,66,30,76,31,134,31,134,30,197,31,40,31,233,31,233,30,21,31,21,30,16,31,202,31,95,31,245,31,209,31,209,30,209,29,20,31,52,31,62,31,51,31,89,31,169,31,169,30,153,31,39,31,1,31,179,31,179,30,50,31,119,31,195,31,57,31,131,31,44,31,237,31,222,31,116,31,116,30,116,29,116,28,116,27,240,31,104,31,8,31,101,31,168,31,168,30,36,31,36,30,60,31,20,31,40,31,35,31,125,31,90,31,90,30,105,31,112,31,156,31,109,31,225,31,84,31,179,31,179,30,59,31,59,30,59,29,6,31,198,31,122,31,183,31,53,31,230,31,23,31,247,31,32,31,32,30,53,31,240,31,240,30,230,31,227,31,164,31,197,31,179,31,179,30,97,31,171,31,173,31,23,31,219,31,137,31,116,31,13,31,236,31,251,31,184,31,73,31,73,30,36,31,224,31,108,31,155,31,67,31,44,31,126,31,211,31,41,31,169,31,128,31,175,31,238,31,154,31,148,31,148,30,231,31,235,31,235,30,15,31,15,30,10,31,171,31,171,30,170,31,68,31,74,31,37,31,185,31,181,31,181,30,181,29,145,31,196,31,189,31,163,31,107,31,77,31,153,31,112,31,112,30,110,31,38,31,154,31,154,30,204,31,155,31,114,31,19,31,46,31,79,31,79,30,92,31,41,31,91,31,91,30,234,31,56,31,227,31,227,30,227,29,155,31,105,31,118,31,142,31,163,31,39,31,134,31,43,31,95,31,95,30,17,31,17,30,70,31,116,31,61,31,61,30,177,31,230,31,48,31,245,31,201,31,202,31,42,31,42,30,227,31,227,30,227,29,227,28,157,31,129,31,244,31,244,30,209,31,153,31,195,31,248,31,149,31,200,31,101,31,67,31,46,31,101,31,31,31,60,31,171,31,171,30,119,31,126,31,21,31,21,30,28,31,43,31,66,31,66,30,24,31,189,31,178,31,137,31,72,31,72,30,71,31,66,31,157,31,4,31,46,31,46,30,221,31,238,31,225,31,169,31,130,31,232,31,26,31,164,31,164,30,132,31,195,31,199,31,199,30,73,31,68,31,246,31,162,31,126,31,126,30,197,31,45,31,45,30,45,29,45,28,191,31,191,30,168,31,168,30,234,31,80,31,235,31,36,31,186,31,186,30,186,29,127,31,60,31,82,31,8,31,222,31,222,30,222,29,52,31,52,30,60,31,131,31,72,31,66,31,118,31,32,31,208,31,208,30,208,29,213,31,113,31,229,31,254,31,60,31,200,31,232,31,212,31,216,31,216,30,37,31,59,31,59,30,164,31,164,30,164,29,94,31,163,31,223,31,205,31,196,31,196,30,196,29,196,28,196,27,110,31,4,31,14,31,166,31,178,31,5,31,5,30,199,31,199,30,79,31,80,31,56,31,191,31,15,31,15,30,184,31,187,31,126,31,121,31,31,31,70,31,148,31,148,30,194,31,149,31,218,31,150,31,118,31,240,31,218,31,189,31,42,31,45,31,126,31,11,31,175,31,206,31,246,31,35,31,73,31,1,31,155,31,202,31,195,31,136,31,136,30,44,31,232,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
