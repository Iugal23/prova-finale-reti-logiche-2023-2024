-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 950;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,232,0,44,0,0,0,165,0,0,0,185,0,140,0,96,0,101,0,0,0,196,0,67,0,14,0,123,0,0,0,0,0,0,0,218,0,237,0,170,0,0,0,78,0,214,0,221,0,59,0,219,0,226,0,104,0,165,0,163,0,173,0,185,0,68,0,95,0,132,0,201,0,109,0,123,0,46,0,83,0,0,0,80,0,211,0,48,0,232,0,151,0,1,0,19,0,109,0,34,0,162,0,45,0,0,0,40,0,0,0,0,0,161,0,23,0,137,0,98,0,129,0,161,0,67,0,52,0,47,0,106,0,204,0,225,0,195,0,147,0,238,0,12,0,0,0,35,0,0,0,99,0,246,0,97,0,204,0,129,0,126,0,168,0,109,0,0,0,16,0,215,0,158,0,157,0,166,0,22,0,247,0,161,0,24,0,151,0,236,0,204,0,21,0,159,0,83,0,235,0,155,0,0,0,229,0,216,0,238,0,104,0,11,0,94,0,188,0,196,0,153,0,161,0,13,0,2,0,57,0,0,0,144,0,0,0,0,0,0,0,191,0,248,0,33,0,116,0,123,0,228,0,94,0,0,0,0,0,131,0,217,0,136,0,91,0,158,0,117,0,105,0,0,0,11,0,206,0,0,0,49,0,79,0,153,0,0,0,210,0,112,0,237,0,76,0,204,0,0,0,109,0,77,0,67,0,0,0,82,0,28,0,18,0,135,0,36,0,74,0,148,0,0,0,95,0,232,0,211,0,102,0,96,0,84,0,0,0,188,0,0,0,0,0,192,0,122,0,63,0,69,0,100,0,187,0,186,0,203,0,239,0,50,0,104,0,0,0,246,0,10,0,135,0,78,0,64,0,183,0,0,0,60,0,145,0,185,0,194,0,0,0,240,0,0,0,0,0,203,0,94,0,220,0,76,0,0,0,160,0,0,0,44,0,233,0,0,0,0,0,191,0,12,0,177,0,0,0,172,0,230,0,82,0,204,0,240,0,92,0,221,0,220,0,80,0,133,0,166,0,191,0,180,0,46,0,67,0,170,0,48,0,216,0,0,0,150,0,12,0,234,0,204,0,25,0,195,0,219,0,0,0,82,0,6,0,102,0,0,0,35,0,90,0,127,0,197,0,163,0,106,0,0,0,112,0,183,0,95,0,253,0,63,0,241,0,16,0,123,0,36,0,197,0,235,0,161,0,101,0,111,0,204,0,80,0,248,0,224,0,105,0,79,0,226,0,103,0,218,0,176,0,109,0,0,0,37,0,0,0,8,0,150,0,198,0,211,0,144,0,54,0,132,0,0,0,57,0,254,0,233,0,0,0,0,0,41,0,40,0,112,0,53,0,221,0,34,0,93,0,0,0,137,0,164,0,0,0,74,0,181,0,111,0,176,0,222,0,19,0,245,0,210,0,8,0,173,0,27,0,156,0,188,0,0,0,0,0,156,0,208,0,21,0,124,0,13,0,243,0,164,0,136,0,72,0,236,0,83,0,29,0,94,0,20,0,213,0,245,0,121,0,210,0,228,0,0,0,187,0,51,0,0,0,0,0,212,0,0,0,239,0,52,0,0,0,11,0,0,0,0,0,0,0,39,0,65,0,0,0,246,0,22,0,224,0,244,0,162,0,0,0,78,0,103,0,0,0,0,0,193,0,63,0,95,0,138,0,9,0,161,0,0,0,210,0,96,0,0,0,99,0,21,0,197,0,73,0,63,0,171,0,242,0,0,0,0,0,0,0,212,0,205,0,0,0,36,0,22,0,214,0,63,0,75,0,55,0,237,0,117,0,141,0,195,0,52,0,241,0,244,0,225,0,210,0,196,0,0,0,0,0,83,0,36,0,174,0,38,0,52,0,242,0,70,0,0,0,180,0,0,0,206,0,0,0,59,0,144,0,0,0,172,0,155,0,245,0,0,0,0,0,57,0,125,0,44,0,78,0,146,0,235,0,0,0,79,0,122,0,200,0,255,0,115,0,183,0,119,0,175,0,251,0,0,0,0,0,184,0,106,0,140,0,100,0,214,0,58,0,0,0,0,0,198,0,216,0,133,0,85,0,201,0,80,0,110,0,164,0,172,0,150,0,252,0,211,0,208,0,0,0,0,0,57,0,94,0,181,0,170,0,118,0,202,0,111,0,154,0,124,0,0,0,29,0,0,0,0,0,192,0,229,0,86,0,71,0,159,0,106,0,149,0,0,0,239,0,0,0,0,0,61,0,163,0,236,0,192,0,117,0,177,0,241,0,0,0,242,0,21,0,216,0,183,0,142,0,230,0,170,0,178,0,160,0,199,0,111,0,148,0,78,0,220,0,38,0,5,0,202,0,28,0,79,0,0,0,0,0,64,0,50,0,96,0,0,0,52,0,150,0,255,0,56,0,200,0,252,0,119,0,55,0,0,0,0,0,0,0,230,0,1,0,204,0,115,0,153,0,3,0,85,0,0,0,0,0,54,0,125,0,159,0,135,0,118,0,196,0,78,0,248,0,146,0,72,0,0,0,251,0,81,0,0,0,33,0,0,0,128,0,92,0,127,0,0,0,63,0,174,0,0,0,0,0,133,0,47,0,86,0,191,0,179,0,41,0,0,0,125,0,0,0,59,0,211,0,0,0,89,0,130,0,184,0,0,0,95,0,0,0,138,0,0,0,0,0,0,0,224,0,52,0,23,0,181,0,181,0,164,0,0,0,186,0,236,0,136,0,133,0,53,0,124,0,9,0,203,0,143,0,35,0,70,0,97,0,0,0,60,0,0,0,0,0,44,0,1,0,167,0,0,0,200,0,189,0,136,0,237,0,140,0,11,0,0,0,38,0,140,0,31,0,183,0,198,0,102,0,31,0,0,0,153,0,101,0,112,0,235,0,181,0,50,0,40,0,0,0,0,0,14,0,108,0,96,0,0,0,150,0,81,0,4,0,12,0,209,0,39,0,0,0,45,0,26,0,80,0,128,0,0,0,253,0,203,0,0,0,21,0,0,0,142,0,81,0,144,0,140,0,161,0,0,0,128,0,104,0,109,0,175,0,0,0,114,0,77,0,148,0,165,0,176,0,22,0,188,0,0,0,198,0,202,0,186,0,26,0,0,0,132,0,0,0,164,0,145,0,176,0,1,0,195,0,0,0,0,0,146,0,101,0,143,0,149,0,216,0,162,0,1,0,76,0,233,0,190,0,241,0,9,0,0,0,78,0,58,0,67,0,245,0,0,0,0,0,95,0,62,0,182,0,235,0,0,0,95,0,255,0,145,0,50,0,253,0,1,0,30,0,101,0,204,0,87,0,185,0,192,0,240,0,0,0,0,0,0,0,201,0,0,0,222,0,0,0,160,0,140,0,197,0,122,0,171,0,90,0,48,0,35,0,179,0,232,0,156,0,0,0,78,0,203,0,151,0,0,0,182,0,0,0,0,0,251,0,27,0,0,0,195,0,10,0,70,0,184,0,0,0,136,0,63,0,191,0,27,0,210,0,26,0,22,0,198,0,13,0,162,0,250,0,142,0,144,0,0,0,96,0,92,0,141,0,52,0,0,0,225,0,92,0,0,0,180,0,0,0,0,0,6,0,199,0,16,0,97,0,215,0,164,0,62,0,134,0,93,0,157,0,24,0,162,0,148,0,219,0,0,0,0,0,224,0,0,0,190,0,0,0,0,0,0,0,29,0,156,0,0,0,8,0,253,0,225,0,3,0,0,0,102,0,149,0,38,0,191,0,239,0,95,0,0,0,137,0,7,0,217,0,117,0,0,0,122,0,53,0,237,0,172,0,165,0,0,0,128,0,227,0,0,0,147,0,171,0,0,0,0,0,144,0,175,0,106,0,118,0,186,0,0,0,152,0,17,0,219,0,2,0,0,0,249,0,233,0,164,0,140,0,47,0,0,0,234,0,254,0,0,0,19,0,0,0,80,0,0,0,124,0,74,0,176,0,253,0,222,0,158,0,97,0,219,0,184,0,250,0,55,0,111,0,0,0,102,0,0,0,223,0,2,0,9,0,0,0,115,0,150,0,0,0,202,0,0,0,169,0,67,0,50,0,201,0,186,0,182,0,105,0,199,0,111,0,135,0,64,0,191,0,96,0,58,0,230,0,0,0,212,0,84,0,39,0,243,0,0,0,112,0,213,0,115,0,56,0,0,0,11,0,196,0,42,0,91,0,137,0,68,0,232,0,157,0,196,0,0,0,222,0,131,0,160,0,1,0,37,0,105,0,1,0,0,0,160,0,0,0,121,0,85,0,239,0,208,0,76,0,240,0,73,0,0,0,95,0);
signal scenario_full  : scenario_type := (0,0,232,31,44,31,44,30,165,31,165,30,185,31,140,31,96,31,101,31,101,30,196,31,67,31,14,31,123,31,123,30,123,29,123,28,218,31,237,31,170,31,170,30,78,31,214,31,221,31,59,31,219,31,226,31,104,31,165,31,163,31,173,31,185,31,68,31,95,31,132,31,201,31,109,31,123,31,46,31,83,31,83,30,80,31,211,31,48,31,232,31,151,31,1,31,19,31,109,31,34,31,162,31,45,31,45,30,40,31,40,30,40,29,161,31,23,31,137,31,98,31,129,31,161,31,67,31,52,31,47,31,106,31,204,31,225,31,195,31,147,31,238,31,12,31,12,30,35,31,35,30,99,31,246,31,97,31,204,31,129,31,126,31,168,31,109,31,109,30,16,31,215,31,158,31,157,31,166,31,22,31,247,31,161,31,24,31,151,31,236,31,204,31,21,31,159,31,83,31,235,31,155,31,155,30,229,31,216,31,238,31,104,31,11,31,94,31,188,31,196,31,153,31,161,31,13,31,2,31,57,31,57,30,144,31,144,30,144,29,144,28,191,31,248,31,33,31,116,31,123,31,228,31,94,31,94,30,94,29,131,31,217,31,136,31,91,31,158,31,117,31,105,31,105,30,11,31,206,31,206,30,49,31,79,31,153,31,153,30,210,31,112,31,237,31,76,31,204,31,204,30,109,31,77,31,67,31,67,30,82,31,28,31,18,31,135,31,36,31,74,31,148,31,148,30,95,31,232,31,211,31,102,31,96,31,84,31,84,30,188,31,188,30,188,29,192,31,122,31,63,31,69,31,100,31,187,31,186,31,203,31,239,31,50,31,104,31,104,30,246,31,10,31,135,31,78,31,64,31,183,31,183,30,60,31,145,31,185,31,194,31,194,30,240,31,240,30,240,29,203,31,94,31,220,31,76,31,76,30,160,31,160,30,44,31,233,31,233,30,233,29,191,31,12,31,177,31,177,30,172,31,230,31,82,31,204,31,240,31,92,31,221,31,220,31,80,31,133,31,166,31,191,31,180,31,46,31,67,31,170,31,48,31,216,31,216,30,150,31,12,31,234,31,204,31,25,31,195,31,219,31,219,30,82,31,6,31,102,31,102,30,35,31,90,31,127,31,197,31,163,31,106,31,106,30,112,31,183,31,95,31,253,31,63,31,241,31,16,31,123,31,36,31,197,31,235,31,161,31,101,31,111,31,204,31,80,31,248,31,224,31,105,31,79,31,226,31,103,31,218,31,176,31,109,31,109,30,37,31,37,30,8,31,150,31,198,31,211,31,144,31,54,31,132,31,132,30,57,31,254,31,233,31,233,30,233,29,41,31,40,31,112,31,53,31,221,31,34,31,93,31,93,30,137,31,164,31,164,30,74,31,181,31,111,31,176,31,222,31,19,31,245,31,210,31,8,31,173,31,27,31,156,31,188,31,188,30,188,29,156,31,208,31,21,31,124,31,13,31,243,31,164,31,136,31,72,31,236,31,83,31,29,31,94,31,20,31,213,31,245,31,121,31,210,31,228,31,228,30,187,31,51,31,51,30,51,29,212,31,212,30,239,31,52,31,52,30,11,31,11,30,11,29,11,28,39,31,65,31,65,30,246,31,22,31,224,31,244,31,162,31,162,30,78,31,103,31,103,30,103,29,193,31,63,31,95,31,138,31,9,31,161,31,161,30,210,31,96,31,96,30,99,31,21,31,197,31,73,31,63,31,171,31,242,31,242,30,242,29,242,28,212,31,205,31,205,30,36,31,22,31,214,31,63,31,75,31,55,31,237,31,117,31,141,31,195,31,52,31,241,31,244,31,225,31,210,31,196,31,196,30,196,29,83,31,36,31,174,31,38,31,52,31,242,31,70,31,70,30,180,31,180,30,206,31,206,30,59,31,144,31,144,30,172,31,155,31,245,31,245,30,245,29,57,31,125,31,44,31,78,31,146,31,235,31,235,30,79,31,122,31,200,31,255,31,115,31,183,31,119,31,175,31,251,31,251,30,251,29,184,31,106,31,140,31,100,31,214,31,58,31,58,30,58,29,198,31,216,31,133,31,85,31,201,31,80,31,110,31,164,31,172,31,150,31,252,31,211,31,208,31,208,30,208,29,57,31,94,31,181,31,170,31,118,31,202,31,111,31,154,31,124,31,124,30,29,31,29,30,29,29,192,31,229,31,86,31,71,31,159,31,106,31,149,31,149,30,239,31,239,30,239,29,61,31,163,31,236,31,192,31,117,31,177,31,241,31,241,30,242,31,21,31,216,31,183,31,142,31,230,31,170,31,178,31,160,31,199,31,111,31,148,31,78,31,220,31,38,31,5,31,202,31,28,31,79,31,79,30,79,29,64,31,50,31,96,31,96,30,52,31,150,31,255,31,56,31,200,31,252,31,119,31,55,31,55,30,55,29,55,28,230,31,1,31,204,31,115,31,153,31,3,31,85,31,85,30,85,29,54,31,125,31,159,31,135,31,118,31,196,31,78,31,248,31,146,31,72,31,72,30,251,31,81,31,81,30,33,31,33,30,128,31,92,31,127,31,127,30,63,31,174,31,174,30,174,29,133,31,47,31,86,31,191,31,179,31,41,31,41,30,125,31,125,30,59,31,211,31,211,30,89,31,130,31,184,31,184,30,95,31,95,30,138,31,138,30,138,29,138,28,224,31,52,31,23,31,181,31,181,31,164,31,164,30,186,31,236,31,136,31,133,31,53,31,124,31,9,31,203,31,143,31,35,31,70,31,97,31,97,30,60,31,60,30,60,29,44,31,1,31,167,31,167,30,200,31,189,31,136,31,237,31,140,31,11,31,11,30,38,31,140,31,31,31,183,31,198,31,102,31,31,31,31,30,153,31,101,31,112,31,235,31,181,31,50,31,40,31,40,30,40,29,14,31,108,31,96,31,96,30,150,31,81,31,4,31,12,31,209,31,39,31,39,30,45,31,26,31,80,31,128,31,128,30,253,31,203,31,203,30,21,31,21,30,142,31,81,31,144,31,140,31,161,31,161,30,128,31,104,31,109,31,175,31,175,30,114,31,77,31,148,31,165,31,176,31,22,31,188,31,188,30,198,31,202,31,186,31,26,31,26,30,132,31,132,30,164,31,145,31,176,31,1,31,195,31,195,30,195,29,146,31,101,31,143,31,149,31,216,31,162,31,1,31,76,31,233,31,190,31,241,31,9,31,9,30,78,31,58,31,67,31,245,31,245,30,245,29,95,31,62,31,182,31,235,31,235,30,95,31,255,31,145,31,50,31,253,31,1,31,30,31,101,31,204,31,87,31,185,31,192,31,240,31,240,30,240,29,240,28,201,31,201,30,222,31,222,30,160,31,140,31,197,31,122,31,171,31,90,31,48,31,35,31,179,31,232,31,156,31,156,30,78,31,203,31,151,31,151,30,182,31,182,30,182,29,251,31,27,31,27,30,195,31,10,31,70,31,184,31,184,30,136,31,63,31,191,31,27,31,210,31,26,31,22,31,198,31,13,31,162,31,250,31,142,31,144,31,144,30,96,31,92,31,141,31,52,31,52,30,225,31,92,31,92,30,180,31,180,30,180,29,6,31,199,31,16,31,97,31,215,31,164,31,62,31,134,31,93,31,157,31,24,31,162,31,148,31,219,31,219,30,219,29,224,31,224,30,190,31,190,30,190,29,190,28,29,31,156,31,156,30,8,31,253,31,225,31,3,31,3,30,102,31,149,31,38,31,191,31,239,31,95,31,95,30,137,31,7,31,217,31,117,31,117,30,122,31,53,31,237,31,172,31,165,31,165,30,128,31,227,31,227,30,147,31,171,31,171,30,171,29,144,31,175,31,106,31,118,31,186,31,186,30,152,31,17,31,219,31,2,31,2,30,249,31,233,31,164,31,140,31,47,31,47,30,234,31,254,31,254,30,19,31,19,30,80,31,80,30,124,31,74,31,176,31,253,31,222,31,158,31,97,31,219,31,184,31,250,31,55,31,111,31,111,30,102,31,102,30,223,31,2,31,9,31,9,30,115,31,150,31,150,30,202,31,202,30,169,31,67,31,50,31,201,31,186,31,182,31,105,31,199,31,111,31,135,31,64,31,191,31,96,31,58,31,230,31,230,30,212,31,84,31,39,31,243,31,243,30,112,31,213,31,115,31,56,31,56,30,11,31,196,31,42,31,91,31,137,31,68,31,232,31,157,31,196,31,196,30,222,31,131,31,160,31,1,31,37,31,105,31,1,31,1,30,160,31,160,30,121,31,85,31,239,31,208,31,76,31,240,31,73,31,73,30,95,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
