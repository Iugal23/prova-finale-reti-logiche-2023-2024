-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 239;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (154,0,237,0,48,0,172,0,0,0,0,0,86,0,222,0,19,0,67,0,119,0,0,0,30,0,0,0,173,0,142,0,184,0,192,0,168,0,199,0,77,0,20,0,0,0,85,0,156,0,154,0,48,0,0,0,24,0,4,0,107,0,229,0,0,0,32,0,0,0,135,0,112,0,159,0,248,0,134,0,182,0,69,0,95,0,155,0,18,0,0,0,110,0,0,0,129,0,95,0,87,0,11,0,202,0,36,0,1,0,0,0,74,0,128,0,133,0,45,0,184,0,0,0,160,0,45,0,0,0,56,0,0,0,0,0,84,0,69,0,25,0,5,0,34,0,113,0,174,0,161,0,0,0,146,0,90,0,235,0,133,0,0,0,79,0,58,0,179,0,211,0,127,0,0,0,0,0,95,0,177,0,0,0,158,0,0,0,158,0,223,0,136,0,0,0,113,0,0,0,51,0,0,0,0,0,116,0,152,0,73,0,51,0,42,0,70,0,225,0,106,0,45,0,178,0,0,0,194,0,137,0,9,0,106,0,222,0,0,0,0,0,84,0,183,0,42,0,95,0,116,0,16,0,87,0,240,0,0,0,237,0,220,0,114,0,48,0,254,0,144,0,20,0,154,0,85,0,0,0,6,0,177,0,76,0,3,0,146,0,0,0,67,0,227,0,248,0,49,0,130,0,21,0,51,0,50,0,0,0,200,0,0,0,77,0,42,0,20,0,176,0,137,0,5,0,234,0,0,0,28,0,0,0,75,0,237,0,0,0,0,0,57,0,113,0,169,0,0,0,153,0,189,0,194,0,115,0,158,0,139,0,148,0,111,0,212,0,38,0,190,0,191,0,49,0,0,0,178,0,0,0,51,0,223,0,0,0,78,0,88,0,8,0,0,0,137,0,236,0,150,0,115,0,253,0,159,0,0,0,0,0,210,0,149,0,213,0,184,0,184,0,180,0,23,0,0,0,117,0,251,0,93,0,252,0,225,0,55,0,172,0,12,0,122,0,197,0,0,0,0,0,57,0,186,0,241,0,186,0,0,0,29,0,161,0,203,0,0,0,0,0,246,0,22,0,0,0);
signal scenario_full  : scenario_type := (154,31,237,31,48,31,172,31,172,30,172,29,86,31,222,31,19,31,67,31,119,31,119,30,30,31,30,30,173,31,142,31,184,31,192,31,168,31,199,31,77,31,20,31,20,30,85,31,156,31,154,31,48,31,48,30,24,31,4,31,107,31,229,31,229,30,32,31,32,30,135,31,112,31,159,31,248,31,134,31,182,31,69,31,95,31,155,31,18,31,18,30,110,31,110,30,129,31,95,31,87,31,11,31,202,31,36,31,1,31,1,30,74,31,128,31,133,31,45,31,184,31,184,30,160,31,45,31,45,30,56,31,56,30,56,29,84,31,69,31,25,31,5,31,34,31,113,31,174,31,161,31,161,30,146,31,90,31,235,31,133,31,133,30,79,31,58,31,179,31,211,31,127,31,127,30,127,29,95,31,177,31,177,30,158,31,158,30,158,31,223,31,136,31,136,30,113,31,113,30,51,31,51,30,51,29,116,31,152,31,73,31,51,31,42,31,70,31,225,31,106,31,45,31,178,31,178,30,194,31,137,31,9,31,106,31,222,31,222,30,222,29,84,31,183,31,42,31,95,31,116,31,16,31,87,31,240,31,240,30,237,31,220,31,114,31,48,31,254,31,144,31,20,31,154,31,85,31,85,30,6,31,177,31,76,31,3,31,146,31,146,30,67,31,227,31,248,31,49,31,130,31,21,31,51,31,50,31,50,30,200,31,200,30,77,31,42,31,20,31,176,31,137,31,5,31,234,31,234,30,28,31,28,30,75,31,237,31,237,30,237,29,57,31,113,31,169,31,169,30,153,31,189,31,194,31,115,31,158,31,139,31,148,31,111,31,212,31,38,31,190,31,191,31,49,31,49,30,178,31,178,30,51,31,223,31,223,30,78,31,88,31,8,31,8,30,137,31,236,31,150,31,115,31,253,31,159,31,159,30,159,29,210,31,149,31,213,31,184,31,184,31,180,31,23,31,23,30,117,31,251,31,93,31,252,31,225,31,55,31,172,31,12,31,122,31,197,31,197,30,197,29,57,31,186,31,241,31,186,31,186,30,29,31,161,31,203,31,203,30,203,29,246,31,22,31,22,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
