-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 335;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,226,0,86,0,105,0,117,0,0,0,0,0,0,0,218,0,225,0,0,0,53,0,185,0,114,0,35,0,206,0,0,0,229,0,77,0,16,0,81,0,0,0,42,0,184,0,0,0,212,0,234,0,198,0,53,0,236,0,179,0,224,0,237,0,0,0,189,0,223,0,99,0,201,0,142,0,233,0,20,0,252,0,210,0,0,0,183,0,75,0,27,0,118,0,133,0,232,0,0,0,81,0,252,0,0,0,153,0,191,0,132,0,223,0,65,0,68,0,214,0,0,0,118,0,159,0,0,0,44,0,152,0,0,0,159,0,38,0,179,0,63,0,145,0,151,0,0,0,5,0,59,0,111,0,106,0,110,0,157,0,213,0,152,0,68,0,184,0,5,0,0,0,88,0,157,0,19,0,22,0,105,0,0,0,0,0,67,0,125,0,0,0,0,0,71,0,0,0,76,0,76,0,49,0,161,0,0,0,26,0,180,0,0,0,136,0,194,0,0,0,168,0,135,0,0,0,145,0,23,0,1,0,207,0,113,0,0,0,131,0,33,0,207,0,184,0,61,0,0,0,0,0,211,0,227,0,0,0,46,0,0,0,60,0,7,0,0,0,131,0,0,0,248,0,53,0,96,0,0,0,0,0,172,0,230,0,213,0,16,0,235,0,102,0,152,0,103,0,57,0,86,0,0,0,246,0,51,0,196,0,0,0,0,0,251,0,75,0,86,0,125,0,183,0,55,0,0,0,186,0,0,0,180,0,27,0,78,0,154,0,72,0,251,0,135,0,205,0,135,0,252,0,168,0,115,0,124,0,44,0,191,0,132,0,0,0,241,0,89,0,98,0,149,0,197,0,254,0,27,0,130,0,108,0,155,0,146,0,196,0,0,0,46,0,139,0,196,0,185,0,186,0,0,0,155,0,110,0,74,0,205,0,132,0,96,0,191,0,19,0,171,0,119,0,111,0,158,0,234,0,237,0,40,0,76,0,37,0,197,0,237,0,159,0,0,0,24,0,216,0,58,0,230,0,140,0,93,0,0,0,250,0,0,0,146,0,148,0,244,0,0,0,35,0,36,0,242,0,79,0,87,0,212,0,233,0,184,0,128,0,194,0,0,0,0,0,60,0,106,0,247,0,161,0,160,0,183,0,197,0,52,0,30,0,17,0,0,0,163,0,61,0,192,0,17,0,115,0,71,0,0,0,144,0,233,0,0,0,28,0,25,0,157,0,24,0,40,0,253,0,22,0,136,0,47,0,0,0,0,0,40,0,133,0,38,0,239,0,2,0,239,0,38,0,238,0,218,0,141,0,143,0,55,0,69,0,79,0,119,0,4,0,0,0,58,0,172,0,0,0,224,0,0,0,203,0,49,0,27,0,9,0,0,0,251,0,126,0,67,0,149,0,0,0,0,0,130,0,37,0,194,0,2,0,149,0,215,0,188,0,36,0,82,0,57,0,51,0,0,0,3,0,206,0,121,0,108,0,181,0,6,0,229,0,58,0,234,0);
signal scenario_full  : scenario_type := (0,0,226,31,86,31,105,31,117,31,117,30,117,29,117,28,218,31,225,31,225,30,53,31,185,31,114,31,35,31,206,31,206,30,229,31,77,31,16,31,81,31,81,30,42,31,184,31,184,30,212,31,234,31,198,31,53,31,236,31,179,31,224,31,237,31,237,30,189,31,223,31,99,31,201,31,142,31,233,31,20,31,252,31,210,31,210,30,183,31,75,31,27,31,118,31,133,31,232,31,232,30,81,31,252,31,252,30,153,31,191,31,132,31,223,31,65,31,68,31,214,31,214,30,118,31,159,31,159,30,44,31,152,31,152,30,159,31,38,31,179,31,63,31,145,31,151,31,151,30,5,31,59,31,111,31,106,31,110,31,157,31,213,31,152,31,68,31,184,31,5,31,5,30,88,31,157,31,19,31,22,31,105,31,105,30,105,29,67,31,125,31,125,30,125,29,71,31,71,30,76,31,76,31,49,31,161,31,161,30,26,31,180,31,180,30,136,31,194,31,194,30,168,31,135,31,135,30,145,31,23,31,1,31,207,31,113,31,113,30,131,31,33,31,207,31,184,31,61,31,61,30,61,29,211,31,227,31,227,30,46,31,46,30,60,31,7,31,7,30,131,31,131,30,248,31,53,31,96,31,96,30,96,29,172,31,230,31,213,31,16,31,235,31,102,31,152,31,103,31,57,31,86,31,86,30,246,31,51,31,196,31,196,30,196,29,251,31,75,31,86,31,125,31,183,31,55,31,55,30,186,31,186,30,180,31,27,31,78,31,154,31,72,31,251,31,135,31,205,31,135,31,252,31,168,31,115,31,124,31,44,31,191,31,132,31,132,30,241,31,89,31,98,31,149,31,197,31,254,31,27,31,130,31,108,31,155,31,146,31,196,31,196,30,46,31,139,31,196,31,185,31,186,31,186,30,155,31,110,31,74,31,205,31,132,31,96,31,191,31,19,31,171,31,119,31,111,31,158,31,234,31,237,31,40,31,76,31,37,31,197,31,237,31,159,31,159,30,24,31,216,31,58,31,230,31,140,31,93,31,93,30,250,31,250,30,146,31,148,31,244,31,244,30,35,31,36,31,242,31,79,31,87,31,212,31,233,31,184,31,128,31,194,31,194,30,194,29,60,31,106,31,247,31,161,31,160,31,183,31,197,31,52,31,30,31,17,31,17,30,163,31,61,31,192,31,17,31,115,31,71,31,71,30,144,31,233,31,233,30,28,31,25,31,157,31,24,31,40,31,253,31,22,31,136,31,47,31,47,30,47,29,40,31,133,31,38,31,239,31,2,31,239,31,38,31,238,31,218,31,141,31,143,31,55,31,69,31,79,31,119,31,4,31,4,30,58,31,172,31,172,30,224,31,224,30,203,31,49,31,27,31,9,31,9,30,251,31,126,31,67,31,149,31,149,30,149,29,130,31,37,31,194,31,2,31,149,31,215,31,188,31,36,31,82,31,57,31,51,31,51,30,3,31,206,31,121,31,108,31,181,31,6,31,229,31,58,31,234,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
