-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 831;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (35,0,183,0,243,0,14,0,102,0,72,0,0,0,54,0,0,0,193,0,127,0,56,0,207,0,134,0,97,0,252,0,157,0,152,0,75,0,28,0,74,0,55,0,196,0,50,0,29,0,27,0,0,0,173,0,0,0,122,0,75,0,155,0,134,0,96,0,0,0,245,0,143,0,64,0,0,0,228,0,111,0,29,0,9,0,0,0,0,0,0,0,50,0,211,0,65,0,0,0,52,0,51,0,96,0,94,0,95,0,0,0,235,0,189,0,0,0,98,0,178,0,162,0,100,0,173,0,0,0,0,0,0,0,201,0,158,0,215,0,234,0,158,0,0,0,133,0,0,0,0,0,148,0,0,0,130,0,187,0,8,0,241,0,248,0,0,0,0,0,186,0,94,0,20,0,0,0,19,0,171,0,76,0,225,0,200,0,0,0,0,0,223,0,2,0,159,0,57,0,0,0,58,0,0,0,224,0,88,0,97,0,86,0,27,0,104,0,0,0,114,0,35,0,0,0,211,0,28,0,101,0,94,0,194,0,160,0,44,0,0,0,0,0,23,0,241,0,103,0,0,0,159,0,206,0,178,0,52,0,209,0,0,0,152,0,99,0,213,0,228,0,0,0,154,0,123,0,195,0,136,0,0,0,13,0,82,0,200,0,126,0,66,0,153,0,118,0,235,0,95,0,243,0,69,0,0,0,221,0,201,0,0,0,0,0,243,0,154,0,206,0,0,0,71,0,0,0,0,0,105,0,0,0,250,0,174,0,139,0,20,0,171,0,68,0,239,0,231,0,0,0,41,0,191,0,138,0,213,0,43,0,227,0,182,0,86,0,37,0,0,0,229,0,178,0,128,0,231,0,97,0,0,0,51,0,0,0,207,0,225,0,11,0,125,0,245,0,0,0,239,0,110,0,30,0,205,0,238,0,0,0,214,0,123,0,55,0,219,0,113,0,4,0,71,0,0,0,86,0,202,0,250,0,156,0,239,0,139,0,55,0,0,0,207,0,85,0,0,0,49,0,0,0,178,0,225,0,0,0,147,0,155,0,93,0,0,0,64,0,231,0,86,0,225,0,70,0,32,0,84,0,198,0,0,0,204,0,0,0,169,0,213,0,163,0,106,0,212,0,4,0,175,0,133,0,69,0,122,0,78,0,0,0,29,0,51,0,253,0,0,0,173,0,127,0,116,0,67,0,26,0,223,0,136,0,252,0,174,0,157,0,0,0,23,0,38,0,250,0,11,0,163,0,249,0,0,0,244,0,181,0,60,0,12,0,137,0,150,0,230,0,173,0,0,0,55,0,124,0,0,0,130,0,137,0,199,0,150,0,72,0,172,0,173,0,0,0,32,0,153,0,108,0,234,0,14,0,116,0,21,0,75,0,11,0,0,0,0,0,240,0,234,0,113,0,18,0,0,0,246,0,193,0,99,0,35,0,137,0,252,0,213,0,0,0,0,0,133,0,34,0,189,0,144,0,13,0,83,0,241,0,135,0,166,0,0,0,60,0,214,0,155,0,67,0,80,0,218,0,222,0,47,0,160,0,119,0,5,0,74,0,77,0,198,0,75,0,0,0,3,0,87,0,105,0,0,0,241,0,79,0,21,0,109,0,0,0,0,0,0,0,31,0,0,0,13,0,69,0,30,0,206,0,174,0,48,0,99,0,27,0,0,0,0,0,0,0,208,0,178,0,109,0,0,0,4,0,0,0,87,0,192,0,71,0,189,0,188,0,55,0,207,0,0,0,221,0,166,0,229,0,43,0,0,0,251,0,38,0,244,0,0,0,155,0,80,0,30,0,0,0,0,0,199,0,198,0,0,0,191,0,65,0,179,0,14,0,251,0,0,0,165,0,33,0,212,0,0,0,0,0,67,0,60,0,111,0,0,0,109,0,51,0,53,0,149,0,0,0,170,0,234,0,149,0,150,0,224,0,198,0,163,0,70,0,58,0,84,0,44,0,41,0,55,0,48,0,64,0,231,0,205,0,0,0,0,0,72,0,195,0,180,0,241,0,216,0,252,0,100,0,22,0,0,0,240,0,0,0,0,0,22,0,110,0,112,0,196,0,24,0,184,0,119,0,6,0,80,0,221,0,184,0,204,0,56,0,0,0,163,0,209,0,54,0,0,0,0,0,232,0,0,0,199,0,130,0,206,0,204,0,42,0,241,0,35,0,215,0,78,0,136,0,162,0,196,0,0,0,200,0,201,0,189,0,39,0,212,0,0,0,63,0,115,0,0,0,239,0,0,0,108,0,130,0,101,0,0,0,29,0,187,0,3,0,6,0,159,0,66,0,0,0,144,0,122,0,195,0,15,0,168,0,249,0,0,0,0,0,0,0,249,0,136,0,56,0,237,0,238,0,82,0,212,0,78,0,55,0,224,0,53,0,169,0,139,0,0,0,113,0,19,0,172,0,247,0,0,0,115,0,21,0,118,0,170,0,100,0,149,0,15,0,11,0,44,0,0,0,32,0,75,0,157,0,116,0,0,0,195,0,0,0,0,0,73,0,50,0,0,0,253,0,142,0,11,0,4,0,108,0,0,0,121,0,0,0,107,0,69,0,197,0,94,0,128,0,57,0,78,0,188,0,110,0,101,0,116,0,37,0,0,0,38,0,70,0,0,0,18,0,0,0,0,0,0,0,0,0,199,0,0,0,249,0,47,0,9,0,0,0,185,0,0,0,121,0,0,0,30,0,227,0,0,0,99,0,0,0,26,0,158,0,201,0,255,0,0,0,119,0,203,0,195,0,20,0,53,0,37,0,0,0,111,0,230,0,0,0,0,0,0,0,0,0,154,0,157,0,117,0,140,0,168,0,0,0,243,0,0,0,198,0,74,0,146,0,68,0,20,0,202,0,0,0,110,0,49,0,0,0,23,0,100,0,40,0,70,0,0,0,0,0,202,0,16,0,0,0,0,0,238,0,91,0,173,0,16,0,131,0,236,0,0,0,0,0,174,0,0,0,59,0,248,0,20,0,84,0,41,0,0,0,235,0,65,0,27,0,132,0,0,0,0,0,165,0,0,0,41,0,128,0,0,0,165,0,116,0,0,0,175,0,173,0,74,0,132,0,254,0,70,0,92,0,0,0,0,0,0,0,20,0,32,0,0,0,121,0,0,0,182,0,98,0,86,0,73,0,214,0,250,0,0,0,9,0,209,0,196,0,99,0,229,0,164,0,0,0,0,0,184,0,105,0,64,0,154,0,65,0,0,0,233,0,24,0,170,0,99,0,130,0,0,0,240,0,36,0,0,0,166,0,0,0,17,0,226,0,234,0,104,0,237,0,38,0,165,0,150,0,107,0,138,0,0,0,23,0,168,0,34,0,0,0,153,0,14,0,251,0,108,0,0,0,0,0,0,0,69,0,235,0,0,0,226,0,81,0,57,0,225,0,108,0,0,0,48,0,133,0,182,0,139,0,168,0,157,0,21,0,107,0,127,0,93,0,198,0,190,0,115,0,0,0,202,0,0,0,204,0,0,0,71,0,35,0,146,0,44,0,6,0,11,0,0,0,45,0,0,0,58,0,64,0,117,0,0,0,203,0,124,0,202,0,89,0,1,0,0,0,26,0,146,0,231,0,61,0,32,0,0,0,0,0,46,0,227,0,41,0,217,0,230,0,162,0,11,0,205,0,0,0,120,0,208,0,131,0,25,0,96,0,110,0,79,0,36,0,221,0,0,0,171,0,146,0,71,0,85,0,146,0,75,0,21,0,0,0,105,0);
signal scenario_full  : scenario_type := (35,31,183,31,243,31,14,31,102,31,72,31,72,30,54,31,54,30,193,31,127,31,56,31,207,31,134,31,97,31,252,31,157,31,152,31,75,31,28,31,74,31,55,31,196,31,50,31,29,31,27,31,27,30,173,31,173,30,122,31,75,31,155,31,134,31,96,31,96,30,245,31,143,31,64,31,64,30,228,31,111,31,29,31,9,31,9,30,9,29,9,28,50,31,211,31,65,31,65,30,52,31,51,31,96,31,94,31,95,31,95,30,235,31,189,31,189,30,98,31,178,31,162,31,100,31,173,31,173,30,173,29,173,28,201,31,158,31,215,31,234,31,158,31,158,30,133,31,133,30,133,29,148,31,148,30,130,31,187,31,8,31,241,31,248,31,248,30,248,29,186,31,94,31,20,31,20,30,19,31,171,31,76,31,225,31,200,31,200,30,200,29,223,31,2,31,159,31,57,31,57,30,58,31,58,30,224,31,88,31,97,31,86,31,27,31,104,31,104,30,114,31,35,31,35,30,211,31,28,31,101,31,94,31,194,31,160,31,44,31,44,30,44,29,23,31,241,31,103,31,103,30,159,31,206,31,178,31,52,31,209,31,209,30,152,31,99,31,213,31,228,31,228,30,154,31,123,31,195,31,136,31,136,30,13,31,82,31,200,31,126,31,66,31,153,31,118,31,235,31,95,31,243,31,69,31,69,30,221,31,201,31,201,30,201,29,243,31,154,31,206,31,206,30,71,31,71,30,71,29,105,31,105,30,250,31,174,31,139,31,20,31,171,31,68,31,239,31,231,31,231,30,41,31,191,31,138,31,213,31,43,31,227,31,182,31,86,31,37,31,37,30,229,31,178,31,128,31,231,31,97,31,97,30,51,31,51,30,207,31,225,31,11,31,125,31,245,31,245,30,239,31,110,31,30,31,205,31,238,31,238,30,214,31,123,31,55,31,219,31,113,31,4,31,71,31,71,30,86,31,202,31,250,31,156,31,239,31,139,31,55,31,55,30,207,31,85,31,85,30,49,31,49,30,178,31,225,31,225,30,147,31,155,31,93,31,93,30,64,31,231,31,86,31,225,31,70,31,32,31,84,31,198,31,198,30,204,31,204,30,169,31,213,31,163,31,106,31,212,31,4,31,175,31,133,31,69,31,122,31,78,31,78,30,29,31,51,31,253,31,253,30,173,31,127,31,116,31,67,31,26,31,223,31,136,31,252,31,174,31,157,31,157,30,23,31,38,31,250,31,11,31,163,31,249,31,249,30,244,31,181,31,60,31,12,31,137,31,150,31,230,31,173,31,173,30,55,31,124,31,124,30,130,31,137,31,199,31,150,31,72,31,172,31,173,31,173,30,32,31,153,31,108,31,234,31,14,31,116,31,21,31,75,31,11,31,11,30,11,29,240,31,234,31,113,31,18,31,18,30,246,31,193,31,99,31,35,31,137,31,252,31,213,31,213,30,213,29,133,31,34,31,189,31,144,31,13,31,83,31,241,31,135,31,166,31,166,30,60,31,214,31,155,31,67,31,80,31,218,31,222,31,47,31,160,31,119,31,5,31,74,31,77,31,198,31,75,31,75,30,3,31,87,31,105,31,105,30,241,31,79,31,21,31,109,31,109,30,109,29,109,28,31,31,31,30,13,31,69,31,30,31,206,31,174,31,48,31,99,31,27,31,27,30,27,29,27,28,208,31,178,31,109,31,109,30,4,31,4,30,87,31,192,31,71,31,189,31,188,31,55,31,207,31,207,30,221,31,166,31,229,31,43,31,43,30,251,31,38,31,244,31,244,30,155,31,80,31,30,31,30,30,30,29,199,31,198,31,198,30,191,31,65,31,179,31,14,31,251,31,251,30,165,31,33,31,212,31,212,30,212,29,67,31,60,31,111,31,111,30,109,31,51,31,53,31,149,31,149,30,170,31,234,31,149,31,150,31,224,31,198,31,163,31,70,31,58,31,84,31,44,31,41,31,55,31,48,31,64,31,231,31,205,31,205,30,205,29,72,31,195,31,180,31,241,31,216,31,252,31,100,31,22,31,22,30,240,31,240,30,240,29,22,31,110,31,112,31,196,31,24,31,184,31,119,31,6,31,80,31,221,31,184,31,204,31,56,31,56,30,163,31,209,31,54,31,54,30,54,29,232,31,232,30,199,31,130,31,206,31,204,31,42,31,241,31,35,31,215,31,78,31,136,31,162,31,196,31,196,30,200,31,201,31,189,31,39,31,212,31,212,30,63,31,115,31,115,30,239,31,239,30,108,31,130,31,101,31,101,30,29,31,187,31,3,31,6,31,159,31,66,31,66,30,144,31,122,31,195,31,15,31,168,31,249,31,249,30,249,29,249,28,249,31,136,31,56,31,237,31,238,31,82,31,212,31,78,31,55,31,224,31,53,31,169,31,139,31,139,30,113,31,19,31,172,31,247,31,247,30,115,31,21,31,118,31,170,31,100,31,149,31,15,31,11,31,44,31,44,30,32,31,75,31,157,31,116,31,116,30,195,31,195,30,195,29,73,31,50,31,50,30,253,31,142,31,11,31,4,31,108,31,108,30,121,31,121,30,107,31,69,31,197,31,94,31,128,31,57,31,78,31,188,31,110,31,101,31,116,31,37,31,37,30,38,31,70,31,70,30,18,31,18,30,18,29,18,28,18,27,199,31,199,30,249,31,47,31,9,31,9,30,185,31,185,30,121,31,121,30,30,31,227,31,227,30,99,31,99,30,26,31,158,31,201,31,255,31,255,30,119,31,203,31,195,31,20,31,53,31,37,31,37,30,111,31,230,31,230,30,230,29,230,28,230,27,154,31,157,31,117,31,140,31,168,31,168,30,243,31,243,30,198,31,74,31,146,31,68,31,20,31,202,31,202,30,110,31,49,31,49,30,23,31,100,31,40,31,70,31,70,30,70,29,202,31,16,31,16,30,16,29,238,31,91,31,173,31,16,31,131,31,236,31,236,30,236,29,174,31,174,30,59,31,248,31,20,31,84,31,41,31,41,30,235,31,65,31,27,31,132,31,132,30,132,29,165,31,165,30,41,31,128,31,128,30,165,31,116,31,116,30,175,31,173,31,74,31,132,31,254,31,70,31,92,31,92,30,92,29,92,28,20,31,32,31,32,30,121,31,121,30,182,31,98,31,86,31,73,31,214,31,250,31,250,30,9,31,209,31,196,31,99,31,229,31,164,31,164,30,164,29,184,31,105,31,64,31,154,31,65,31,65,30,233,31,24,31,170,31,99,31,130,31,130,30,240,31,36,31,36,30,166,31,166,30,17,31,226,31,234,31,104,31,237,31,38,31,165,31,150,31,107,31,138,31,138,30,23,31,168,31,34,31,34,30,153,31,14,31,251,31,108,31,108,30,108,29,108,28,69,31,235,31,235,30,226,31,81,31,57,31,225,31,108,31,108,30,48,31,133,31,182,31,139,31,168,31,157,31,21,31,107,31,127,31,93,31,198,31,190,31,115,31,115,30,202,31,202,30,204,31,204,30,71,31,35,31,146,31,44,31,6,31,11,31,11,30,45,31,45,30,58,31,64,31,117,31,117,30,203,31,124,31,202,31,89,31,1,31,1,30,26,31,146,31,231,31,61,31,32,31,32,30,32,29,46,31,227,31,41,31,217,31,230,31,162,31,11,31,205,31,205,30,120,31,208,31,131,31,25,31,96,31,110,31,79,31,36,31,221,31,221,30,171,31,146,31,71,31,85,31,146,31,75,31,21,31,21,30,105,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
