-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_709 is
end project_tb_709;

architecture project_tb_arch_709 of project_tb_709 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 288;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (238,0,186,0,85,0,32,0,158,0,0,0,8,0,43,0,10,0,73,0,33,0,206,0,175,0,14,0,0,0,73,0,102,0,37,0,0,0,0,0,179,0,40,0,243,0,0,0,240,0,0,0,103,0,0,0,94,0,89,0,199,0,0,0,0,0,85,0,22,0,4,0,27,0,244,0,62,0,43,0,226,0,0,0,0,0,0,0,0,0,0,0,125,0,199,0,100,0,202,0,94,0,194,0,156,0,239,0,119,0,0,0,108,0,79,0,219,0,184,0,198,0,161,0,218,0,246,0,0,0,87,0,90,0,160,0,195,0,167,0,231,0,45,0,67,0,134,0,24,0,0,0,97,0,59,0,0,0,0,0,121,0,89,0,50,0,167,0,234,0,123,0,171,0,244,0,0,0,0,0,184,0,184,0,0,0,30,0,140,0,0,0,60,0,158,0,0,0,173,0,0,0,170,0,53,0,237,0,1,0,178,0,114,0,236,0,15,0,176,0,204,0,143,0,233,0,245,0,0,0,0,0,172,0,1,0,214,0,38,0,216,0,2,0,136,0,87,0,144,0,229,0,28,0,0,0,201,0,72,0,213,0,119,0,0,0,0,0,192,0,165,0,196,0,97,0,0,0,37,0,206,0,0,0,46,0,122,0,3,0,214,0,92,0,0,0,86,0,0,0,73,0,31,0,94,0,230,0,208,0,22,0,0,0,102,0,30,0,158,0,193,0,246,0,194,0,248,0,27,0,156,0,51,0,40,0,0,0,1,0,243,0,103,0,0,0,101,0,207,0,0,0,0,0,0,0,202,0,0,0,13,0,32,0,210,0,20,0,235,0,65,0,56,0,255,0,0,0,225,0,135,0,0,0,0,0,248,0,75,0,170,0,100,0,0,0,237,0,0,0,214,0,7,0,251,0,171,0,65,0,236,0,165,0,68,0,0,0,135,0,0,0,189,0,0,0,211,0,87,0,147,0,0,0,209,0,62,0,99,0,168,0,0,0,27,0,0,0,0,0,224,0,0,0,52,0,38,0,29,0,180,0,0,0,0,0,0,0,0,0,0,0,27,0,107,0,126,0,38,0,22,0,108,0,141,0,121,0,42,0,94,0,166,0,0,0,183,0,136,0,117,0,32,0,162,0,96,0,124,0,240,0,3,0,0,0,118,0,12,0,0,0,29,0,0,0,243,0,0,0,35,0,61,0,0,0,131,0,167,0,249,0,229,0,22,0,175,0,42,0,28,0,0,0,22,0,0,0,85,0,0,0,48,0,0,0,129,0,0,0,0,0,94,0,90,0);
signal scenario_full  : scenario_type := (238,31,186,31,85,31,32,31,158,31,158,30,8,31,43,31,10,31,73,31,33,31,206,31,175,31,14,31,14,30,73,31,102,31,37,31,37,30,37,29,179,31,40,31,243,31,243,30,240,31,240,30,103,31,103,30,94,31,89,31,199,31,199,30,199,29,85,31,22,31,4,31,27,31,244,31,62,31,43,31,226,31,226,30,226,29,226,28,226,27,226,26,125,31,199,31,100,31,202,31,94,31,194,31,156,31,239,31,119,31,119,30,108,31,79,31,219,31,184,31,198,31,161,31,218,31,246,31,246,30,87,31,90,31,160,31,195,31,167,31,231,31,45,31,67,31,134,31,24,31,24,30,97,31,59,31,59,30,59,29,121,31,89,31,50,31,167,31,234,31,123,31,171,31,244,31,244,30,244,29,184,31,184,31,184,30,30,31,140,31,140,30,60,31,158,31,158,30,173,31,173,30,170,31,53,31,237,31,1,31,178,31,114,31,236,31,15,31,176,31,204,31,143,31,233,31,245,31,245,30,245,29,172,31,1,31,214,31,38,31,216,31,2,31,136,31,87,31,144,31,229,31,28,31,28,30,201,31,72,31,213,31,119,31,119,30,119,29,192,31,165,31,196,31,97,31,97,30,37,31,206,31,206,30,46,31,122,31,3,31,214,31,92,31,92,30,86,31,86,30,73,31,31,31,94,31,230,31,208,31,22,31,22,30,102,31,30,31,158,31,193,31,246,31,194,31,248,31,27,31,156,31,51,31,40,31,40,30,1,31,243,31,103,31,103,30,101,31,207,31,207,30,207,29,207,28,202,31,202,30,13,31,32,31,210,31,20,31,235,31,65,31,56,31,255,31,255,30,225,31,135,31,135,30,135,29,248,31,75,31,170,31,100,31,100,30,237,31,237,30,214,31,7,31,251,31,171,31,65,31,236,31,165,31,68,31,68,30,135,31,135,30,189,31,189,30,211,31,87,31,147,31,147,30,209,31,62,31,99,31,168,31,168,30,27,31,27,30,27,29,224,31,224,30,52,31,38,31,29,31,180,31,180,30,180,29,180,28,180,27,180,26,27,31,107,31,126,31,38,31,22,31,108,31,141,31,121,31,42,31,94,31,166,31,166,30,183,31,136,31,117,31,32,31,162,31,96,31,124,31,240,31,3,31,3,30,118,31,12,31,12,30,29,31,29,30,243,31,243,30,35,31,61,31,61,30,131,31,167,31,249,31,229,31,22,31,175,31,42,31,28,31,28,30,22,31,22,30,85,31,85,30,48,31,48,30,129,31,129,30,129,29,94,31,90,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
