-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_612 is
end project_tb_612;

architecture project_tb_arch_612 of project_tb_612 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 777;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (48,0,0,0,118,0,153,0,253,0,168,0,223,0,214,0,27,0,233,0,34,0,0,0,167,0,45,0,38,0,157,0,252,0,245,0,146,0,245,0,60,0,16,0,230,0,224,0,194,0,83,0,61,0,106,0,184,0,87,0,207,0,0,0,79,0,162,0,70,0,96,0,0,0,139,0,115,0,29,0,198,0,0,0,151,0,107,0,0,0,147,0,56,0,165,0,0,0,136,0,219,0,148,0,37,0,207,0,232,0,234,0,247,0,228,0,38,0,88,0,238,0,136,0,194,0,163,0,67,0,185,0,248,0,0,0,184,0,161,0,159,0,149,0,0,0,236,0,82,0,64,0,170,0,222,0,94,0,151,0,0,0,216,0,58,0,190,0,176,0,72,0,51,0,0,0,143,0,6,0,41,0,0,0,226,0,171,0,213,0,226,0,56,0,0,0,76,0,158,0,181,0,184,0,228,0,88,0,217,0,119,0,160,0,129,0,15,0,0,0,63,0,178,0,0,0,159,0,110,0,65,0,147,0,50,0,10,0,12,0,0,0,17,0,5,0,181,0,175,0,79,0,236,0,79,0,48,0,167,0,67,0,110,0,57,0,243,0,81,0,61,0,0,0,51,0,129,0,66,0,156,0,208,0,116,0,43,0,2,0,219,0,0,0,192,0,221,0,87,0,155,0,6,0,155,0,155,0,166,0,119,0,82,0,0,0,180,0,163,0,177,0,207,0,124,0,253,0,126,0,59,0,109,0,0,0,0,0,0,0,193,0,0,0,188,0,11,0,144,0,17,0,0,0,185,0,99,0,186,0,16,0,0,0,106,0,183,0,251,0,185,0,0,0,62,0,0,0,0,0,226,0,184,0,19,0,114,0,78,0,36,0,101,0,0,0,85,0,206,0,191,0,84,0,0,0,40,0,14,0,107,0,198,0,16,0,187,0,0,0,56,0,0,0,198,0,0,0,0,0,60,0,116,0,120,0,0,0,246,0,203,0,223,0,0,0,40,0,0,0,0,0,126,0,29,0,187,0,0,0,198,0,116,0,100,0,0,0,0,0,11,0,236,0,45,0,0,0,247,0,0,0,0,0,207,0,0,0,0,0,88,0,255,0,179,0,48,0,234,0,0,0,211,0,151,0,237,0,149,0,52,0,97,0,0,0,217,0,196,0,191,0,142,0,241,0,200,0,120,0,119,0,2,0,97,0,84,0,139,0,206,0,173,0,0,0,174,0,120,0,56,0,147,0,181,0,145,0,170,0,0,0,0,0,206,0,230,0,133,0,50,0,232,0,32,0,60,0,0,0,67,0,0,0,246,0,197,0,109,0,187,0,133,0,116,0,151,0,38,0,208,0,0,0,70,0,75,0,0,0,0,0,47,0,0,0,58,0,204,0,177,0,26,0,203,0,174,0,249,0,0,0,25,0,56,0,115,0,24,0,0,0,0,0,98,0,61,0,172,0,0,0,0,0,135,0,127,0,8,0,170,0,178,0,122,0,224,0,37,0,0,0,224,0,63,0,151,0,105,0,0,0,0,0,115,0,151,0,168,0,58,0,90,0,99,0,45,0,44,0,254,0,0,0,206,0,127,0,0,0,195,0,57,0,0,0,231,0,0,0,245,0,0,0,155,0,0,0,145,0,219,0,222,0,0,0,131,0,10,0,171,0,213,0,110,0,51,0,0,0,36,0,81,0,195,0,0,0,94,0,50,0,215,0,48,0,8,0,228,0,160,0,0,0,0,0,0,0,54,0,242,0,158,0,35,0,79,0,204,0,209,0,216,0,0,0,0,0,170,0,119,0,0,0,124,0,0,0,250,0,47,0,217,0,140,0,0,0,162,0,1,0,0,0,44,0,48,0,169,0,99,0,187,0,193,0,117,0,106,0,212,0,185,0,160,0,206,0,100,0,39,0,210,0,0,0,32,0,0,0,213,0,25,0,187,0,139,0,174,0,125,0,232,0,107,0,46,0,0,0,251,0,0,0,113,0,5,0,0,0,76,0,182,0,86,0,111,0,183,0,240,0,216,0,32,0,189,0,0,0,0,0,53,0,129,0,0,0,0,0,134,0,0,0,110,0,227,0,24,0,250,0,50,0,33,0,205,0,238,0,68,0,42,0,101,0,201,0,68,0,113,0,196,0,51,0,179,0,0,0,89,0,228,0,0,0,155,0,25,0,121,0,48,0,49,0,0,0,29,0,245,0,0,0,72,0,110,0,253,0,204,0,47,0,182,0,145,0,61,0,101,0,152,0,38,0,0,0,112,0,64,0,221,0,177,0,81,0,0,0,63,0,215,0,25,0,168,0,2,0,19,0,0,0,222,0,232,0,218,0,87,0,28,0,22,0,13,0,225,0,105,0,95,0,0,0,199,0,0,0,80,0,75,0,195,0,0,0,64,0,204,0,218,0,6,0,171,0,102,0,22,0,197,0,254,0,10,0,149,0,108,0,0,0,129,0,0,0,51,0,0,0,34,0,0,0,35,0,167,0,27,0,148,0,162,0,88,0,130,0,24,0,0,0,210,0,0,0,61,0,208,0,160,0,164,0,26,0,0,0,211,0,103,0,0,0,11,0,209,0,171,0,97,0,120,0,184,0,40,0,215,0,9,0,81,0,155,0,0,0,45,0,204,0,187,0,0,0,45,0,194,0,155,0,127,0,88,0,89,0,0,0,17,0,0,0,87,0,112,0,15,0,80,0,179,0,165,0,168,0,241,0,117,0,0,0,111,0,235,0,131,0,5,0,240,0,123,0,113,0,197,0,0,0,0,0,61,0,15,0,25,0,95,0,54,0,61,0,33,0,0,0,144,0,133,0,235,0,0,0,249,0,177,0,74,0,229,0,164,0,0,0,0,0,0,0,167,0,193,0,37,0,184,0,101,0,0,0,50,0,74,0,9,0,141,0,224,0,25,0,0,0,24,0,201,0,15,0,76,0,0,0,118,0,0,0,206,0,0,0,142,0,149,0,100,0,11,0,8,0,149,0,230,0,215,0,85,0,47,0,248,0,217,0,237,0,205,0,21,0,145,0,0,0,211,0,0,0,0,0,237,0,193,0,239,0,16,0,87,0,165,0,0,0,0,0,119,0,41,0,132,0,0,0,224,0,23,0,38,0,116,0,0,0,86,0,3,0,175,0,0,0,150,0,0,0,167,0,0,0,127,0,202,0,255,0,121,0,0,0,223,0,252,0,77,0,89,0,0,0,84,0,50,0,185,0,0,0,177,0,0,0,21,0,0,0,0,0,43,0,89,0,36,0,17,0,93,0,24,0,0,0,8,0,0,0,10,0,142,0,102,0,0,0,77,0,102,0,99,0,129,0,146,0,195,0,0,0,93,0,42,0,72,0,0,0,196,0,56,0,48,0,90,0,89,0,114,0,0,0,0,0,117,0,0,0,0,0,80,0,187,0,0,0,184,0,41,0,27,0,247,0,160,0,212,0,99,0,48,0,126,0,79,0,57,0,44,0,230,0,71,0,0,0);
signal scenario_full  : scenario_type := (48,31,48,30,118,31,153,31,253,31,168,31,223,31,214,31,27,31,233,31,34,31,34,30,167,31,45,31,38,31,157,31,252,31,245,31,146,31,245,31,60,31,16,31,230,31,224,31,194,31,83,31,61,31,106,31,184,31,87,31,207,31,207,30,79,31,162,31,70,31,96,31,96,30,139,31,115,31,29,31,198,31,198,30,151,31,107,31,107,30,147,31,56,31,165,31,165,30,136,31,219,31,148,31,37,31,207,31,232,31,234,31,247,31,228,31,38,31,88,31,238,31,136,31,194,31,163,31,67,31,185,31,248,31,248,30,184,31,161,31,159,31,149,31,149,30,236,31,82,31,64,31,170,31,222,31,94,31,151,31,151,30,216,31,58,31,190,31,176,31,72,31,51,31,51,30,143,31,6,31,41,31,41,30,226,31,171,31,213,31,226,31,56,31,56,30,76,31,158,31,181,31,184,31,228,31,88,31,217,31,119,31,160,31,129,31,15,31,15,30,63,31,178,31,178,30,159,31,110,31,65,31,147,31,50,31,10,31,12,31,12,30,17,31,5,31,181,31,175,31,79,31,236,31,79,31,48,31,167,31,67,31,110,31,57,31,243,31,81,31,61,31,61,30,51,31,129,31,66,31,156,31,208,31,116,31,43,31,2,31,219,31,219,30,192,31,221,31,87,31,155,31,6,31,155,31,155,31,166,31,119,31,82,31,82,30,180,31,163,31,177,31,207,31,124,31,253,31,126,31,59,31,109,31,109,30,109,29,109,28,193,31,193,30,188,31,11,31,144,31,17,31,17,30,185,31,99,31,186,31,16,31,16,30,106,31,183,31,251,31,185,31,185,30,62,31,62,30,62,29,226,31,184,31,19,31,114,31,78,31,36,31,101,31,101,30,85,31,206,31,191,31,84,31,84,30,40,31,14,31,107,31,198,31,16,31,187,31,187,30,56,31,56,30,198,31,198,30,198,29,60,31,116,31,120,31,120,30,246,31,203,31,223,31,223,30,40,31,40,30,40,29,126,31,29,31,187,31,187,30,198,31,116,31,100,31,100,30,100,29,11,31,236,31,45,31,45,30,247,31,247,30,247,29,207,31,207,30,207,29,88,31,255,31,179,31,48,31,234,31,234,30,211,31,151,31,237,31,149,31,52,31,97,31,97,30,217,31,196,31,191,31,142,31,241,31,200,31,120,31,119,31,2,31,97,31,84,31,139,31,206,31,173,31,173,30,174,31,120,31,56,31,147,31,181,31,145,31,170,31,170,30,170,29,206,31,230,31,133,31,50,31,232,31,32,31,60,31,60,30,67,31,67,30,246,31,197,31,109,31,187,31,133,31,116,31,151,31,38,31,208,31,208,30,70,31,75,31,75,30,75,29,47,31,47,30,58,31,204,31,177,31,26,31,203,31,174,31,249,31,249,30,25,31,56,31,115,31,24,31,24,30,24,29,98,31,61,31,172,31,172,30,172,29,135,31,127,31,8,31,170,31,178,31,122,31,224,31,37,31,37,30,224,31,63,31,151,31,105,31,105,30,105,29,115,31,151,31,168,31,58,31,90,31,99,31,45,31,44,31,254,31,254,30,206,31,127,31,127,30,195,31,57,31,57,30,231,31,231,30,245,31,245,30,155,31,155,30,145,31,219,31,222,31,222,30,131,31,10,31,171,31,213,31,110,31,51,31,51,30,36,31,81,31,195,31,195,30,94,31,50,31,215,31,48,31,8,31,228,31,160,31,160,30,160,29,160,28,54,31,242,31,158,31,35,31,79,31,204,31,209,31,216,31,216,30,216,29,170,31,119,31,119,30,124,31,124,30,250,31,47,31,217,31,140,31,140,30,162,31,1,31,1,30,44,31,48,31,169,31,99,31,187,31,193,31,117,31,106,31,212,31,185,31,160,31,206,31,100,31,39,31,210,31,210,30,32,31,32,30,213,31,25,31,187,31,139,31,174,31,125,31,232,31,107,31,46,31,46,30,251,31,251,30,113,31,5,31,5,30,76,31,182,31,86,31,111,31,183,31,240,31,216,31,32,31,189,31,189,30,189,29,53,31,129,31,129,30,129,29,134,31,134,30,110,31,227,31,24,31,250,31,50,31,33,31,205,31,238,31,68,31,42,31,101,31,201,31,68,31,113,31,196,31,51,31,179,31,179,30,89,31,228,31,228,30,155,31,25,31,121,31,48,31,49,31,49,30,29,31,245,31,245,30,72,31,110,31,253,31,204,31,47,31,182,31,145,31,61,31,101,31,152,31,38,31,38,30,112,31,64,31,221,31,177,31,81,31,81,30,63,31,215,31,25,31,168,31,2,31,19,31,19,30,222,31,232,31,218,31,87,31,28,31,22,31,13,31,225,31,105,31,95,31,95,30,199,31,199,30,80,31,75,31,195,31,195,30,64,31,204,31,218,31,6,31,171,31,102,31,22,31,197,31,254,31,10,31,149,31,108,31,108,30,129,31,129,30,51,31,51,30,34,31,34,30,35,31,167,31,27,31,148,31,162,31,88,31,130,31,24,31,24,30,210,31,210,30,61,31,208,31,160,31,164,31,26,31,26,30,211,31,103,31,103,30,11,31,209,31,171,31,97,31,120,31,184,31,40,31,215,31,9,31,81,31,155,31,155,30,45,31,204,31,187,31,187,30,45,31,194,31,155,31,127,31,88,31,89,31,89,30,17,31,17,30,87,31,112,31,15,31,80,31,179,31,165,31,168,31,241,31,117,31,117,30,111,31,235,31,131,31,5,31,240,31,123,31,113,31,197,31,197,30,197,29,61,31,15,31,25,31,95,31,54,31,61,31,33,31,33,30,144,31,133,31,235,31,235,30,249,31,177,31,74,31,229,31,164,31,164,30,164,29,164,28,167,31,193,31,37,31,184,31,101,31,101,30,50,31,74,31,9,31,141,31,224,31,25,31,25,30,24,31,201,31,15,31,76,31,76,30,118,31,118,30,206,31,206,30,142,31,149,31,100,31,11,31,8,31,149,31,230,31,215,31,85,31,47,31,248,31,217,31,237,31,205,31,21,31,145,31,145,30,211,31,211,30,211,29,237,31,193,31,239,31,16,31,87,31,165,31,165,30,165,29,119,31,41,31,132,31,132,30,224,31,23,31,38,31,116,31,116,30,86,31,3,31,175,31,175,30,150,31,150,30,167,31,167,30,127,31,202,31,255,31,121,31,121,30,223,31,252,31,77,31,89,31,89,30,84,31,50,31,185,31,185,30,177,31,177,30,21,31,21,30,21,29,43,31,89,31,36,31,17,31,93,31,24,31,24,30,8,31,8,30,10,31,142,31,102,31,102,30,77,31,102,31,99,31,129,31,146,31,195,31,195,30,93,31,42,31,72,31,72,30,196,31,56,31,48,31,90,31,89,31,114,31,114,30,114,29,117,31,117,30,117,29,80,31,187,31,187,30,184,31,41,31,27,31,247,31,160,31,212,31,99,31,48,31,126,31,79,31,57,31,44,31,230,31,71,31,71,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
