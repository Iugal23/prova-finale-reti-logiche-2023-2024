-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 364;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,184,0,139,0,69,0,0,0,56,0,0,0,183,0,190,0,218,0,0,0,50,0,101,0,231,0,109,0,66,0,247,0,0,0,76,0,198,0,64,0,138,0,57,0,0,0,55,0,90,0,96,0,64,0,131,0,0,0,7,0,0,0,0,0,83,0,6,0,195,0,117,0,218,0,71,0,33,0,167,0,133,0,0,0,0,0,190,0,2,0,137,0,131,0,31,0,166,0,217,0,0,0,225,0,17,0,216,0,96,0,221,0,119,0,0,0,104,0,123,0,0,0,0,0,230,0,205,0,213,0,189,0,91,0,0,0,247,0,169,0,0,0,204,0,0,0,100,0,141,0,178,0,248,0,216,0,190,0,100,0,216,0,58,0,47,0,34,0,187,0,53,0,84,0,86,0,11,0,168,0,0,0,230,0,61,0,123,0,0,0,38,0,141,0,204,0,96,0,40,0,138,0,187,0,0,0,89,0,137,0,210,0,231,0,22,0,6,0,0,0,0,0,138,0,12,0,0,0,116,0,130,0,0,0,67,0,136,0,71,0,26,0,164,0,29,0,238,0,0,0,222,0,50,0,250,0,0,0,216,0,146,0,73,0,0,0,131,0,114,0,0,0,175,0,174,0,100,0,154,0,228,0,113,0,0,0,130,0,126,0,0,0,245,0,1,0,223,0,238,0,237,0,227,0,228,0,216,0,122,0,23,0,222,0,209,0,219,0,0,0,52,0,107,0,0,0,209,0,19,0,150,0,218,0,162,0,249,0,43,0,59,0,0,0,0,0,194,0,0,0,107,0,64,0,197,0,167,0,122,0,147,0,177,0,0,0,48,0,75,0,153,0,251,0,109,0,193,0,7,0,128,0,184,0,0,0,59,0,56,0,202,0,87,0,0,0,0,0,37,0,203,0,0,0,171,0,213,0,187,0,0,0,0,0,14,0,195,0,183,0,183,0,172,0,0,0,251,0,81,0,29,0,0,0,120,0,32,0,116,0,99,0,167,0,19,0,0,0,0,0,120,0,202,0,0,0,71,0,44,0,128,0,107,0,231,0,90,0,221,0,70,0,112,0,0,0,205,0,9,0,160,0,0,0,174,0,204,0,251,0,149,0,162,0,0,0,27,0,190,0,71,0,150,0,0,0,227,0,240,0,8,0,0,0,199,0,200,0,39,0,44,0,65,0,0,0,30,0,109,0,89,0,250,0,0,0,0,0,94,0,116,0,6,0,220,0,80,0,116,0,213,0,242,0,0,0,187,0,218,0,199,0,0,0,199,0,0,0,147,0,105,0,0,0,12,0,133,0,186,0,42,0,160,0,114,0,51,0,172,0,34,0,212,0,144,0,18,0,0,0,78,0,0,0,0,0,92,0,6,0,228,0,74,0,62,0,98,0,162,0,0,0,186,0,0,0,220,0,0,0,52,0,80,0,37,0,196,0,95,0,188,0,169,0,0,0,30,0,11,0,0,0,249,0,0,0,0,0,0,0,0,0,98,0,98,0,87,0,136,0,0,0,237,0,221,0,210,0,156,0,70,0,125,0,117,0,129,0,119,0,29,0,24,0,88,0,23,0,98,0,42,0,113,0,107,0,178,0,0,0,11,0,61,0,232,0,210,0,231,0,76,0,0,0,190,0);
signal scenario_full  : scenario_type := (0,0,184,31,139,31,69,31,69,30,56,31,56,30,183,31,190,31,218,31,218,30,50,31,101,31,231,31,109,31,66,31,247,31,247,30,76,31,198,31,64,31,138,31,57,31,57,30,55,31,90,31,96,31,64,31,131,31,131,30,7,31,7,30,7,29,83,31,6,31,195,31,117,31,218,31,71,31,33,31,167,31,133,31,133,30,133,29,190,31,2,31,137,31,131,31,31,31,166,31,217,31,217,30,225,31,17,31,216,31,96,31,221,31,119,31,119,30,104,31,123,31,123,30,123,29,230,31,205,31,213,31,189,31,91,31,91,30,247,31,169,31,169,30,204,31,204,30,100,31,141,31,178,31,248,31,216,31,190,31,100,31,216,31,58,31,47,31,34,31,187,31,53,31,84,31,86,31,11,31,168,31,168,30,230,31,61,31,123,31,123,30,38,31,141,31,204,31,96,31,40,31,138,31,187,31,187,30,89,31,137,31,210,31,231,31,22,31,6,31,6,30,6,29,138,31,12,31,12,30,116,31,130,31,130,30,67,31,136,31,71,31,26,31,164,31,29,31,238,31,238,30,222,31,50,31,250,31,250,30,216,31,146,31,73,31,73,30,131,31,114,31,114,30,175,31,174,31,100,31,154,31,228,31,113,31,113,30,130,31,126,31,126,30,245,31,1,31,223,31,238,31,237,31,227,31,228,31,216,31,122,31,23,31,222,31,209,31,219,31,219,30,52,31,107,31,107,30,209,31,19,31,150,31,218,31,162,31,249,31,43,31,59,31,59,30,59,29,194,31,194,30,107,31,64,31,197,31,167,31,122,31,147,31,177,31,177,30,48,31,75,31,153,31,251,31,109,31,193,31,7,31,128,31,184,31,184,30,59,31,56,31,202,31,87,31,87,30,87,29,37,31,203,31,203,30,171,31,213,31,187,31,187,30,187,29,14,31,195,31,183,31,183,31,172,31,172,30,251,31,81,31,29,31,29,30,120,31,32,31,116,31,99,31,167,31,19,31,19,30,19,29,120,31,202,31,202,30,71,31,44,31,128,31,107,31,231,31,90,31,221,31,70,31,112,31,112,30,205,31,9,31,160,31,160,30,174,31,204,31,251,31,149,31,162,31,162,30,27,31,190,31,71,31,150,31,150,30,227,31,240,31,8,31,8,30,199,31,200,31,39,31,44,31,65,31,65,30,30,31,109,31,89,31,250,31,250,30,250,29,94,31,116,31,6,31,220,31,80,31,116,31,213,31,242,31,242,30,187,31,218,31,199,31,199,30,199,31,199,30,147,31,105,31,105,30,12,31,133,31,186,31,42,31,160,31,114,31,51,31,172,31,34,31,212,31,144,31,18,31,18,30,78,31,78,30,78,29,92,31,6,31,228,31,74,31,62,31,98,31,162,31,162,30,186,31,186,30,220,31,220,30,52,31,80,31,37,31,196,31,95,31,188,31,169,31,169,30,30,31,11,31,11,30,249,31,249,30,249,29,249,28,249,27,98,31,98,31,87,31,136,31,136,30,237,31,221,31,210,31,156,31,70,31,125,31,117,31,129,31,119,31,29,31,24,31,88,31,23,31,98,31,42,31,113,31,107,31,178,31,178,30,11,31,61,31,232,31,210,31,231,31,76,31,76,30,190,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
