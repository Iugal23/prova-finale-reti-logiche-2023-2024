-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_289 is
end project_tb_289;

architecture project_tb_arch_289 of project_tb_289 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 587;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (195,0,0,0,46,0,245,0,193,0,41,0,225,0,85,0,102,0,111,0,158,0,176,0,0,0,8,0,0,0,0,0,10,0,134,0,0,0,0,0,124,0,211,0,189,0,0,0,162,0,161,0,91,0,72,0,220,0,111,0,0,0,0,0,81,0,42,0,64,0,0,0,214,0,0,0,141,0,94,0,46,0,0,0,99,0,144,0,241,0,134,0,45,0,146,0,0,0,39,0,208,0,0,0,38,0,90,0,79,0,0,0,0,0,22,0,168,0,0,0,247,0,223,0,26,0,117,0,0,0,102,0,12,0,204,0,0,0,112,0,102,0,179,0,186,0,54,0,60,0,246,0,0,0,109,0,0,0,178,0,102,0,0,0,53,0,168,0,189,0,45,0,144,0,0,0,204,0,133,0,75,0,43,0,136,0,228,0,0,0,34,0,0,0,0,0,49,0,70,0,229,0,150,0,141,0,15,0,201,0,50,0,240,0,0,0,183,0,203,0,0,0,158,0,74,0,0,0,120,0,0,0,48,0,161,0,0,0,151,0,0,0,0,0,0,0,49,0,19,0,230,0,74,0,66,0,238,0,92,0,7,0,79,0,139,0,49,0,175,0,214,0,1,0,125,0,94,0,168,0,193,0,143,0,117,0,201,0,157,0,36,0,0,0,0,0,99,0,0,0,0,0,189,0,38,0,68,0,224,0,208,0,108,0,0,0,0,0,155,0,231,0,43,0,106,0,113,0,131,0,24,0,136,0,27,0,34,0,85,0,92,0,0,0,245,0,0,0,5,0,21,0,208,0,5,0,0,0,0,0,0,0,132,0,172,0,166,0,241,0,1,0,110,0,0,0,101,0,4,0,187,0,0,0,143,0,2,0,0,0,16,0,162,0,215,0,100,0,27,0,50,0,0,0,172,0,221,0,0,0,20,0,0,0,175,0,0,0,151,0,0,0,41,0,34,0,190,0,148,0,101,0,226,0,0,0,178,0,81,0,156,0,0,0,55,0,149,0,38,0,78,0,210,0,198,0,11,0,0,0,39,0,20,0,82,0,195,0,178,0,204,0,173,0,0,0,185,0,0,0,220,0,156,0,139,0,153,0,0,0,212,0,0,0,242,0,51,0,78,0,0,0,139,0,226,0,229,0,127,0,222,0,111,0,0,0,150,0,75,0,26,0,174,0,216,0,101,0,192,0,185,0,203,0,173,0,224,0,83,0,24,0,253,0,248,0,237,0,19,0,0,0,175,0,31,0,62,0,178,0,117,0,115,0,156,0,0,0,111,0,245,0,41,0,177,0,0,0,12,0,131,0,181,0,57,0,77,0,106,0,148,0,247,0,252,0,231,0,0,0,51,0,221,0,0,0,0,0,223,0,89,0,197,0,65,0,211,0,104,0,78,0,76,0,0,0,66,0,0,0,0,0,126,0,79,0,129,0,85,0,61,0,59,0,102,0,60,0,245,0,207,0,240,0,169,0,39,0,185,0,79,0,215,0,0,0,141,0,95,0,0,0,71,0,216,0,10,0,10,0,88,0,0,0,156,0,171,0,132,0,248,0,148,0,194,0,45,0,170,0,162,0,0,0,243,0,57,0,20,0,39,0,15,0,148,0,208,0,49,0,157,0,252,0,38,0,25,0,0,0,0,0,0,0,0,0,76,0,91,0,0,0,28,0,165,0,101,0,123,0,190,0,221,0,185,0,28,0,171,0,88,0,147,0,34,0,105,0,54,0,123,0,193,0,0,0,46,0,74,0,0,0,49,0,183,0,180,0,34,0,66,0,236,0,85,0,189,0,0,0,214,0,0,0,113,0,0,0,1,0,107,0,0,0,29,0,0,0,112,0,0,0,86,0,242,0,189,0,11,0,225,0,28,0,161,0,191,0,214,0,102,0,0,0,181,0,155,0,0,0,216,0,0,0,33,0,179,0,130,0,123,0,0,0,18,0,123,0,0,0,90,0,20,0,228,0,141,0,56,0,181,0,14,0,3,0,83,0,64,0,0,0,73,0,231,0,30,0,161,0,250,0,0,0,255,0,237,0,31,0,251,0,247,0,244,0,134,0,249,0,0,0,37,0,212,0,220,0,71,0,142,0,46,0,148,0,152,0,55,0,185,0,199,0,183,0,49,0,75,0,0,0,196,0,143,0,107,0,248,0,214,0,0,0,65,0,115,0,129,0,242,0,207,0,54,0,0,0,143,0,0,0,240,0,145,0,150,0,0,0,43,0,0,0,120,0,0,0,0,0,0,0,34,0,120,0,227,0,82,0,19,0,185,0,55,0,208,0,130,0,230,0,186,0,126,0,0,0,32,0,51,0,231,0,15,0,10,0,135,0,141,0,68,0,125,0,0,0,7,0,0,0,125,0,200,0,73,0,83,0,7,0,71,0,217,0,255,0,0,0,0,0,240,0,0,0,141,0,239,0,48,0,0,0,181,0,83,0,192,0,41,0,148,0,173,0,142,0,55,0,202,0,171,0,0,0,120,0,255,0,206,0,190,0,196,0,0,0,91,0,30,0,37,0,64,0,0,0,6,0,235,0,206,0,177,0,9,0,59,0,0,0,0,0,241,0,161,0,0,0,248,0,10,0,73,0,238,0,197,0,84,0,75,0,51,0,0,0,244,0,0,0,83,0);
signal scenario_full  : scenario_type := (195,31,195,30,46,31,245,31,193,31,41,31,225,31,85,31,102,31,111,31,158,31,176,31,176,30,8,31,8,30,8,29,10,31,134,31,134,30,134,29,124,31,211,31,189,31,189,30,162,31,161,31,91,31,72,31,220,31,111,31,111,30,111,29,81,31,42,31,64,31,64,30,214,31,214,30,141,31,94,31,46,31,46,30,99,31,144,31,241,31,134,31,45,31,146,31,146,30,39,31,208,31,208,30,38,31,90,31,79,31,79,30,79,29,22,31,168,31,168,30,247,31,223,31,26,31,117,31,117,30,102,31,12,31,204,31,204,30,112,31,102,31,179,31,186,31,54,31,60,31,246,31,246,30,109,31,109,30,178,31,102,31,102,30,53,31,168,31,189,31,45,31,144,31,144,30,204,31,133,31,75,31,43,31,136,31,228,31,228,30,34,31,34,30,34,29,49,31,70,31,229,31,150,31,141,31,15,31,201,31,50,31,240,31,240,30,183,31,203,31,203,30,158,31,74,31,74,30,120,31,120,30,48,31,161,31,161,30,151,31,151,30,151,29,151,28,49,31,19,31,230,31,74,31,66,31,238,31,92,31,7,31,79,31,139,31,49,31,175,31,214,31,1,31,125,31,94,31,168,31,193,31,143,31,117,31,201,31,157,31,36,31,36,30,36,29,99,31,99,30,99,29,189,31,38,31,68,31,224,31,208,31,108,31,108,30,108,29,155,31,231,31,43,31,106,31,113,31,131,31,24,31,136,31,27,31,34,31,85,31,92,31,92,30,245,31,245,30,5,31,21,31,208,31,5,31,5,30,5,29,5,28,132,31,172,31,166,31,241,31,1,31,110,31,110,30,101,31,4,31,187,31,187,30,143,31,2,31,2,30,16,31,162,31,215,31,100,31,27,31,50,31,50,30,172,31,221,31,221,30,20,31,20,30,175,31,175,30,151,31,151,30,41,31,34,31,190,31,148,31,101,31,226,31,226,30,178,31,81,31,156,31,156,30,55,31,149,31,38,31,78,31,210,31,198,31,11,31,11,30,39,31,20,31,82,31,195,31,178,31,204,31,173,31,173,30,185,31,185,30,220,31,156,31,139,31,153,31,153,30,212,31,212,30,242,31,51,31,78,31,78,30,139,31,226,31,229,31,127,31,222,31,111,31,111,30,150,31,75,31,26,31,174,31,216,31,101,31,192,31,185,31,203,31,173,31,224,31,83,31,24,31,253,31,248,31,237,31,19,31,19,30,175,31,31,31,62,31,178,31,117,31,115,31,156,31,156,30,111,31,245,31,41,31,177,31,177,30,12,31,131,31,181,31,57,31,77,31,106,31,148,31,247,31,252,31,231,31,231,30,51,31,221,31,221,30,221,29,223,31,89,31,197,31,65,31,211,31,104,31,78,31,76,31,76,30,66,31,66,30,66,29,126,31,79,31,129,31,85,31,61,31,59,31,102,31,60,31,245,31,207,31,240,31,169,31,39,31,185,31,79,31,215,31,215,30,141,31,95,31,95,30,71,31,216,31,10,31,10,31,88,31,88,30,156,31,171,31,132,31,248,31,148,31,194,31,45,31,170,31,162,31,162,30,243,31,57,31,20,31,39,31,15,31,148,31,208,31,49,31,157,31,252,31,38,31,25,31,25,30,25,29,25,28,25,27,76,31,91,31,91,30,28,31,165,31,101,31,123,31,190,31,221,31,185,31,28,31,171,31,88,31,147,31,34,31,105,31,54,31,123,31,193,31,193,30,46,31,74,31,74,30,49,31,183,31,180,31,34,31,66,31,236,31,85,31,189,31,189,30,214,31,214,30,113,31,113,30,1,31,107,31,107,30,29,31,29,30,112,31,112,30,86,31,242,31,189,31,11,31,225,31,28,31,161,31,191,31,214,31,102,31,102,30,181,31,155,31,155,30,216,31,216,30,33,31,179,31,130,31,123,31,123,30,18,31,123,31,123,30,90,31,20,31,228,31,141,31,56,31,181,31,14,31,3,31,83,31,64,31,64,30,73,31,231,31,30,31,161,31,250,31,250,30,255,31,237,31,31,31,251,31,247,31,244,31,134,31,249,31,249,30,37,31,212,31,220,31,71,31,142,31,46,31,148,31,152,31,55,31,185,31,199,31,183,31,49,31,75,31,75,30,196,31,143,31,107,31,248,31,214,31,214,30,65,31,115,31,129,31,242,31,207,31,54,31,54,30,143,31,143,30,240,31,145,31,150,31,150,30,43,31,43,30,120,31,120,30,120,29,120,28,34,31,120,31,227,31,82,31,19,31,185,31,55,31,208,31,130,31,230,31,186,31,126,31,126,30,32,31,51,31,231,31,15,31,10,31,135,31,141,31,68,31,125,31,125,30,7,31,7,30,125,31,200,31,73,31,83,31,7,31,71,31,217,31,255,31,255,30,255,29,240,31,240,30,141,31,239,31,48,31,48,30,181,31,83,31,192,31,41,31,148,31,173,31,142,31,55,31,202,31,171,31,171,30,120,31,255,31,206,31,190,31,196,31,196,30,91,31,30,31,37,31,64,31,64,30,6,31,235,31,206,31,177,31,9,31,59,31,59,30,59,29,241,31,161,31,161,30,248,31,10,31,73,31,238,31,197,31,84,31,75,31,51,31,51,30,244,31,244,30,83,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
