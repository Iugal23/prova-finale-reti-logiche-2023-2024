-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_120 is
end project_tb_120;

architecture project_tb_arch_120 of project_tb_120 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 889;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,90,0,239,0,249,0,224,0,224,0,0,0,0,0,10,0,144,0,101,0,36,0,230,0,132,0,160,0,0,0,22,0,80,0,32,0,123,0,91,0,199,0,189,0,211,0,123,0,195,0,0,0,206,0,196,0,121,0,0,0,123,0,223,0,80,0,218,0,215,0,45,0,254,0,0,0,154,0,112,0,46,0,0,0,70,0,0,0,0,0,117,0,0,0,228,0,0,0,118,0,160,0,225,0,67,0,133,0,58,0,209,0,205,0,86,0,79,0,66,0,201,0,163,0,42,0,214,0,0,0,57,0,190,0,166,0,245,0,245,0,137,0,132,0,190,0,57,0,0,0,203,0,71,0,100,0,248,0,235,0,200,0,46,0,112,0,0,0,159,0,25,0,0,0,106,0,0,0,129,0,0,0,75,0,0,0,147,0,104,0,162,0,249,0,153,0,86,0,82,0,55,0,9,0,5,0,255,0,47,0,181,0,0,0,229,0,51,0,234,0,240,0,0,0,0,0,179,0,84,0,0,0,0,0,235,0,112,0,43,0,0,0,179,0,236,0,0,0,145,0,242,0,165,0,230,0,144,0,107,0,239,0,131,0,201,0,166,0,206,0,0,0,188,0,165,0,0,0,62,0,58,0,120,0,72,0,189,0,179,0,0,0,130,0,67,0,143,0,176,0,122,0,153,0,253,0,189,0,207,0,0,0,0,0,3,0,70,0,119,0,51,0,156,0,193,0,14,0,146,0,0,0,185,0,0,0,210,0,174,0,143,0,28,0,0,0,183,0,173,0,159,0,161,0,0,0,61,0,91,0,0,0,14,0,46,0,3,0,115,0,0,0,243,0,0,0,0,0,21,0,0,0,245,0,0,0,80,0,0,0,188,0,42,0,82,0,185,0,59,0,98,0,0,0,0,0,0,0,245,0,116,0,0,0,113,0,124,0,214,0,192,0,166,0,201,0,58,0,0,0,105,0,38,0,119,0,232,0,153,0,107,0,43,0,124,0,185,0,84,0,58,0,98,0,144,0,0,0,106,0,62,0,0,0,148,0,232,0,73,0,152,0,161,0,122,0,133,0,0,0,79,0,0,0,250,0,95,0,106,0,139,0,39,0,114,0,0,0,225,0,197,0,107,0,20,0,249,0,200,0,11,0,220,0,174,0,61,0,18,0,177,0,70,0,77,0,88,0,164,0,0,0,201,0,200,0,235,0,0,0,78,0,188,0,236,0,16,0,0,0,12,0,189,0,0,0,242,0,108,0,0,0,231,0,73,0,159,0,6,0,107,0,216,0,0,0,240,0,243,0,240,0,100,0,233,0,9,0,80,0,0,0,42,0,0,0,220,0,209,0,209,0,0,0,0,0,9,0,0,0,63,0,61,0,0,0,5,0,210,0,148,0,164,0,0,0,87,0,0,0,60,0,160,0,223,0,255,0,163,0,252,0,137,0,0,0,73,0,221,0,0,0,248,0,0,0,0,0,0,0,35,0,124,0,108,0,89,0,168,0,0,0,0,0,7,0,37,0,232,0,0,0,59,0,115,0,221,0,84,0,69,0,167,0,202,0,0,0,159,0,77,0,0,0,233,0,0,0,253,0,88,0,17,0,32,0,8,0,150,0,86,0,228,0,152,0,51,0,0,0,53,0,134,0,0,0,71,0,253,0,105,0,61,0,232,0,136,0,180,0,195,0,170,0,21,0,20,0,63,0,251,0,57,0,188,0,52,0,0,0,245,0,207,0,89,0,174,0,169,0,29,0,113,0,196,0,0,0,173,0,15,0,25,0,0,0,124,0,59,0,237,0,79,0,33,0,60,0,0,0,0,0,113,0,0,0,105,0,151,0,44,0,96,0,122,0,0,0,100,0,76,0,208,0,50,0,0,0,100,0,83,0,111,0,92,0,0,0,0,0,77,0,186,0,123,0,120,0,232,0,0,0,220,0,68,0,0,0,142,0,87,0,28,0,227,0,26,0,115,0,58,0,0,0,24,0,54,0,0,0,153,0,207,0,6,0,203,0,146,0,169,0,189,0,109,0,136,0,167,0,254,0,164,0,132,0,212,0,215,0,71,0,160,0,65,0,0,0,67,0,201,0,0,0,52,0,0,0,208,0,221,0,213,0,125,0,0,0,233,0,93,0,243,0,12,0,157,0,100,0,201,0,173,0,81,0,245,0,12,0,206,0,214,0,42,0,0,0,0,0,4,0,222,0,94,0,60,0,4,0,138,0,204,0,111,0,0,0,196,0,38,0,23,0,185,0,0,0,17,0,0,0,0,0,216,0,0,0,0,0,99,0,20,0,121,0,0,0,119,0,165,0,137,0,0,0,211,0,0,0,94,0,172,0,80,0,0,0,0,0,41,0,213,0,61,0,0,0,0,0,69,0,111,0,63,0,7,0,0,0,36,0,75,0,44,0,0,0,38,0,206,0,169,0,21,0,33,0,9,0,0,0,181,0,173,0,64,0,94,0,103,0,204,0,127,0,217,0,95,0,0,0,0,0,25,0,247,0,63,0,0,0,150,0,83,0,176,0,0,0,153,0,218,0,223,0,74,0,76,0,0,0,160,0,168,0,97,0,15,0,157,0,118,0,0,0,229,0,9,0,13,0,79,0,0,0,199,0,73,0,53,0,33,0,173,0,0,0,205,0,115,0,107,0,20,0,125,0,0,0,164,0,156,0,3,0,91,0,245,0,0,0,69,0,0,0,160,0,216,0,19,0,119,0,0,0,117,0,131,0,0,0,212,0,215,0,0,0,117,0,0,0,54,0,247,0,170,0,99,0,116,0,125,0,81,0,0,0,0,0,40,0,50,0,0,0,133,0,54,0,0,0,7,0,232,0,0,0,138,0,114,0,36,0,177,0,242,0,202,0,0,0,0,0,8,0,0,0,71,0,187,0,90,0,0,0,35,0,0,0,10,0,17,0,0,0,201,0,42,0,59,0,168,0,173,0,147,0,8,0,0,0,153,0,249,0,0,0,90,0,0,0,232,0,84,0,123,0,30,0,213,0,0,0,92,0,71,0,2,0,232,0,223,0,0,0,0,0,0,0,56,0,143,0,126,0,251,0,148,0,0,0,51,0,254,0,0,0,67,0,0,0,0,0,141,0,113,0,88,0,133,0,0,0,118,0,255,0,136,0,170,0,250,0,135,0,17,0,73,0,194,0,48,0,76,0,22,0,225,0,0,0,163,0,77,0,26,0,21,0,200,0,212,0,252,0,201,0,1,0,118,0,118,0,234,0,9,0,103,0,75,0,217,0,144,0,151,0,105,0,216,0,103,0,0,0,48,0,241,0,123,0,108,0,202,0,149,0,0,0,159,0,195,0,183,0,242,0,234,0,173,0,34,0,56,0,61,0,1,0,142,0,146,0,7,0,123,0,195,0,91,0,86,0,214,0,72,0,254,0,0,0,65,0,36,0,68,0,200,0,4,0,165,0,60,0,9,0,0,0,194,0,3,0,42,0,171,0,0,0,129,0,217,0,99,0,0,0,222,0,0,0,164,0,0,0,96,0,76,0,229,0,163,0,122,0,58,0,0,0,49,0,5,0,0,0,194,0,22,0,36,0,30,0,152,0,11,0,41,0,195,0,104,0,156,0,0,0,96,0,141,0,127,0,53,0,216,0,212,0,115,0,112,0,213,0,8,0,209,0,0,0,0,0,231,0,21,0,0,0,239,0,114,0,254,0,9,0,133,0,239,0,150,0,35,0,131,0,105,0,0,0,0,0,199,0,56,0,88,0,231,0,0,0,212,0,88,0,3,0,0,0,198,0,222,0,233,0,79,0,0,0,61,0,27,0,0,0,0,0,0,0,242,0,162,0,3,0,140,0,15,0,193,0,161,0,48,0,252,0,20,0,32,0,187,0,115,0,71,0,0,0,24,0,18,0,0,0,94,0,178,0,0,0,30,0,0,0,0,0,192,0,142,0,200,0,227,0,74,0,206,0,191,0,0,0,112,0,173,0,0,0,66,0);
signal scenario_full  : scenario_type := (0,0,0,0,90,31,239,31,249,31,224,31,224,31,224,30,224,29,10,31,144,31,101,31,36,31,230,31,132,31,160,31,160,30,22,31,80,31,32,31,123,31,91,31,199,31,189,31,211,31,123,31,195,31,195,30,206,31,196,31,121,31,121,30,123,31,223,31,80,31,218,31,215,31,45,31,254,31,254,30,154,31,112,31,46,31,46,30,70,31,70,30,70,29,117,31,117,30,228,31,228,30,118,31,160,31,225,31,67,31,133,31,58,31,209,31,205,31,86,31,79,31,66,31,201,31,163,31,42,31,214,31,214,30,57,31,190,31,166,31,245,31,245,31,137,31,132,31,190,31,57,31,57,30,203,31,71,31,100,31,248,31,235,31,200,31,46,31,112,31,112,30,159,31,25,31,25,30,106,31,106,30,129,31,129,30,75,31,75,30,147,31,104,31,162,31,249,31,153,31,86,31,82,31,55,31,9,31,5,31,255,31,47,31,181,31,181,30,229,31,51,31,234,31,240,31,240,30,240,29,179,31,84,31,84,30,84,29,235,31,112,31,43,31,43,30,179,31,236,31,236,30,145,31,242,31,165,31,230,31,144,31,107,31,239,31,131,31,201,31,166,31,206,31,206,30,188,31,165,31,165,30,62,31,58,31,120,31,72,31,189,31,179,31,179,30,130,31,67,31,143,31,176,31,122,31,153,31,253,31,189,31,207,31,207,30,207,29,3,31,70,31,119,31,51,31,156,31,193,31,14,31,146,31,146,30,185,31,185,30,210,31,174,31,143,31,28,31,28,30,183,31,173,31,159,31,161,31,161,30,61,31,91,31,91,30,14,31,46,31,3,31,115,31,115,30,243,31,243,30,243,29,21,31,21,30,245,31,245,30,80,31,80,30,188,31,42,31,82,31,185,31,59,31,98,31,98,30,98,29,98,28,245,31,116,31,116,30,113,31,124,31,214,31,192,31,166,31,201,31,58,31,58,30,105,31,38,31,119,31,232,31,153,31,107,31,43,31,124,31,185,31,84,31,58,31,98,31,144,31,144,30,106,31,62,31,62,30,148,31,232,31,73,31,152,31,161,31,122,31,133,31,133,30,79,31,79,30,250,31,95,31,106,31,139,31,39,31,114,31,114,30,225,31,197,31,107,31,20,31,249,31,200,31,11,31,220,31,174,31,61,31,18,31,177,31,70,31,77,31,88,31,164,31,164,30,201,31,200,31,235,31,235,30,78,31,188,31,236,31,16,31,16,30,12,31,189,31,189,30,242,31,108,31,108,30,231,31,73,31,159,31,6,31,107,31,216,31,216,30,240,31,243,31,240,31,100,31,233,31,9,31,80,31,80,30,42,31,42,30,220,31,209,31,209,31,209,30,209,29,9,31,9,30,63,31,61,31,61,30,5,31,210,31,148,31,164,31,164,30,87,31,87,30,60,31,160,31,223,31,255,31,163,31,252,31,137,31,137,30,73,31,221,31,221,30,248,31,248,30,248,29,248,28,35,31,124,31,108,31,89,31,168,31,168,30,168,29,7,31,37,31,232,31,232,30,59,31,115,31,221,31,84,31,69,31,167,31,202,31,202,30,159,31,77,31,77,30,233,31,233,30,253,31,88,31,17,31,32,31,8,31,150,31,86,31,228,31,152,31,51,31,51,30,53,31,134,31,134,30,71,31,253,31,105,31,61,31,232,31,136,31,180,31,195,31,170,31,21,31,20,31,63,31,251,31,57,31,188,31,52,31,52,30,245,31,207,31,89,31,174,31,169,31,29,31,113,31,196,31,196,30,173,31,15,31,25,31,25,30,124,31,59,31,237,31,79,31,33,31,60,31,60,30,60,29,113,31,113,30,105,31,151,31,44,31,96,31,122,31,122,30,100,31,76,31,208,31,50,31,50,30,100,31,83,31,111,31,92,31,92,30,92,29,77,31,186,31,123,31,120,31,232,31,232,30,220,31,68,31,68,30,142,31,87,31,28,31,227,31,26,31,115,31,58,31,58,30,24,31,54,31,54,30,153,31,207,31,6,31,203,31,146,31,169,31,189,31,109,31,136,31,167,31,254,31,164,31,132,31,212,31,215,31,71,31,160,31,65,31,65,30,67,31,201,31,201,30,52,31,52,30,208,31,221,31,213,31,125,31,125,30,233,31,93,31,243,31,12,31,157,31,100,31,201,31,173,31,81,31,245,31,12,31,206,31,214,31,42,31,42,30,42,29,4,31,222,31,94,31,60,31,4,31,138,31,204,31,111,31,111,30,196,31,38,31,23,31,185,31,185,30,17,31,17,30,17,29,216,31,216,30,216,29,99,31,20,31,121,31,121,30,119,31,165,31,137,31,137,30,211,31,211,30,94,31,172,31,80,31,80,30,80,29,41,31,213,31,61,31,61,30,61,29,69,31,111,31,63,31,7,31,7,30,36,31,75,31,44,31,44,30,38,31,206,31,169,31,21,31,33,31,9,31,9,30,181,31,173,31,64,31,94,31,103,31,204,31,127,31,217,31,95,31,95,30,95,29,25,31,247,31,63,31,63,30,150,31,83,31,176,31,176,30,153,31,218,31,223,31,74,31,76,31,76,30,160,31,168,31,97,31,15,31,157,31,118,31,118,30,229,31,9,31,13,31,79,31,79,30,199,31,73,31,53,31,33,31,173,31,173,30,205,31,115,31,107,31,20,31,125,31,125,30,164,31,156,31,3,31,91,31,245,31,245,30,69,31,69,30,160,31,216,31,19,31,119,31,119,30,117,31,131,31,131,30,212,31,215,31,215,30,117,31,117,30,54,31,247,31,170,31,99,31,116,31,125,31,81,31,81,30,81,29,40,31,50,31,50,30,133,31,54,31,54,30,7,31,232,31,232,30,138,31,114,31,36,31,177,31,242,31,202,31,202,30,202,29,8,31,8,30,71,31,187,31,90,31,90,30,35,31,35,30,10,31,17,31,17,30,201,31,42,31,59,31,168,31,173,31,147,31,8,31,8,30,153,31,249,31,249,30,90,31,90,30,232,31,84,31,123,31,30,31,213,31,213,30,92,31,71,31,2,31,232,31,223,31,223,30,223,29,223,28,56,31,143,31,126,31,251,31,148,31,148,30,51,31,254,31,254,30,67,31,67,30,67,29,141,31,113,31,88,31,133,31,133,30,118,31,255,31,136,31,170,31,250,31,135,31,17,31,73,31,194,31,48,31,76,31,22,31,225,31,225,30,163,31,77,31,26,31,21,31,200,31,212,31,252,31,201,31,1,31,118,31,118,31,234,31,9,31,103,31,75,31,217,31,144,31,151,31,105,31,216,31,103,31,103,30,48,31,241,31,123,31,108,31,202,31,149,31,149,30,159,31,195,31,183,31,242,31,234,31,173,31,34,31,56,31,61,31,1,31,142,31,146,31,7,31,123,31,195,31,91,31,86,31,214,31,72,31,254,31,254,30,65,31,36,31,68,31,200,31,4,31,165,31,60,31,9,31,9,30,194,31,3,31,42,31,171,31,171,30,129,31,217,31,99,31,99,30,222,31,222,30,164,31,164,30,96,31,76,31,229,31,163,31,122,31,58,31,58,30,49,31,5,31,5,30,194,31,22,31,36,31,30,31,152,31,11,31,41,31,195,31,104,31,156,31,156,30,96,31,141,31,127,31,53,31,216,31,212,31,115,31,112,31,213,31,8,31,209,31,209,30,209,29,231,31,21,31,21,30,239,31,114,31,254,31,9,31,133,31,239,31,150,31,35,31,131,31,105,31,105,30,105,29,199,31,56,31,88,31,231,31,231,30,212,31,88,31,3,31,3,30,198,31,222,31,233,31,79,31,79,30,61,31,27,31,27,30,27,29,27,28,242,31,162,31,3,31,140,31,15,31,193,31,161,31,48,31,252,31,20,31,32,31,187,31,115,31,71,31,71,30,24,31,18,31,18,30,94,31,178,31,178,30,30,31,30,30,30,29,192,31,142,31,200,31,227,31,74,31,206,31,191,31,191,30,112,31,173,31,173,30,66,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
