-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 966;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (40,0,116,0,154,0,254,0,198,0,13,0,2,0,0,0,0,0,81,0,181,0,233,0,60,0,42,0,80,0,74,0,187,0,10,0,0,0,245,0,132,0,252,0,223,0,9,0,213,0,0,0,90,0,0,0,223,0,0,0,0,0,161,0,141,0,52,0,225,0,0,0,90,0,143,0,191,0,0,0,87,0,201,0,0,0,66,0,105,0,7,0,81,0,56,0,12,0,153,0,28,0,252,0,189,0,77,0,0,0,48,0,174,0,113,0,249,0,82,0,145,0,184,0,189,0,149,0,132,0,248,0,72,0,85,0,66,0,116,0,11,0,55,0,0,0,19,0,146,0,0,0,0,0,144,0,0,0,105,0,159,0,51,0,181,0,190,0,90,0,255,0,0,0,238,0,34,0,0,0,133,0,175,0,101,0,79,0,0,0,219,0,141,0,12,0,0,0,181,0,0,0,128,0,207,0,87,0,0,0,0,0,4,0,0,0,81,0,0,0,188,0,54,0,22,0,0,0,114,0,193,0,0,0,203,0,92,0,229,0,76,0,75,0,56,0,21,0,237,0,57,0,49,0,140,0,151,0,206,0,118,0,0,0,0,0,124,0,166,0,164,0,0,0,129,0,0,0,248,0,184,0,165,0,61,0,245,0,0,0,189,0,242,0,33,0,166,0,102,0,0,0,193,0,0,0,20,0,68,0,175,0,186,0,0,0,216,0,80,0,224,0,0,0,18,0,192,0,51,0,116,0,140,0,20,0,171,0,127,0,8,0,108,0,173,0,134,0,19,0,201,0,163,0,194,0,199,0,0,0,75,0,210,0,8,0,203,0,61,0,149,0,251,0,242,0,0,0,231,0,129,0,0,0,9,0,0,0,238,0,218,0,120,0,0,0,227,0,110,0,20,0,0,0,0,0,74,0,210,0,73,0,179,0,237,0,0,0,0,0,89,0,3,0,238,0,215,0,131,0,241,0,169,0,18,0,61,0,108,0,102,0,189,0,89,0,223,0,222,0,40,0,149,0,30,0,91,0,32,0,12,0,149,0,144,0,52,0,249,0,0,0,230,0,0,0,156,0,124,0,188,0,203,0,172,0,216,0,0,0,82,0,52,0,0,0,101,0,145,0,78,0,238,0,112,0,7,0,0,0,210,0,208,0,0,0,251,0,243,0,0,0,193,0,130,0,157,0,91,0,0,0,0,0,236,0,5,0,92,0,54,0,0,0,0,0,89,0,94,0,96,0,93,0,29,0,0,0,117,0,238,0,184,0,91,0,165,0,1,0,182,0,197,0,219,0,89,0,185,0,151,0,193,0,158,0,213,0,69,0,132,0,30,0,129,0,0,0,243,0,78,0,137,0,194,0,186,0,111,0,210,0,34,0,22,0,35,0,195,0,163,0,0,0,229,0,122,0,159,0,161,0,113,0,51,0,207,0,214,0,0,0,66,0,122,0,224,0,76,0,44,0,0,0,234,0,156,0,0,0,164,0,54,0,26,0,204,0,32,0,183,0,15,0,0,0,146,0,248,0,159,0,46,0,0,0,150,0,21,0,4,0,144,0,61,0,58,0,171,0,0,0,243,0,213,0,231,0,116,0,123,0,115,0,13,0,0,0,151,0,200,0,107,0,234,0,197,0,70,0,25,0,88,0,0,0,81,0,177,0,100,0,113,0,187,0,46,0,0,0,15,0,191,0,0,0,135,0,251,0,36,0,107,0,11,0,0,0,51,0,0,0,107,0,186,0,68,0,103,0,124,0,189,0,107,0,12,0,14,0,229,0,0,0,42,0,0,0,50,0,116,0,226,0,42,0,68,0,200,0,241,0,0,0,41,0,153,0,195,0,172,0,144,0,154,0,234,0,95,0,72,0,68,0,0,0,136,0,42,0,226,0,206,0,145,0,66,0,114,0,240,0,253,0,177,0,203,0,167,0,100,0,186,0,248,0,123,0,0,0,0,0,136,0,0,0,84,0,24,0,0,0,0,0,106,0,135,0,244,0,0,0,18,0,96,0,0,0,156,0,111,0,25,0,98,0,107,0,0,0,0,0,92,0,22,0,151,0,66,0,233,0,184,0,0,0,59,0,223,0,64,0,33,0,237,0,180,0,0,0,186,0,0,0,180,0,255,0,251,0,75,0,0,0,26,0,195,0,212,0,17,0,0,0,130,0,155,0,204,0,117,0,49,0,0,0,47,0,121,0,0,0,0,0,0,0,83,0,0,0,117,0,78,0,0,0,29,0,11,0,211,0,177,0,0,0,240,0,112,0,0,0,202,0,0,0,235,0,0,0,149,0,108,0,152,0,39,0,191,0,0,0,0,0,225,0,105,0,208,0,0,0,175,0,0,0,73,0,159,0,248,0,0,0,64,0,208,0,237,0,50,0,6,0,239,0,40,0,107,0,178,0,25,0,68,0,61,0,0,0,173,0,0,0,224,0,220,0,127,0,59,0,71,0,81,0,116,0,141,0,0,0,59,0,132,0,240,0,56,0,149,0,49,0,105,0,0,0,184,0,127,0,247,0,82,0,0,0,37,0,67,0,0,0,101,0,122,0,163,0,222,0,82,0,28,0,0,0,89,0,80,0,154,0,62,0,202,0,0,0,1,0,144,0,154,0,145,0,114,0,246,0,237,0,98,0,117,0,0,0,224,0,0,0,73,0,196,0,114,0,0,0,224,0,208,0,101,0,237,0,182,0,137,0,0,0,239,0,0,0,124,0,0,0,0,0,0,0,68,0,195,0,186,0,6,0,137,0,209,0,180,0,244,0,237,0,0,0,161,0,0,0,101,0,234,0,82,0,229,0,21,0,119,0,111,0,0,0,76,0,22,0,70,0,21,0,178,0,235,0,79,0,181,0,6,0,0,0,129,0,0,0,0,0,223,0,101,0,27,0,245,0,27,0,228,0,107,0,0,0,0,0,115,0,0,0,230,0,100,0,185,0,209,0,103,0,82,0,251,0,126,0,80,0,245,0,198,0,0,0,0,0,168,0,176,0,33,0,163,0,29,0,22,0,134,0,163,0,114,0,187,0,0,0,120,0,204,0,168,0,42,0,185,0,0,0,115,0,0,0,154,0,199,0,93,0,16,0,218,0,121,0,0,0,34,0,148,0,79,0,79,0,180,0,213,0,105,0,0,0,182,0,115,0,6,0,113,0,52,0,0,0,38,0,175,0,0,0,141,0,228,0,96,0,4,0,0,0,0,0,209,0,200,0,153,0,0,0,0,0,73,0,172,0,99,0,34,0,0,0,248,0,0,0,141,0,223,0,119,0,16,0,77,0,0,0,132,0,177,0,250,0,242,0,109,0,221,0,175,0,216,0,20,0,0,0,84,0,67,0,129,0,115,0,0,0,71,0,69,0,238,0,68,0,32,0,204,0,157,0,161,0,0,0,3,0,64,0,72,0,241,0,206,0,248,0,35,0,0,0,234,0,48,0,172,0,0,0,168,0,0,0,225,0,57,0,163,0,0,0,104,0,27,0,45,0,0,0,166,0,143,0,54,0,207,0,243,0,162,0,232,0,0,0,0,0,214,0,2,0,66,0,0,0,7,0,28,0,5,0,193,0,0,0,101,0,0,0,168,0,0,0,225,0,0,0,72,0,5,0,249,0,89,0,0,0,0,0,0,0,43,0,208,0,62,0,133,0,206,0,125,0,0,0,48,0,0,0,0,0,82,0,0,0,159,0,248,0,106,0,3,0,0,0,108,0,133,0,27,0,57,0,16,0,143,0,235,0,176,0,43,0,57,0,0,0,151,0,168,0,0,0,238,0,99,0,119,0,148,0,15,0,184,0,67,0,75,0,0,0,202,0,16,0,9,0,52,0,148,0,108,0,161,0,0,0,145,0,31,0,148,0,245,0,59,0,0,0,38,0,57,0,176,0,205,0,134,0,0,0,49,0,218,0,233,0,134,0,235,0,0,0,131,0,104,0,0,0,75,0,32,0,110,0,215,0,0,0,244,0,241,0,0,0,0,0,140,0,75,0,31,0,0,0,207,0,241,0,253,0,34,0,111,0,171,0,0,0,249,0,187,0,183,0,96,0,147,0,161,0,106,0,129,0,232,0,63,0,0,0,57,0,30,0,23,0,72,0,249,0,0,0,0,0,84,0,175,0,123,0,55,0,0,0,222,0,148,0,220,0,181,0,103,0,0,0,52,0,29,0,225,0,161,0,0,0,0,0,198,0,201,0,120,0,16,0,76,0,235,0,45,0,91,0,0,0,226,0,159,0,120,0,239,0,159,0,245,0,49,0,0,0,245,0,0,0,0,0,0,0,74,0,231,0,0,0,70,0,207,0,0,0,239,0,109,0,77,0,253,0,0,0);
signal scenario_full  : scenario_type := (40,31,116,31,154,31,254,31,198,31,13,31,2,31,2,30,2,29,81,31,181,31,233,31,60,31,42,31,80,31,74,31,187,31,10,31,10,30,245,31,132,31,252,31,223,31,9,31,213,31,213,30,90,31,90,30,223,31,223,30,223,29,161,31,141,31,52,31,225,31,225,30,90,31,143,31,191,31,191,30,87,31,201,31,201,30,66,31,105,31,7,31,81,31,56,31,12,31,153,31,28,31,252,31,189,31,77,31,77,30,48,31,174,31,113,31,249,31,82,31,145,31,184,31,189,31,149,31,132,31,248,31,72,31,85,31,66,31,116,31,11,31,55,31,55,30,19,31,146,31,146,30,146,29,144,31,144,30,105,31,159,31,51,31,181,31,190,31,90,31,255,31,255,30,238,31,34,31,34,30,133,31,175,31,101,31,79,31,79,30,219,31,141,31,12,31,12,30,181,31,181,30,128,31,207,31,87,31,87,30,87,29,4,31,4,30,81,31,81,30,188,31,54,31,22,31,22,30,114,31,193,31,193,30,203,31,92,31,229,31,76,31,75,31,56,31,21,31,237,31,57,31,49,31,140,31,151,31,206,31,118,31,118,30,118,29,124,31,166,31,164,31,164,30,129,31,129,30,248,31,184,31,165,31,61,31,245,31,245,30,189,31,242,31,33,31,166,31,102,31,102,30,193,31,193,30,20,31,68,31,175,31,186,31,186,30,216,31,80,31,224,31,224,30,18,31,192,31,51,31,116,31,140,31,20,31,171,31,127,31,8,31,108,31,173,31,134,31,19,31,201,31,163,31,194,31,199,31,199,30,75,31,210,31,8,31,203,31,61,31,149,31,251,31,242,31,242,30,231,31,129,31,129,30,9,31,9,30,238,31,218,31,120,31,120,30,227,31,110,31,20,31,20,30,20,29,74,31,210,31,73,31,179,31,237,31,237,30,237,29,89,31,3,31,238,31,215,31,131,31,241,31,169,31,18,31,61,31,108,31,102,31,189,31,89,31,223,31,222,31,40,31,149,31,30,31,91,31,32,31,12,31,149,31,144,31,52,31,249,31,249,30,230,31,230,30,156,31,124,31,188,31,203,31,172,31,216,31,216,30,82,31,52,31,52,30,101,31,145,31,78,31,238,31,112,31,7,31,7,30,210,31,208,31,208,30,251,31,243,31,243,30,193,31,130,31,157,31,91,31,91,30,91,29,236,31,5,31,92,31,54,31,54,30,54,29,89,31,94,31,96,31,93,31,29,31,29,30,117,31,238,31,184,31,91,31,165,31,1,31,182,31,197,31,219,31,89,31,185,31,151,31,193,31,158,31,213,31,69,31,132,31,30,31,129,31,129,30,243,31,78,31,137,31,194,31,186,31,111,31,210,31,34,31,22,31,35,31,195,31,163,31,163,30,229,31,122,31,159,31,161,31,113,31,51,31,207,31,214,31,214,30,66,31,122,31,224,31,76,31,44,31,44,30,234,31,156,31,156,30,164,31,54,31,26,31,204,31,32,31,183,31,15,31,15,30,146,31,248,31,159,31,46,31,46,30,150,31,21,31,4,31,144,31,61,31,58,31,171,31,171,30,243,31,213,31,231,31,116,31,123,31,115,31,13,31,13,30,151,31,200,31,107,31,234,31,197,31,70,31,25,31,88,31,88,30,81,31,177,31,100,31,113,31,187,31,46,31,46,30,15,31,191,31,191,30,135,31,251,31,36,31,107,31,11,31,11,30,51,31,51,30,107,31,186,31,68,31,103,31,124,31,189,31,107,31,12,31,14,31,229,31,229,30,42,31,42,30,50,31,116,31,226,31,42,31,68,31,200,31,241,31,241,30,41,31,153,31,195,31,172,31,144,31,154,31,234,31,95,31,72,31,68,31,68,30,136,31,42,31,226,31,206,31,145,31,66,31,114,31,240,31,253,31,177,31,203,31,167,31,100,31,186,31,248,31,123,31,123,30,123,29,136,31,136,30,84,31,24,31,24,30,24,29,106,31,135,31,244,31,244,30,18,31,96,31,96,30,156,31,111,31,25,31,98,31,107,31,107,30,107,29,92,31,22,31,151,31,66,31,233,31,184,31,184,30,59,31,223,31,64,31,33,31,237,31,180,31,180,30,186,31,186,30,180,31,255,31,251,31,75,31,75,30,26,31,195,31,212,31,17,31,17,30,130,31,155,31,204,31,117,31,49,31,49,30,47,31,121,31,121,30,121,29,121,28,83,31,83,30,117,31,78,31,78,30,29,31,11,31,211,31,177,31,177,30,240,31,112,31,112,30,202,31,202,30,235,31,235,30,149,31,108,31,152,31,39,31,191,31,191,30,191,29,225,31,105,31,208,31,208,30,175,31,175,30,73,31,159,31,248,31,248,30,64,31,208,31,237,31,50,31,6,31,239,31,40,31,107,31,178,31,25,31,68,31,61,31,61,30,173,31,173,30,224,31,220,31,127,31,59,31,71,31,81,31,116,31,141,31,141,30,59,31,132,31,240,31,56,31,149,31,49,31,105,31,105,30,184,31,127,31,247,31,82,31,82,30,37,31,67,31,67,30,101,31,122,31,163,31,222,31,82,31,28,31,28,30,89,31,80,31,154,31,62,31,202,31,202,30,1,31,144,31,154,31,145,31,114,31,246,31,237,31,98,31,117,31,117,30,224,31,224,30,73,31,196,31,114,31,114,30,224,31,208,31,101,31,237,31,182,31,137,31,137,30,239,31,239,30,124,31,124,30,124,29,124,28,68,31,195,31,186,31,6,31,137,31,209,31,180,31,244,31,237,31,237,30,161,31,161,30,101,31,234,31,82,31,229,31,21,31,119,31,111,31,111,30,76,31,22,31,70,31,21,31,178,31,235,31,79,31,181,31,6,31,6,30,129,31,129,30,129,29,223,31,101,31,27,31,245,31,27,31,228,31,107,31,107,30,107,29,115,31,115,30,230,31,100,31,185,31,209,31,103,31,82,31,251,31,126,31,80,31,245,31,198,31,198,30,198,29,168,31,176,31,33,31,163,31,29,31,22,31,134,31,163,31,114,31,187,31,187,30,120,31,204,31,168,31,42,31,185,31,185,30,115,31,115,30,154,31,199,31,93,31,16,31,218,31,121,31,121,30,34,31,148,31,79,31,79,31,180,31,213,31,105,31,105,30,182,31,115,31,6,31,113,31,52,31,52,30,38,31,175,31,175,30,141,31,228,31,96,31,4,31,4,30,4,29,209,31,200,31,153,31,153,30,153,29,73,31,172,31,99,31,34,31,34,30,248,31,248,30,141,31,223,31,119,31,16,31,77,31,77,30,132,31,177,31,250,31,242,31,109,31,221,31,175,31,216,31,20,31,20,30,84,31,67,31,129,31,115,31,115,30,71,31,69,31,238,31,68,31,32,31,204,31,157,31,161,31,161,30,3,31,64,31,72,31,241,31,206,31,248,31,35,31,35,30,234,31,48,31,172,31,172,30,168,31,168,30,225,31,57,31,163,31,163,30,104,31,27,31,45,31,45,30,166,31,143,31,54,31,207,31,243,31,162,31,232,31,232,30,232,29,214,31,2,31,66,31,66,30,7,31,28,31,5,31,193,31,193,30,101,31,101,30,168,31,168,30,225,31,225,30,72,31,5,31,249,31,89,31,89,30,89,29,89,28,43,31,208,31,62,31,133,31,206,31,125,31,125,30,48,31,48,30,48,29,82,31,82,30,159,31,248,31,106,31,3,31,3,30,108,31,133,31,27,31,57,31,16,31,143,31,235,31,176,31,43,31,57,31,57,30,151,31,168,31,168,30,238,31,99,31,119,31,148,31,15,31,184,31,67,31,75,31,75,30,202,31,16,31,9,31,52,31,148,31,108,31,161,31,161,30,145,31,31,31,148,31,245,31,59,31,59,30,38,31,57,31,176,31,205,31,134,31,134,30,49,31,218,31,233,31,134,31,235,31,235,30,131,31,104,31,104,30,75,31,32,31,110,31,215,31,215,30,244,31,241,31,241,30,241,29,140,31,75,31,31,31,31,30,207,31,241,31,253,31,34,31,111,31,171,31,171,30,249,31,187,31,183,31,96,31,147,31,161,31,106,31,129,31,232,31,63,31,63,30,57,31,30,31,23,31,72,31,249,31,249,30,249,29,84,31,175,31,123,31,55,31,55,30,222,31,148,31,220,31,181,31,103,31,103,30,52,31,29,31,225,31,161,31,161,30,161,29,198,31,201,31,120,31,16,31,76,31,235,31,45,31,91,31,91,30,226,31,159,31,120,31,239,31,159,31,245,31,49,31,49,30,245,31,245,30,245,29,245,28,74,31,231,31,231,30,70,31,207,31,207,30,239,31,109,31,77,31,253,31,253,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
