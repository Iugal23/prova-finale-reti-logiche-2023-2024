-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_806 is
end project_tb_806;

architecture project_tb_arch_806 of project_tb_806 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 316;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,73,0,0,0,252,0,237,0,4,0,69,0,81,0,0,0,0,0,13,0,148,0,23,0,0,0,0,0,0,0,189,0,78,0,54,0,83,0,120,0,210,0,126,0,48,0,0,0,157,0,13,0,0,0,253,0,59,0,0,0,171,0,194,0,0,0,220,0,122,0,0,0,40,0,143,0,12,0,209,0,165,0,0,0,22,0,82,0,9,0,171,0,11,0,32,0,246,0,124,0,0,0,126,0,176,0,0,0,33,0,221,0,52,0,0,0,0,0,175,0,0,0,61,0,150,0,177,0,225,0,0,0,236,0,183,0,33,0,159,0,0,0,77,0,62,0,179,0,249,0,221,0,201,0,113,0,220,0,146,0,47,0,0,0,0,0,143,0,81,0,177,0,61,0,52,0,0,0,54,0,190,0,115,0,75,0,122,0,245,0,52,0,132,0,34,0,204,0,227,0,125,0,86,0,0,0,14,0,32,0,0,0,113,0,0,0,0,0,55,0,16,0,31,0,114,0,207,0,76,0,94,0,192,0,0,0,0,0,205,0,0,0,0,0,0,0,0,0,129,0,175,0,166,0,245,0,80,0,202,0,131,0,102,0,84,0,55,0,93,0,80,0,17,0,200,0,191,0,0,0,226,0,178,0,242,0,224,0,196,0,0,0,85,0,115,0,132,0,47,0,75,0,227,0,168,0,150,0,221,0,130,0,250,0,0,0,0,0,144,0,8,0,215,0,8,0,120,0,0,0,192,0,42,0,103,0,111,0,236,0,121,0,0,0,90,0,102,0,153,0,167,0,14,0,191,0,0,0,197,0,0,0,194,0,62,0,0,0,0,0,35,0,8,0,21,0,0,0,203,0,41,0,87,0,0,0,0,0,0,0,19,0,161,0,0,0,129,0,190,0,47,0,0,0,211,0,0,0,172,0,0,0,17,0,66,0,234,0,81,0,220,0,165,0,111,0,0,0,0,0,199,0,159,0,18,0,244,0,0,0,249,0,0,0,211,0,75,0,193,0,0,0,189,0,137,0,0,0,30,0,217,0,107,0,206,0,0,0,36,0,113,0,187,0,0,0,0,0,114,0,223,0,223,0,158,0,0,0,0,0,232,0,191,0,0,0,122,0,144,0,218,0,178,0,28,0,34,0,69,0,0,0,23,0,144,0,55,0,24,0,122,0,0,0,13,0,134,0,0,0,158,0,103,0,217,0,67,0,0,0,0,0,179,0,239,0,0,0,0,0,68,0,12,0,146,0,216,0,222,0,38,0,150,0,227,0,111,0,36,0,119,0,221,0,120,0,101,0,136,0,1,0,163,0,171,0,169,0,64,0,60,0,133,0,167,0,0,0,0,0,226,0,143,0,0,0,0,0,77,0,0,0,187,0,121,0,0,0,207,0,200,0,0,0,194,0,164,0,0,0);
signal scenario_full  : scenario_type := (0,0,73,31,73,30,252,31,237,31,4,31,69,31,81,31,81,30,81,29,13,31,148,31,23,31,23,30,23,29,23,28,189,31,78,31,54,31,83,31,120,31,210,31,126,31,48,31,48,30,157,31,13,31,13,30,253,31,59,31,59,30,171,31,194,31,194,30,220,31,122,31,122,30,40,31,143,31,12,31,209,31,165,31,165,30,22,31,82,31,9,31,171,31,11,31,32,31,246,31,124,31,124,30,126,31,176,31,176,30,33,31,221,31,52,31,52,30,52,29,175,31,175,30,61,31,150,31,177,31,225,31,225,30,236,31,183,31,33,31,159,31,159,30,77,31,62,31,179,31,249,31,221,31,201,31,113,31,220,31,146,31,47,31,47,30,47,29,143,31,81,31,177,31,61,31,52,31,52,30,54,31,190,31,115,31,75,31,122,31,245,31,52,31,132,31,34,31,204,31,227,31,125,31,86,31,86,30,14,31,32,31,32,30,113,31,113,30,113,29,55,31,16,31,31,31,114,31,207,31,76,31,94,31,192,31,192,30,192,29,205,31,205,30,205,29,205,28,205,27,129,31,175,31,166,31,245,31,80,31,202,31,131,31,102,31,84,31,55,31,93,31,80,31,17,31,200,31,191,31,191,30,226,31,178,31,242,31,224,31,196,31,196,30,85,31,115,31,132,31,47,31,75,31,227,31,168,31,150,31,221,31,130,31,250,31,250,30,250,29,144,31,8,31,215,31,8,31,120,31,120,30,192,31,42,31,103,31,111,31,236,31,121,31,121,30,90,31,102,31,153,31,167,31,14,31,191,31,191,30,197,31,197,30,194,31,62,31,62,30,62,29,35,31,8,31,21,31,21,30,203,31,41,31,87,31,87,30,87,29,87,28,19,31,161,31,161,30,129,31,190,31,47,31,47,30,211,31,211,30,172,31,172,30,17,31,66,31,234,31,81,31,220,31,165,31,111,31,111,30,111,29,199,31,159,31,18,31,244,31,244,30,249,31,249,30,211,31,75,31,193,31,193,30,189,31,137,31,137,30,30,31,217,31,107,31,206,31,206,30,36,31,113,31,187,31,187,30,187,29,114,31,223,31,223,31,158,31,158,30,158,29,232,31,191,31,191,30,122,31,144,31,218,31,178,31,28,31,34,31,69,31,69,30,23,31,144,31,55,31,24,31,122,31,122,30,13,31,134,31,134,30,158,31,103,31,217,31,67,31,67,30,67,29,179,31,239,31,239,30,239,29,68,31,12,31,146,31,216,31,222,31,38,31,150,31,227,31,111,31,36,31,119,31,221,31,120,31,101,31,136,31,1,31,163,31,171,31,169,31,64,31,60,31,133,31,167,31,167,30,167,29,226,31,143,31,143,30,143,29,77,31,77,30,187,31,121,31,121,30,207,31,200,31,200,30,194,31,164,31,164,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
