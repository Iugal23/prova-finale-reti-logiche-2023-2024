-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_210 is
end project_tb_210;

architecture project_tb_arch_210 of project_tb_210 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1012;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (42,0,0,0,68,0,60,0,96,0,0,0,42,0,119,0,231,0,0,0,100,0,0,0,0,0,205,0,213,0,16,0,0,0,122,0,3,0,27,0,78,0,171,0,0,0,0,0,187,0,155,0,73,0,177,0,0,0,171,0,72,0,184,0,103,0,160,0,0,0,93,0,0,0,126,0,99,0,0,0,59,0,19,0,0,0,0,0,0,0,250,0,88,0,91,0,209,0,208,0,37,0,171,0,62,0,188,0,0,0,60,0,0,0,107,0,158,0,185,0,0,0,0,0,53,0,210,0,238,0,52,0,69,0,13,0,59,0,191,0,227,0,45,0,138,0,98,0,132,0,0,0,0,0,200,0,0,0,215,0,0,0,61,0,10,0,87,0,0,0,29,0,36,0,230,0,23,0,88,0,0,0,255,0,0,0,167,0,0,0,0,0,39,0,71,0,0,0,0,0,205,0,79,0,216,0,0,0,135,0,140,0,126,0,240,0,179,0,0,0,67,0,76,0,63,0,152,0,211,0,40,0,112,0,95,0,0,0,183,0,149,0,224,0,195,0,0,0,36,0,148,0,213,0,177,0,212,0,0,0,230,0,28,0,67,0,0,0,0,0,2,0,73,0,0,0,160,0,112,0,0,0,27,0,48,0,0,0,120,0,177,0,163,0,104,0,60,0,119,0,65,0,201,0,233,0,0,0,178,0,0,0,154,0,0,0,0,0,103,0,255,0,243,0,190,0,227,0,132,0,1,0,212,0,182,0,33,0,49,0,0,0,138,0,72,0,231,0,222,0,59,0,252,0,107,0,199,0,52,0,167,0,34,0,6,0,137,0,111,0,192,0,248,0,85,0,88,0,166,0,51,0,0,0,6,0,4,0,1,0,116,0,177,0,15,0,0,0,0,0,2,0,205,0,253,0,133,0,27,0,131,0,20,0,160,0,99,0,138,0,129,0,111,0,218,0,251,0,214,0,235,0,118,0,0,0,71,0,86,0,0,0,86,0,216,0,126,0,43,0,111,0,0,0,6,0,3,0,0,0,171,0,0,0,245,0,29,0,80,0,52,0,0,0,0,0,0,0,1,0,131,0,144,0,63,0,78,0,0,0,184,0,225,0,239,0,225,0,35,0,45,0,94,0,66,0,12,0,171,0,0,0,0,0,13,0,157,0,0,0,0,0,0,0,190,0,148,0,0,0,0,0,215,0,25,0,81,0,118,0,62,0,71,0,0,0,0,0,68,0,58,0,57,0,155,0,118,0,17,0,167,0,91,0,208,0,0,0,228,0,0,0,0,0,112,0,0,0,233,0,188,0,77,0,0,0,193,0,17,0,68,0,182,0,78,0,0,0,135,0,98,0,97,0,39,0,32,0,204,0,207,0,7,0,27,0,0,0,158,0,184,0,0,0,184,0,0,0,111,0,28,0,233,0,77,0,240,0,129,0,133,0,52,0,0,0,138,0,0,0,79,0,54,0,88,0,63,0,213,0,78,0,0,0,0,0,204,0,0,0,138,0,12,0,0,0,57,0,131,0,109,0,131,0,46,0,118,0,218,0,173,0,136,0,146,0,215,0,187,0,25,0,124,0,225,0,191,0,20,0,155,0,0,0,120,0,141,0,2,0,207,0,224,0,158,0,54,0,217,0,194,0,51,0,24,0,0,0,148,0,203,0,101,0,0,0,207,0,149,0,9,0,12,0,110,0,80,0,213,0,78,0,61,0,0,0,0,0,63,0,173,0,161,0,170,0,132,0,176,0,169,0,248,0,0,0,229,0,101,0,174,0,104,0,130,0,0,0,161,0,128,0,6,0,17,0,12,0,0,0,141,0,172,0,78,0,20,0,63,0,70,0,118,0,0,0,35,0,13,0,214,0,0,0,156,0,240,0,85,0,175,0,88,0,224,0,126,0,6,0,173,0,161,0,0,0,207,0,140,0,3,0,145,0,71,0,0,0,0,0,140,0,11,0,250,0,73,0,157,0,2,0,245,0,5,0,241,0,208,0,0,0,105,0,228,0,240,0,202,0,97,0,242,0,0,0,95,0,121,0,179,0,83,0,75,0,185,0,137,0,47,0,48,0,0,0,0,0,64,0,231,0,55,0,69,0,254,0,143,0,42,0,0,0,11,0,0,0,132,0,66,0,170,0,120,0,173,0,71,0,214,0,3,0,218,0,0,0,250,0,128,0,16,0,130,0,0,0,180,0,175,0,0,0,190,0,57,0,78,0,196,0,0,0,68,0,250,0,0,0,0,0,89,0,0,0,86,0,0,0,97,0,89,0,208,0,240,0,0,0,85,0,244,0,60,0,0,0,0,0,245,0,0,0,92,0,0,0,199,0,88,0,228,0,189,0,152,0,171,0,0,0,191,0,0,0,33,0,233,0,85,0,0,0,248,0,20,0,0,0,55,0,250,0,212,0,86,0,31,0,233,0,0,0,167,0,231,0,100,0,123,0,21,0,241,0,113,0,0,0,50,0,107,0,252,0,254,0,132,0,76,0,0,0,0,0,164,0,118,0,0,0,48,0,177,0,124,0,5,0,248,0,251,0,123,0,247,0,199,0,0,0,87,0,38,0,126,0,38,0,43,0,121,0,0,0,54,0,122,0,162,0,89,0,137,0,69,0,0,0,70,0,66,0,27,0,129,0,0,0,203,0,174,0,209,0,196,0,129,0,118,0,0,0,215,0,20,0,72,0,189,0,29,0,27,0,121,0,4,0,0,0,47,0,255,0,138,0,159,0,211,0,164,0,0,0,237,0,59,0,206,0,120,0,0,0,232,0,104,0,0,0,235,0,242,0,250,0,221,0,70,0,93,0,212,0,246,0,123,0,141,0,241,0,249,0,36,0,19,0,105,0,171,0,253,0,208,0,225,0,220,0,0,0,0,0,0,0,4,0,182,0,0,0,255,0,233,0,19,0,71,0,117,0,39,0,254,0,25,0,0,0,169,0,0,0,74,0,0,0,55,0,31,0,8,0,0,0,14,0,10,0,120,0,75,0,0,0,0,0,125,0,10,0,50,0,0,0,204,0,212,0,210,0,57,0,138,0,224,0,90,0,5,0,117,0,253,0,248,0,176,0,39,0,52,0,105,0,168,0,194,0,217,0,116,0,0,0,128,0,0,0,202,0,95,0,216,0,223,0,125,0,170,0,28,0,221,0,197,0,211,0,56,0,87,0,18,0,164,0,249,0,0,0,169,0,110,0,191,0,145,0,0,0,103,0,162,0,129,0,85,0,6,0,95,0,225,0,130,0,112,0,0,0,159,0,251,0,0,0,0,0,1,0,191,0,0,0,78,0,50,0,29,0,211,0,77,0,136,0,0,0,0,0,209,0,158,0,71,0,188,0,2,0,125,0,0,0,255,0,187,0,27,0,96,0,131,0,27,0,97,0,81,0,24,0,0,0,0,0,71,0,0,0,56,0,231,0,68,0,142,0,247,0,0,0,0,0,175,0,12,0,176,0,205,0,89,0,55,0,237,0,0,0,82,0,228,0,0,0,212,0,85,0,17,0,37,0,85,0,175,0,156,0,162,0,41,0,0,0,23,0,28,0,75,0,159,0,233,0,203,0,0,0,0,0,182,0,43,0,232,0,235,0,0,0,61,0,86,0,66,0,29,0,70,0,0,0,24,0,0,0,191,0,0,0,107,0,125,0,173,0,0,0,217,0,137,0,236,0,187,0,161,0,0,0,237,0,206,0,0,0,227,0,236,0,80,0,20,0,47,0,0,0,88,0,0,0,29,0,68,0,0,0,67,0,88,0,0,0,0,0,124,0,0,0,242,0,191,0,39,0,0,0,0,0,3,0,123,0,44,0,98,0,120,0,236,0,22,0,192,0,0,0,104,0,96,0,0,0,236,0,242,0,157,0,80,0,238,0,245,0,165,0,39,0,80,0,139,0,0,0,8,0,232,0,247,0,232,0,243,0,105,0,0,0,0,0,92,0,184,0,64,0,0,0,93,0,118,0,177,0,6,0,235,0,22,0,0,0,89,0,206,0,23,0,59,0,156,0,116,0,0,0,224,0,255,0,0,0,118,0,81,0,52,0,227,0,48,0,165,0,109,0,214,0,9,0,0,0,0,0,95,0,253,0,50,0,133,0,7,0,7,0,2,0,133,0,239,0,0,0,0,0,187,0,0,0,106,0,0,0,0,0,162,0,108,0,0,0,50,0,126,0,34,0,0,0,85,0,224,0,0,0,175,0,69,0,88,0,0,0,253,0,56,0,77,0,11,0,117,0,111,0,0,0,189,0,90,0,179,0,153,0,136,0,127,0,234,0,0,0,89,0,92,0,0,0,110,0,179,0,78,0,11,0,19,0,51,0,0,0,208,0,28,0,239,0,4,0,0,0,56,0,0,0,155,0,0,0,88,0,113,0,65,0,68,0,0,0,91,0,39,0,0,0,6,0,206,0,157,0,107,0,48,0,177,0,117,0,231,0,56,0,175,0,144,0,44,0,0,0,202,0,251,0,0,0,0,0,4,0,23,0,251,0,118,0,0,0,201,0,243,0,84,0,0,0,133,0,98,0,7,0);
signal scenario_full  : scenario_type := (42,31,42,30,68,31,60,31,96,31,96,30,42,31,119,31,231,31,231,30,100,31,100,30,100,29,205,31,213,31,16,31,16,30,122,31,3,31,27,31,78,31,171,31,171,30,171,29,187,31,155,31,73,31,177,31,177,30,171,31,72,31,184,31,103,31,160,31,160,30,93,31,93,30,126,31,99,31,99,30,59,31,19,31,19,30,19,29,19,28,250,31,88,31,91,31,209,31,208,31,37,31,171,31,62,31,188,31,188,30,60,31,60,30,107,31,158,31,185,31,185,30,185,29,53,31,210,31,238,31,52,31,69,31,13,31,59,31,191,31,227,31,45,31,138,31,98,31,132,31,132,30,132,29,200,31,200,30,215,31,215,30,61,31,10,31,87,31,87,30,29,31,36,31,230,31,23,31,88,31,88,30,255,31,255,30,167,31,167,30,167,29,39,31,71,31,71,30,71,29,205,31,79,31,216,31,216,30,135,31,140,31,126,31,240,31,179,31,179,30,67,31,76,31,63,31,152,31,211,31,40,31,112,31,95,31,95,30,183,31,149,31,224,31,195,31,195,30,36,31,148,31,213,31,177,31,212,31,212,30,230,31,28,31,67,31,67,30,67,29,2,31,73,31,73,30,160,31,112,31,112,30,27,31,48,31,48,30,120,31,177,31,163,31,104,31,60,31,119,31,65,31,201,31,233,31,233,30,178,31,178,30,154,31,154,30,154,29,103,31,255,31,243,31,190,31,227,31,132,31,1,31,212,31,182,31,33,31,49,31,49,30,138,31,72,31,231,31,222,31,59,31,252,31,107,31,199,31,52,31,167,31,34,31,6,31,137,31,111,31,192,31,248,31,85,31,88,31,166,31,51,31,51,30,6,31,4,31,1,31,116,31,177,31,15,31,15,30,15,29,2,31,205,31,253,31,133,31,27,31,131,31,20,31,160,31,99,31,138,31,129,31,111,31,218,31,251,31,214,31,235,31,118,31,118,30,71,31,86,31,86,30,86,31,216,31,126,31,43,31,111,31,111,30,6,31,3,31,3,30,171,31,171,30,245,31,29,31,80,31,52,31,52,30,52,29,52,28,1,31,131,31,144,31,63,31,78,31,78,30,184,31,225,31,239,31,225,31,35,31,45,31,94,31,66,31,12,31,171,31,171,30,171,29,13,31,157,31,157,30,157,29,157,28,190,31,148,31,148,30,148,29,215,31,25,31,81,31,118,31,62,31,71,31,71,30,71,29,68,31,58,31,57,31,155,31,118,31,17,31,167,31,91,31,208,31,208,30,228,31,228,30,228,29,112,31,112,30,233,31,188,31,77,31,77,30,193,31,17,31,68,31,182,31,78,31,78,30,135,31,98,31,97,31,39,31,32,31,204,31,207,31,7,31,27,31,27,30,158,31,184,31,184,30,184,31,184,30,111,31,28,31,233,31,77,31,240,31,129,31,133,31,52,31,52,30,138,31,138,30,79,31,54,31,88,31,63,31,213,31,78,31,78,30,78,29,204,31,204,30,138,31,12,31,12,30,57,31,131,31,109,31,131,31,46,31,118,31,218,31,173,31,136,31,146,31,215,31,187,31,25,31,124,31,225,31,191,31,20,31,155,31,155,30,120,31,141,31,2,31,207,31,224,31,158,31,54,31,217,31,194,31,51,31,24,31,24,30,148,31,203,31,101,31,101,30,207,31,149,31,9,31,12,31,110,31,80,31,213,31,78,31,61,31,61,30,61,29,63,31,173,31,161,31,170,31,132,31,176,31,169,31,248,31,248,30,229,31,101,31,174,31,104,31,130,31,130,30,161,31,128,31,6,31,17,31,12,31,12,30,141,31,172,31,78,31,20,31,63,31,70,31,118,31,118,30,35,31,13,31,214,31,214,30,156,31,240,31,85,31,175,31,88,31,224,31,126,31,6,31,173,31,161,31,161,30,207,31,140,31,3,31,145,31,71,31,71,30,71,29,140,31,11,31,250,31,73,31,157,31,2,31,245,31,5,31,241,31,208,31,208,30,105,31,228,31,240,31,202,31,97,31,242,31,242,30,95,31,121,31,179,31,83,31,75,31,185,31,137,31,47,31,48,31,48,30,48,29,64,31,231,31,55,31,69,31,254,31,143,31,42,31,42,30,11,31,11,30,132,31,66,31,170,31,120,31,173,31,71,31,214,31,3,31,218,31,218,30,250,31,128,31,16,31,130,31,130,30,180,31,175,31,175,30,190,31,57,31,78,31,196,31,196,30,68,31,250,31,250,30,250,29,89,31,89,30,86,31,86,30,97,31,89,31,208,31,240,31,240,30,85,31,244,31,60,31,60,30,60,29,245,31,245,30,92,31,92,30,199,31,88,31,228,31,189,31,152,31,171,31,171,30,191,31,191,30,33,31,233,31,85,31,85,30,248,31,20,31,20,30,55,31,250,31,212,31,86,31,31,31,233,31,233,30,167,31,231,31,100,31,123,31,21,31,241,31,113,31,113,30,50,31,107,31,252,31,254,31,132,31,76,31,76,30,76,29,164,31,118,31,118,30,48,31,177,31,124,31,5,31,248,31,251,31,123,31,247,31,199,31,199,30,87,31,38,31,126,31,38,31,43,31,121,31,121,30,54,31,122,31,162,31,89,31,137,31,69,31,69,30,70,31,66,31,27,31,129,31,129,30,203,31,174,31,209,31,196,31,129,31,118,31,118,30,215,31,20,31,72,31,189,31,29,31,27,31,121,31,4,31,4,30,47,31,255,31,138,31,159,31,211,31,164,31,164,30,237,31,59,31,206,31,120,31,120,30,232,31,104,31,104,30,235,31,242,31,250,31,221,31,70,31,93,31,212,31,246,31,123,31,141,31,241,31,249,31,36,31,19,31,105,31,171,31,253,31,208,31,225,31,220,31,220,30,220,29,220,28,4,31,182,31,182,30,255,31,233,31,19,31,71,31,117,31,39,31,254,31,25,31,25,30,169,31,169,30,74,31,74,30,55,31,31,31,8,31,8,30,14,31,10,31,120,31,75,31,75,30,75,29,125,31,10,31,50,31,50,30,204,31,212,31,210,31,57,31,138,31,224,31,90,31,5,31,117,31,253,31,248,31,176,31,39,31,52,31,105,31,168,31,194,31,217,31,116,31,116,30,128,31,128,30,202,31,95,31,216,31,223,31,125,31,170,31,28,31,221,31,197,31,211,31,56,31,87,31,18,31,164,31,249,31,249,30,169,31,110,31,191,31,145,31,145,30,103,31,162,31,129,31,85,31,6,31,95,31,225,31,130,31,112,31,112,30,159,31,251,31,251,30,251,29,1,31,191,31,191,30,78,31,50,31,29,31,211,31,77,31,136,31,136,30,136,29,209,31,158,31,71,31,188,31,2,31,125,31,125,30,255,31,187,31,27,31,96,31,131,31,27,31,97,31,81,31,24,31,24,30,24,29,71,31,71,30,56,31,231,31,68,31,142,31,247,31,247,30,247,29,175,31,12,31,176,31,205,31,89,31,55,31,237,31,237,30,82,31,228,31,228,30,212,31,85,31,17,31,37,31,85,31,175,31,156,31,162,31,41,31,41,30,23,31,28,31,75,31,159,31,233,31,203,31,203,30,203,29,182,31,43,31,232,31,235,31,235,30,61,31,86,31,66,31,29,31,70,31,70,30,24,31,24,30,191,31,191,30,107,31,125,31,173,31,173,30,217,31,137,31,236,31,187,31,161,31,161,30,237,31,206,31,206,30,227,31,236,31,80,31,20,31,47,31,47,30,88,31,88,30,29,31,68,31,68,30,67,31,88,31,88,30,88,29,124,31,124,30,242,31,191,31,39,31,39,30,39,29,3,31,123,31,44,31,98,31,120,31,236,31,22,31,192,31,192,30,104,31,96,31,96,30,236,31,242,31,157,31,80,31,238,31,245,31,165,31,39,31,80,31,139,31,139,30,8,31,232,31,247,31,232,31,243,31,105,31,105,30,105,29,92,31,184,31,64,31,64,30,93,31,118,31,177,31,6,31,235,31,22,31,22,30,89,31,206,31,23,31,59,31,156,31,116,31,116,30,224,31,255,31,255,30,118,31,81,31,52,31,227,31,48,31,165,31,109,31,214,31,9,31,9,30,9,29,95,31,253,31,50,31,133,31,7,31,7,31,2,31,133,31,239,31,239,30,239,29,187,31,187,30,106,31,106,30,106,29,162,31,108,31,108,30,50,31,126,31,34,31,34,30,85,31,224,31,224,30,175,31,69,31,88,31,88,30,253,31,56,31,77,31,11,31,117,31,111,31,111,30,189,31,90,31,179,31,153,31,136,31,127,31,234,31,234,30,89,31,92,31,92,30,110,31,179,31,78,31,11,31,19,31,51,31,51,30,208,31,28,31,239,31,4,31,4,30,56,31,56,30,155,31,155,30,88,31,113,31,65,31,68,31,68,30,91,31,39,31,39,30,6,31,206,31,157,31,107,31,48,31,177,31,117,31,231,31,56,31,175,31,144,31,44,31,44,30,202,31,251,31,251,30,251,29,4,31,23,31,251,31,118,31,118,30,201,31,243,31,84,31,84,30,133,31,98,31,7,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
