-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_673 is
end project_tb_673;

architecture project_tb_arch_673 of project_tb_673 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 706;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,35,0,178,0,57,0,183,0,0,0,212,0,249,0,0,0,182,0,100,0,41,0,0,0,205,0,240,0,133,0,126,0,58,0,19,0,100,0,28,0,0,0,0,0,51,0,228,0,53,0,115,0,68,0,0,0,5,0,136,0,88,0,195,0,21,0,84,0,83,0,102,0,54,0,215,0,133,0,33,0,123,0,140,0,17,0,0,0,0,0,68,0,0,0,55,0,114,0,180,0,49,0,53,0,241,0,169,0,58,0,0,0,231,0,191,0,231,0,46,0,242,0,26,0,25,0,130,0,0,0,205,0,24,0,131,0,251,0,122,0,18,0,48,0,82,0,232,0,115,0,0,0,90,0,0,0,181,0,215,0,29,0,5,0,0,0,68,0,175,0,0,0,85,0,189,0,148,0,13,0,41,0,178,0,0,0,62,0,194,0,215,0,0,0,10,0,126,0,204,0,0,0,127,0,187,0,133,0,95,0,114,0,149,0,11,0,127,0,0,0,204,0,62,0,39,0,203,0,135,0,114,0,132,0,181,0,0,0,97,0,178,0,137,0,0,0,157,0,238,0,0,0,23,0,42,0,208,0,43,0,247,0,222,0,190,0,181,0,162,0,119,0,82,0,31,0,34,0,0,0,138,0,213,0,123,0,0,0,51,0,11,0,0,0,153,0,106,0,0,0,0,0,5,0,0,0,0,0,0,0,205,0,1,0,154,0,230,0,0,0,207,0,248,0,3,0,195,0,140,0,0,0,212,0,0,0,159,0,69,0,147,0,0,0,0,0,0,0,121,0,211,0,175,0,68,0,87,0,0,0,0,0,150,0,43,0,36,0,0,0,211,0,211,0,98,0,242,0,147,0,124,0,0,0,144,0,0,0,66,0,67,0,19,0,182,0,190,0,0,0,179,0,40,0,63,0,85,0,165,0,85,0,13,0,11,0,176,0,162,0,226,0,222,0,102,0,105,0,0,0,184,0,119,0,0,0,132,0,188,0,60,0,32,0,174,0,194,0,35,0,218,0,0,0,184,0,41,0,101,0,122,0,88,0,100,0,149,0,198,0,0,0,0,0,87,0,182,0,138,0,92,0,167,0,0,0,0,0,0,0,15,0,5,0,236,0,88,0,192,0,253,0,245,0,0,0,135,0,149,0,158,0,35,0,251,0,165,0,42,0,123,0,0,0,119,0,0,0,79,0,244,0,246,0,239,0,117,0,110,0,213,0,0,0,0,0,108,0,59,0,114,0,205,0,146,0,56,0,14,0,0,0,0,0,200,0,193,0,85,0,136,0,0,0,122,0,0,0,206,0,192,0,202,0,0,0,169,0,122,0,93,0,47,0,222,0,4,0,238,0,159,0,125,0,77,0,0,0,176,0,233,0,0,0,133,0,74,0,133,0,212,0,137,0,94,0,183,0,0,0,89,0,198,0,4,0,0,0,139,0,227,0,64,0,233,0,0,0,230,0,88,0,222,0,207,0,157,0,252,0,87,0,210,0,0,0,84,0,0,0,244,0,85,0,237,0,26,0,66,0,0,0,142,0,0,0,1,0,66,0,0,0,225,0,174,0,170,0,4,0,206,0,71,0,122,0,225,0,0,0,183,0,7,0,7,0,213,0,127,0,0,0,244,0,177,0,187,0,244,0,228,0,0,0,192,0,0,0,176,0,240,0,3,0,206,0,69,0,247,0,0,0,0,0,0,0,242,0,200,0,214,0,248,0,215,0,26,0,123,0,10,0,148,0,247,0,29,0,0,0,81,0,27,0,40,0,166,0,184,0,80,0,47,0,0,0,246,0,145,0,166,0,23,0,138,0,244,0,91,0,12,0,0,0,225,0,87,0,12,0,0,0,228,0,0,0,253,0,86,0,244,0,153,0,0,0,170,0,0,0,160,0,31,0,67,0,242,0,250,0,36,0,52,0,156,0,79,0,209,0,166,0,0,0,20,0,0,0,57,0,0,0,111,0,72,0,81,0,175,0,236,0,246,0,48,0,88,0,230,0,12,0,245,0,215,0,0,0,0,0,116,0,49,0,130,0,0,0,39,0,65,0,224,0,0,0,242,0,0,0,36,0,29,0,237,0,131,0,119,0,218,0,161,0,87,0,0,0,0,0,146,0,48,0,91,0,247,0,149,0,51,0,122,0,234,0,89,0,170,0,201,0,0,0,168,0,175,0,205,0,111,0,0,0,0,0,249,0,151,0,219,0,4,0,215,0,53,0,0,0,217,0,31,0,248,0,56,0,206,0,167,0,0,0,45,0,178,0,192,0,38,0,54,0,106,0,73,0,71,0,118,0,105,0,0,0,150,0,158,0,0,0,224,0,139,0,239,0,81,0,11,0,139,0,8,0,239,0,235,0,190,0,0,0,88,0,227,0,212,0,47,0,0,0,205,0,120,0,12,0,52,0,250,0,124,0,205,0,219,0,128,0,248,0,65,0,122,0,96,0,160,0,0,0,120,0,23,0,67,0,0,0,245,0,0,0,0,0,239,0,25,0,195,0,0,0,88,0,177,0,0,0,142,0,165,0,0,0,35,0,0,0,28,0,74,0,24,0,226,0,57,0,53,0,232,0,82,0,175,0,108,0,0,0,0,0,45,0,89,0,80,0,102,0,141,0,0,0,0,0,237,0,13,0,12,0,253,0,75,0,205,0,213,0,245,0,203,0,91,0,106,0,248,0,154,0,21,0,0,0,0,0,93,0,5,0,0,0,246,0,147,0,0,0,0,0,171,0,0,0,114,0,0,0,13,0,203,0,251,0,11,0,158,0,0,0,222,0,0,0,184,0,245,0,138,0,0,0,160,0,20,0,0,0,134,0,33,0,124,0,106,0,0,0,239,0,78,0,37,0,216,0,23,0,0,0,192,0,122,0,234,0,0,0,33,0,7,0,108,0,114,0,0,0,164,0,126,0,0,0,163,0,0,0,236,0,237,0,141,0,144,0,58,0,60,0,165,0,237,0,169,0,46,0,89,0,56,0,0,0,237,0,4,0,152,0,19,0,94,0,200,0,199,0,232,0,0,0,65,0,0,0,99,0,47,0,0,0,121,0,150,0,0,0,118,0,83,0,231,0,168,0,21,0,35,0,61,0,198,0,93,0,146,0,94,0,163,0,212,0,21,0,126,0,98,0,245,0,0,0,98,0,0,0,47,0,76,0,182,0);
signal scenario_full  : scenario_type := (0,0,35,31,178,31,57,31,183,31,183,30,212,31,249,31,249,30,182,31,100,31,41,31,41,30,205,31,240,31,133,31,126,31,58,31,19,31,100,31,28,31,28,30,28,29,51,31,228,31,53,31,115,31,68,31,68,30,5,31,136,31,88,31,195,31,21,31,84,31,83,31,102,31,54,31,215,31,133,31,33,31,123,31,140,31,17,31,17,30,17,29,68,31,68,30,55,31,114,31,180,31,49,31,53,31,241,31,169,31,58,31,58,30,231,31,191,31,231,31,46,31,242,31,26,31,25,31,130,31,130,30,205,31,24,31,131,31,251,31,122,31,18,31,48,31,82,31,232,31,115,31,115,30,90,31,90,30,181,31,215,31,29,31,5,31,5,30,68,31,175,31,175,30,85,31,189,31,148,31,13,31,41,31,178,31,178,30,62,31,194,31,215,31,215,30,10,31,126,31,204,31,204,30,127,31,187,31,133,31,95,31,114,31,149,31,11,31,127,31,127,30,204,31,62,31,39,31,203,31,135,31,114,31,132,31,181,31,181,30,97,31,178,31,137,31,137,30,157,31,238,31,238,30,23,31,42,31,208,31,43,31,247,31,222,31,190,31,181,31,162,31,119,31,82,31,31,31,34,31,34,30,138,31,213,31,123,31,123,30,51,31,11,31,11,30,153,31,106,31,106,30,106,29,5,31,5,30,5,29,5,28,205,31,1,31,154,31,230,31,230,30,207,31,248,31,3,31,195,31,140,31,140,30,212,31,212,30,159,31,69,31,147,31,147,30,147,29,147,28,121,31,211,31,175,31,68,31,87,31,87,30,87,29,150,31,43,31,36,31,36,30,211,31,211,31,98,31,242,31,147,31,124,31,124,30,144,31,144,30,66,31,67,31,19,31,182,31,190,31,190,30,179,31,40,31,63,31,85,31,165,31,85,31,13,31,11,31,176,31,162,31,226,31,222,31,102,31,105,31,105,30,184,31,119,31,119,30,132,31,188,31,60,31,32,31,174,31,194,31,35,31,218,31,218,30,184,31,41,31,101,31,122,31,88,31,100,31,149,31,198,31,198,30,198,29,87,31,182,31,138,31,92,31,167,31,167,30,167,29,167,28,15,31,5,31,236,31,88,31,192,31,253,31,245,31,245,30,135,31,149,31,158,31,35,31,251,31,165,31,42,31,123,31,123,30,119,31,119,30,79,31,244,31,246,31,239,31,117,31,110,31,213,31,213,30,213,29,108,31,59,31,114,31,205,31,146,31,56,31,14,31,14,30,14,29,200,31,193,31,85,31,136,31,136,30,122,31,122,30,206,31,192,31,202,31,202,30,169,31,122,31,93,31,47,31,222,31,4,31,238,31,159,31,125,31,77,31,77,30,176,31,233,31,233,30,133,31,74,31,133,31,212,31,137,31,94,31,183,31,183,30,89,31,198,31,4,31,4,30,139,31,227,31,64,31,233,31,233,30,230,31,88,31,222,31,207,31,157,31,252,31,87,31,210,31,210,30,84,31,84,30,244,31,85,31,237,31,26,31,66,31,66,30,142,31,142,30,1,31,66,31,66,30,225,31,174,31,170,31,4,31,206,31,71,31,122,31,225,31,225,30,183,31,7,31,7,31,213,31,127,31,127,30,244,31,177,31,187,31,244,31,228,31,228,30,192,31,192,30,176,31,240,31,3,31,206,31,69,31,247,31,247,30,247,29,247,28,242,31,200,31,214,31,248,31,215,31,26,31,123,31,10,31,148,31,247,31,29,31,29,30,81,31,27,31,40,31,166,31,184,31,80,31,47,31,47,30,246,31,145,31,166,31,23,31,138,31,244,31,91,31,12,31,12,30,225,31,87,31,12,31,12,30,228,31,228,30,253,31,86,31,244,31,153,31,153,30,170,31,170,30,160,31,31,31,67,31,242,31,250,31,36,31,52,31,156,31,79,31,209,31,166,31,166,30,20,31,20,30,57,31,57,30,111,31,72,31,81,31,175,31,236,31,246,31,48,31,88,31,230,31,12,31,245,31,215,31,215,30,215,29,116,31,49,31,130,31,130,30,39,31,65,31,224,31,224,30,242,31,242,30,36,31,29,31,237,31,131,31,119,31,218,31,161,31,87,31,87,30,87,29,146,31,48,31,91,31,247,31,149,31,51,31,122,31,234,31,89,31,170,31,201,31,201,30,168,31,175,31,205,31,111,31,111,30,111,29,249,31,151,31,219,31,4,31,215,31,53,31,53,30,217,31,31,31,248,31,56,31,206,31,167,31,167,30,45,31,178,31,192,31,38,31,54,31,106,31,73,31,71,31,118,31,105,31,105,30,150,31,158,31,158,30,224,31,139,31,239,31,81,31,11,31,139,31,8,31,239,31,235,31,190,31,190,30,88,31,227,31,212,31,47,31,47,30,205,31,120,31,12,31,52,31,250,31,124,31,205,31,219,31,128,31,248,31,65,31,122,31,96,31,160,31,160,30,120,31,23,31,67,31,67,30,245,31,245,30,245,29,239,31,25,31,195,31,195,30,88,31,177,31,177,30,142,31,165,31,165,30,35,31,35,30,28,31,74,31,24,31,226,31,57,31,53,31,232,31,82,31,175,31,108,31,108,30,108,29,45,31,89,31,80,31,102,31,141,31,141,30,141,29,237,31,13,31,12,31,253,31,75,31,205,31,213,31,245,31,203,31,91,31,106,31,248,31,154,31,21,31,21,30,21,29,93,31,5,31,5,30,246,31,147,31,147,30,147,29,171,31,171,30,114,31,114,30,13,31,203,31,251,31,11,31,158,31,158,30,222,31,222,30,184,31,245,31,138,31,138,30,160,31,20,31,20,30,134,31,33,31,124,31,106,31,106,30,239,31,78,31,37,31,216,31,23,31,23,30,192,31,122,31,234,31,234,30,33,31,7,31,108,31,114,31,114,30,164,31,126,31,126,30,163,31,163,30,236,31,237,31,141,31,144,31,58,31,60,31,165,31,237,31,169,31,46,31,89,31,56,31,56,30,237,31,4,31,152,31,19,31,94,31,200,31,199,31,232,31,232,30,65,31,65,30,99,31,47,31,47,30,121,31,150,31,150,30,118,31,83,31,231,31,168,31,21,31,35,31,61,31,198,31,93,31,146,31,94,31,163,31,212,31,21,31,126,31,98,31,245,31,245,30,98,31,98,30,47,31,76,31,182,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
