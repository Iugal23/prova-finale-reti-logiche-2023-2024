-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 996;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,114,0,0,0,0,0,46,0,35,0,179,0,11,0,129,0,84,0,174,0,0,0,182,0,28,0,174,0,43,0,178,0,64,0,173,0,0,0,83,0,197,0,0,0,201,0,138,0,219,0,128,0,137,0,152,0,171,0,216,0,238,0,10,0,0,0,241,0,92,0,44,0,109,0,89,0,68,0,60,0,41,0,63,0,90,0,142,0,160,0,80,0,184,0,66,0,15,0,252,0,139,0,73,0,212,0,45,0,231,0,52,0,0,0,237,0,0,0,47,0,160,0,69,0,46,0,60,0,0,0,66,0,0,0,108,0,151,0,169,0,43,0,217,0,9,0,230,0,233,0,253,0,147,0,211,0,150,0,206,0,167,0,195,0,255,0,0,0,230,0,18,0,0,0,107,0,24,0,188,0,88,0,120,0,186,0,204,0,166,0,153,0,157,0,196,0,47,0,147,0,60,0,231,0,237,0,218,0,155,0,17,0,0,0,0,0,0,0,151,0,42,0,249,0,0,0,0,0,72,0,175,0,205,0,108,0,0,0,81,0,101,0,0,0,148,0,116,0,248,0,31,0,0,0,0,0,0,0,9,0,0,0,56,0,0,0,223,0,32,0,230,0,165,0,117,0,50,0,39,0,9,0,31,0,97,0,162,0,7,0,151,0,200,0,84,0,244,0,0,0,20,0,192,0,0,0,7,0,127,0,179,0,180,0,47,0,39,0,111,0,176,0,34,0,93,0,0,0,223,0,18,0,35,0,142,0,255,0,98,0,30,0,78,0,233,0,192,0,0,0,0,0,10,0,0,0,48,0,223,0,70,0,165,0,51,0,0,0,165,0,190,0,115,0,0,0,0,0,239,0,190,0,0,0,54,0,0,0,137,0,41,0,138,0,162,0,191,0,164,0,0,0,184,0,167,0,165,0,0,0,225,0,194,0,0,0,165,0,72,0,73,0,174,0,37,0,132,0,251,0,188,0,0,0,184,0,190,0,37,0,67,0,0,0,66,0,0,0,114,0,16,0,139,0,35,0,133,0,89,0,176,0,181,0,192,0,45,0,106,0,77,0,145,0,103,0,205,0,46,0,124,0,180,0,0,0,108,0,93,0,56,0,43,0,4,0,143,0,45,0,0,0,154,0,176,0,197,0,0,0,147,0,254,0,236,0,0,0,254,0,82,0,32,0,111,0,180,0,161,0,162,0,111,0,112,0,2,0,27,0,31,0,198,0,40,0,164,0,231,0,64,0,0,0,0,0,157,0,148,0,120,0,220,0,125,0,188,0,147,0,0,0,157,0,0,0,0,0,192,0,225,0,130,0,0,0,228,0,156,0,173,0,19,0,224,0,44,0,236,0,215,0,144,0,33,0,249,0,37,0,224,0,255,0,110,0,150,0,194,0,240,0,0,0,133,0,39,0,163,0,221,0,0,0,151,0,22,0,146,0,0,0,242,0,191,0,5,0,88,0,139,0,200,0,42,0,0,0,0,0,224,0,127,0,132,0,138,0,13,0,222,0,56,0,83,0,207,0,201,0,91,0,0,0,0,0,0,0,105,0,250,0,81,0,57,0,215,0,0,0,121,0,175,0,0,0,138,0,81,0,66,0,0,0,239,0,21,0,102,0,254,0,106,0,66,0,65,0,78,0,97,0,225,0,192,0,35,0,0,0,160,0,160,0,87,0,247,0,91,0,174,0,108,0,74,0,123,0,180,0,0,0,229,0,199,0,179,0,214,0,49,0,17,0,22,0,188,0,179,0,63,0,0,0,163,0,0,0,211,0,56,0,214,0,249,0,0,0,0,0,121,0,122,0,121,0,64,0,240,0,251,0,74,0,72,0,145,0,236,0,53,0,95,0,0,0,112,0,92,0,62,0,110,0,145,0,211,0,0,0,41,0,28,0,170,0,151,0,0,0,59,0,54,0,171,0,57,0,25,0,253,0,26,0,101,0,45,0,158,0,0,0,221,0,211,0,181,0,82,0,0,0,14,0,0,0,204,0,234,0,219,0,109,0,182,0,116,0,25,0,184,0,87,0,202,0,83,0,108,0,41,0,0,0,218,0,133,0,182,0,56,0,130,0,244,0,0,0,0,0,53,0,194,0,87,0,175,0,0,0,153,0,0,0,232,0,253,0,206,0,210,0,52,0,86,0,0,0,148,0,45,0,0,0,121,0,51,0,203,0,56,0,145,0,0,0,245,0,181,0,14,0,159,0,75,0,81,0,0,0,194,0,93,0,247,0,227,0,252,0,11,0,252,0,0,0,162,0,59,0,224,0,215,0,17,0,30,0,202,0,233,0,66,0,167,0,0,0,127,0,0,0,0,0,0,0,142,0,55,0,234,0,50,0,243,0,145,0,137,0,0,0,168,0,215,0,209,0,234,0,47,0,37,0,106,0,148,0,216,0,183,0,73,0,76,0,12,0,73,0,223,0,97,0,168,0,0,0,183,0,93,0,0,0,122,0,201,0,244,0,0,0,94,0,58,0,0,0,173,0,152,0,183,0,213,0,0,0,0,0,157,0,199,0,131,0,0,0,0,0,117,0,0,0,111,0,127,0,195,0,184,0,0,0,151,0,53,0,163,0,86,0,125,0,0,0,84,0,81,0,126,0,199,0,191,0,0,0,227,0,208,0,0,0,17,0,20,0,190,0,190,0,187,0,132,0,223,0,0,0,227,0,0,0,0,0,228,0,0,0,22,0,237,0,157,0,70,0,88,0,18,0,55,0,0,0,176,0,184,0,0,0,19,0,63,0,200,0,192,0,48,0,17,0,18,0,143,0,0,0,11,0,237,0,220,0,213,0,0,0,81,0,0,0,241,0,207,0,98,0,226,0,211,0,0,0,230,0,7,0,44,0,219,0,109,0,47,0,123,0,125,0,129,0,205,0,139,0,0,0,95,0,65,0,0,0,174,0,175,0,136,0,194,0,8,0,194,0,0,0,68,0,68,0,170,0,62,0,139,0,173,0,135,0,34,0,15,0,174,0,113,0,3,0,0,0,0,0,140,0,144,0,178,0,112,0,109,0,0,0,22,0,193,0,144,0,134,0,231,0,120,0,111,0,81,0,132,0,25,0,240,0,33,0,42,0,60,0,12,0,74,0,199,0,94,0,0,0,98,0,0,0,158,0,77,0,157,0,88,0,58,0,39,0,5,0,6,0,116,0,201,0,0,0,83,0,27,0,186,0,171,0,0,0,0,0,214,0,116,0,148,0,241,0,152,0,108,0,0,0,109,0,31,0,248,0,205,0,138,0,197,0,101,0,213,0,222,0,79,0,1,0,195,0,136,0,154,0,174,0,57,0,0,0,124,0,147,0,0,0,117,0,20,0,0,0,228,0,60,0,0,0,68,0,29,0,146,0,0,0,110,0,234,0,236,0,49,0,255,0,0,0,0,0,201,0,253,0,115,0,70,0,101,0,0,0,134,0,155,0,96,0,231,0,109,0,0,0,76,0,52,0,126,0,224,0,48,0,56,0,0,0,212,0,75,0,18,0,224,0,0,0,23,0,135,0,83,0,167,0,201,0,49,0,186,0,0,0,99,0,0,0,96,0,22,0,169,0,202,0,177,0,253,0,112,0,50,0,0,0,50,0,28,0,192,0,25,0,91,0,0,0,171,0,180,0,70,0,31,0,0,0,63,0,167,0,99,0,105,0,160,0,113,0,217,0,2,0,166,0,0,0,130,0,101,0,0,0,0,0,80,0,103,0,44,0,212,0,83,0,0,0,149,0,0,0,215,0,216,0,225,0,17,0,157,0,3,0,193,0,156,0,45,0,31,0,147,0,12,0,0,0,156,0,30,0,47,0,48,0,176,0,47,0,7,0,0,0,216,0,92,0,67,0,190,0,37,0,145,0,0,0,38,0,242,0,63,0,0,0,188,0,88,0,203,0,159,0,109,0,3,0,101,0,237,0,80,0,120,0,54,0,0,0,63,0,137,0,144,0,111,0,138,0,0,0,199,0,0,0,173,0,66,0,36,0,124,0,191,0,0,0,0,0,11,0,184,0,21,0,242,0,105,0,203,0,89,0,55,0,238,0,133,0,228,0,88,0,112,0,248,0,81,0,241,0,0,0,142,0,132,0,0,0,121,0,2,0,181,0,0,0,19,0,4,0,0,0,96,0,123,0,205,0,217,0,12,0,0,0,219,0,191,0,6,0,85,0,9,0,216,0,0,0,0,0,112,0,132,0,74,0,36,0,118,0,168,0,68,0,125,0,177,0,89,0,158,0,239,0,160,0,0,0,11,0,0,0,29,0,86,0,240,0,229,0,0,0,0,0,0,0,0,0,201,0,11,0,0,0,115,0,0,0,0,0,0,0,91,0,26,0,12,0,215,0,0,0,7,0,0,0,25,0,173,0,0,0,57,0,42,0,0,0,38,0,207,0,229,0,219,0,204,0,105,0,155,0,251,0,166,0,39,0,0,0,189,0,13,0,9,0,31,0,101,0,82,0,106,0);
signal scenario_full  : scenario_type := (0,0,114,31,114,30,114,29,46,31,35,31,179,31,11,31,129,31,84,31,174,31,174,30,182,31,28,31,174,31,43,31,178,31,64,31,173,31,173,30,83,31,197,31,197,30,201,31,138,31,219,31,128,31,137,31,152,31,171,31,216,31,238,31,10,31,10,30,241,31,92,31,44,31,109,31,89,31,68,31,60,31,41,31,63,31,90,31,142,31,160,31,80,31,184,31,66,31,15,31,252,31,139,31,73,31,212,31,45,31,231,31,52,31,52,30,237,31,237,30,47,31,160,31,69,31,46,31,60,31,60,30,66,31,66,30,108,31,151,31,169,31,43,31,217,31,9,31,230,31,233,31,253,31,147,31,211,31,150,31,206,31,167,31,195,31,255,31,255,30,230,31,18,31,18,30,107,31,24,31,188,31,88,31,120,31,186,31,204,31,166,31,153,31,157,31,196,31,47,31,147,31,60,31,231,31,237,31,218,31,155,31,17,31,17,30,17,29,17,28,151,31,42,31,249,31,249,30,249,29,72,31,175,31,205,31,108,31,108,30,81,31,101,31,101,30,148,31,116,31,248,31,31,31,31,30,31,29,31,28,9,31,9,30,56,31,56,30,223,31,32,31,230,31,165,31,117,31,50,31,39,31,9,31,31,31,97,31,162,31,7,31,151,31,200,31,84,31,244,31,244,30,20,31,192,31,192,30,7,31,127,31,179,31,180,31,47,31,39,31,111,31,176,31,34,31,93,31,93,30,223,31,18,31,35,31,142,31,255,31,98,31,30,31,78,31,233,31,192,31,192,30,192,29,10,31,10,30,48,31,223,31,70,31,165,31,51,31,51,30,165,31,190,31,115,31,115,30,115,29,239,31,190,31,190,30,54,31,54,30,137,31,41,31,138,31,162,31,191,31,164,31,164,30,184,31,167,31,165,31,165,30,225,31,194,31,194,30,165,31,72,31,73,31,174,31,37,31,132,31,251,31,188,31,188,30,184,31,190,31,37,31,67,31,67,30,66,31,66,30,114,31,16,31,139,31,35,31,133,31,89,31,176,31,181,31,192,31,45,31,106,31,77,31,145,31,103,31,205,31,46,31,124,31,180,31,180,30,108,31,93,31,56,31,43,31,4,31,143,31,45,31,45,30,154,31,176,31,197,31,197,30,147,31,254,31,236,31,236,30,254,31,82,31,32,31,111,31,180,31,161,31,162,31,111,31,112,31,2,31,27,31,31,31,198,31,40,31,164,31,231,31,64,31,64,30,64,29,157,31,148,31,120,31,220,31,125,31,188,31,147,31,147,30,157,31,157,30,157,29,192,31,225,31,130,31,130,30,228,31,156,31,173,31,19,31,224,31,44,31,236,31,215,31,144,31,33,31,249,31,37,31,224,31,255,31,110,31,150,31,194,31,240,31,240,30,133,31,39,31,163,31,221,31,221,30,151,31,22,31,146,31,146,30,242,31,191,31,5,31,88,31,139,31,200,31,42,31,42,30,42,29,224,31,127,31,132,31,138,31,13,31,222,31,56,31,83,31,207,31,201,31,91,31,91,30,91,29,91,28,105,31,250,31,81,31,57,31,215,31,215,30,121,31,175,31,175,30,138,31,81,31,66,31,66,30,239,31,21,31,102,31,254,31,106,31,66,31,65,31,78,31,97,31,225,31,192,31,35,31,35,30,160,31,160,31,87,31,247,31,91,31,174,31,108,31,74,31,123,31,180,31,180,30,229,31,199,31,179,31,214,31,49,31,17,31,22,31,188,31,179,31,63,31,63,30,163,31,163,30,211,31,56,31,214,31,249,31,249,30,249,29,121,31,122,31,121,31,64,31,240,31,251,31,74,31,72,31,145,31,236,31,53,31,95,31,95,30,112,31,92,31,62,31,110,31,145,31,211,31,211,30,41,31,28,31,170,31,151,31,151,30,59,31,54,31,171,31,57,31,25,31,253,31,26,31,101,31,45,31,158,31,158,30,221,31,211,31,181,31,82,31,82,30,14,31,14,30,204,31,234,31,219,31,109,31,182,31,116,31,25,31,184,31,87,31,202,31,83,31,108,31,41,31,41,30,218,31,133,31,182,31,56,31,130,31,244,31,244,30,244,29,53,31,194,31,87,31,175,31,175,30,153,31,153,30,232,31,253,31,206,31,210,31,52,31,86,31,86,30,148,31,45,31,45,30,121,31,51,31,203,31,56,31,145,31,145,30,245,31,181,31,14,31,159,31,75,31,81,31,81,30,194,31,93,31,247,31,227,31,252,31,11,31,252,31,252,30,162,31,59,31,224,31,215,31,17,31,30,31,202,31,233,31,66,31,167,31,167,30,127,31,127,30,127,29,127,28,142,31,55,31,234,31,50,31,243,31,145,31,137,31,137,30,168,31,215,31,209,31,234,31,47,31,37,31,106,31,148,31,216,31,183,31,73,31,76,31,12,31,73,31,223,31,97,31,168,31,168,30,183,31,93,31,93,30,122,31,201,31,244,31,244,30,94,31,58,31,58,30,173,31,152,31,183,31,213,31,213,30,213,29,157,31,199,31,131,31,131,30,131,29,117,31,117,30,111,31,127,31,195,31,184,31,184,30,151,31,53,31,163,31,86,31,125,31,125,30,84,31,81,31,126,31,199,31,191,31,191,30,227,31,208,31,208,30,17,31,20,31,190,31,190,31,187,31,132,31,223,31,223,30,227,31,227,30,227,29,228,31,228,30,22,31,237,31,157,31,70,31,88,31,18,31,55,31,55,30,176,31,184,31,184,30,19,31,63,31,200,31,192,31,48,31,17,31,18,31,143,31,143,30,11,31,237,31,220,31,213,31,213,30,81,31,81,30,241,31,207,31,98,31,226,31,211,31,211,30,230,31,7,31,44,31,219,31,109,31,47,31,123,31,125,31,129,31,205,31,139,31,139,30,95,31,65,31,65,30,174,31,175,31,136,31,194,31,8,31,194,31,194,30,68,31,68,31,170,31,62,31,139,31,173,31,135,31,34,31,15,31,174,31,113,31,3,31,3,30,3,29,140,31,144,31,178,31,112,31,109,31,109,30,22,31,193,31,144,31,134,31,231,31,120,31,111,31,81,31,132,31,25,31,240,31,33,31,42,31,60,31,12,31,74,31,199,31,94,31,94,30,98,31,98,30,158,31,77,31,157,31,88,31,58,31,39,31,5,31,6,31,116,31,201,31,201,30,83,31,27,31,186,31,171,31,171,30,171,29,214,31,116,31,148,31,241,31,152,31,108,31,108,30,109,31,31,31,248,31,205,31,138,31,197,31,101,31,213,31,222,31,79,31,1,31,195,31,136,31,154,31,174,31,57,31,57,30,124,31,147,31,147,30,117,31,20,31,20,30,228,31,60,31,60,30,68,31,29,31,146,31,146,30,110,31,234,31,236,31,49,31,255,31,255,30,255,29,201,31,253,31,115,31,70,31,101,31,101,30,134,31,155,31,96,31,231,31,109,31,109,30,76,31,52,31,126,31,224,31,48,31,56,31,56,30,212,31,75,31,18,31,224,31,224,30,23,31,135,31,83,31,167,31,201,31,49,31,186,31,186,30,99,31,99,30,96,31,22,31,169,31,202,31,177,31,253,31,112,31,50,31,50,30,50,31,28,31,192,31,25,31,91,31,91,30,171,31,180,31,70,31,31,31,31,30,63,31,167,31,99,31,105,31,160,31,113,31,217,31,2,31,166,31,166,30,130,31,101,31,101,30,101,29,80,31,103,31,44,31,212,31,83,31,83,30,149,31,149,30,215,31,216,31,225,31,17,31,157,31,3,31,193,31,156,31,45,31,31,31,147,31,12,31,12,30,156,31,30,31,47,31,48,31,176,31,47,31,7,31,7,30,216,31,92,31,67,31,190,31,37,31,145,31,145,30,38,31,242,31,63,31,63,30,188,31,88,31,203,31,159,31,109,31,3,31,101,31,237,31,80,31,120,31,54,31,54,30,63,31,137,31,144,31,111,31,138,31,138,30,199,31,199,30,173,31,66,31,36,31,124,31,191,31,191,30,191,29,11,31,184,31,21,31,242,31,105,31,203,31,89,31,55,31,238,31,133,31,228,31,88,31,112,31,248,31,81,31,241,31,241,30,142,31,132,31,132,30,121,31,2,31,181,31,181,30,19,31,4,31,4,30,96,31,123,31,205,31,217,31,12,31,12,30,219,31,191,31,6,31,85,31,9,31,216,31,216,30,216,29,112,31,132,31,74,31,36,31,118,31,168,31,68,31,125,31,177,31,89,31,158,31,239,31,160,31,160,30,11,31,11,30,29,31,86,31,240,31,229,31,229,30,229,29,229,28,229,27,201,31,11,31,11,30,115,31,115,30,115,29,115,28,91,31,26,31,12,31,215,31,215,30,7,31,7,30,25,31,173,31,173,30,57,31,42,31,42,30,38,31,207,31,229,31,219,31,204,31,105,31,155,31,251,31,166,31,39,31,39,30,189,31,13,31,9,31,31,31,101,31,82,31,106,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
