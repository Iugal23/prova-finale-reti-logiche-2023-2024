-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 623;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (102,0,165,0,196,0,111,0,44,0,167,0,163,0,128,0,191,0,198,0,109,0,83,0,141,0,140,0,0,0,0,0,0,0,204,0,81,0,184,0,94,0,83,0,0,0,191,0,86,0,241,0,78,0,2,0,237,0,201,0,127,0,252,0,120,0,195,0,54,0,226,0,138,0,0,0,147,0,0,0,206,0,33,0,68,0,157,0,80,0,110,0,0,0,53,0,0,0,148,0,0,0,186,0,187,0,5,0,146,0,65,0,245,0,218,0,186,0,68,0,153,0,38,0,246,0,0,0,57,0,119,0,73,0,40,0,65,0,0,0,45,0,50,0,0,0,32,0,50,0,0,0,27,0,236,0,131,0,103,0,21,0,1,0,0,0,50,0,150,0,76,0,176,0,0,0,187,0,200,0,2,0,197,0,196,0,19,0,179,0,64,0,0,0,207,0,135,0,1,0,154,0,166,0,132,0,5,0,99,0,188,0,170,0,98,0,101,0,181,0,57,0,2,0,107,0,185,0,0,0,196,0,86,0,230,0,61,0,147,0,214,0,228,0,136,0,76,0,195,0,135,0,132,0,0,0,67,0,204,0,0,0,121,0,0,0,252,0,111,0,209,0,204,0,0,0,0,0,120,0,60,0,54,0,255,0,77,0,0,0,168,0,42,0,21,0,112,0,0,0,228,0,232,0,77,0,27,0,72,0,0,0,69,0,32,0,217,0,0,0,0,0,5,0,137,0,117,0,0,0,29,0,216,0,24,0,33,0,113,0,97,0,215,0,186,0,113,0,239,0,30,0,233,0,120,0,0,0,165,0,89,0,223,0,168,0,101,0,23,0,195,0,180,0,5,0,157,0,5,0,36,0,229,0,40,0,125,0,118,0,0,0,0,0,216,0,0,0,222,0,123,0,139,0,162,0,0,0,45,0,0,0,144,0,138,0,165,0,120,0,20,0,195,0,86,0,78,0,72,0,77,0,59,0,243,0,89,0,247,0,36,0,0,0,41,0,141,0,57,0,152,0,139,0,0,0,107,0,0,0,87,0,69,0,27,0,101,0,0,0,0,0,255,0,151,0,255,0,0,0,231,0,0,0,93,0,154,0,118,0,0,0,106,0,0,0,168,0,150,0,114,0,207,0,0,0,22,0,0,0,0,0,107,0,233,0,170,0,0,0,23,0,116,0,219,0,201,0,33,0,22,0,0,0,126,0,25,0,103,0,54,0,0,0,60,0,77,0,0,0,13,0,128,0,112,0,152,0,136,0,139,0,201,0,219,0,0,0,157,0,75,0,133,0,54,0,0,0,179,0,207,0,59,0,12,0,0,0,93,0,0,0,0,0,0,0,28,0,26,0,0,0,104,0,10,0,149,0,8,0,50,0,170,0,36,0,183,0,29,0,0,0,162,0,19,0,96,0,33,0,170,0,0,0,195,0,249,0,0,0,19,0,0,0,152,0,0,0,0,0,63,0,195,0,0,0,87,0,194,0,170,0,240,0,0,0,147,0,0,0,0,0,193,0,83,0,33,0,91,0,0,0,206,0,26,0,4,0,117,0,4,0,153,0,0,0,26,0,48,0,7,0,0,0,162,0,0,0,213,0,206,0,238,0,27,0,150,0,17,0,212,0,238,0,143,0,0,0,215,0,185,0,148,0,239,0,19,0,92,0,57,0,148,0,125,0,33,0,168,0,1,0,156,0,255,0,177,0,43,0,190,0,0,0,96,0,103,0,102,0,182,0,88,0,151,0,169,0,45,0,108,0,9,0,0,0,183,0,70,0,107,0,12,0,241,0,81,0,0,0,20,0,253,0,196,0,143,0,0,0,117,0,56,0,0,0,191,0,123,0,130,0,248,0,59,0,253,0,0,0,195,0,19,0,216,0,0,0,95,0,0,0,0,0,235,0,3,0,62,0,130,0,0,0,85,0,230,0,32,0,220,0,50,0,156,0,190,0,172,0,47,0,0,0,0,0,151,0,0,0,148,0,199,0,67,0,131,0,114,0,0,0,57,0,243,0,0,0,0,0,50,0,0,0,99,0,159,0,233,0,42,0,0,0,109,0,0,0,218,0,149,0,150,0,191,0,66,0,91,0,139,0,78,0,26,0,12,0,48,0,79,0,0,0,0,0,185,0,0,0,0,0,0,0,155,0,179,0,0,0,16,0,0,0,236,0,221,0,27,0,44,0,0,0,252,0,56,0,67,0,41,0,226,0,217,0,30,0,245,0,105,0,152,0,0,0,0,0,197,0,192,0,165,0,143,0,82,0,0,0,94,0,144,0,207,0,0,0,131,0,164,0,0,0,0,0,234,0,146,0,168,0,0,0,222,0,235,0,185,0,237,0,0,0,229,0,104,0,187,0,62,0,155,0,0,0,47,0,60,0,43,0,0,0,83,0,89,0,2,0,95,0,1,0,18,0,224,0,108,0,0,0,190,0,160,0,220,0,244,0,0,0,33,0,0,0,225,0,221,0,216,0,86,0,211,0,0,0,54,0,0,0,157,0,125,0,17,0,22,0,0,0,72,0,227,0,211,0,239,0,185,0,0,0,170,0,0,0,0,0,174,0,120,0,48,0,119,0,132,0,113,0,163,0,85,0,0,0,0,0,143,0,246,0,82,0,29,0,58,0,0,0,171,0,67,0,148,0,187,0,124,0,0,0,157,0,0,0,0,0,56,0,215,0,28,0,229,0,0,0,0,0,142,0,0,0,252,0,83,0,133,0,21,0,170,0,116,0,64,0,32,0,68,0,161,0,142,0,84,0,254,0,213,0,9,0,132,0,0,0,70,0,37,0,9,0);
signal scenario_full  : scenario_type := (102,31,165,31,196,31,111,31,44,31,167,31,163,31,128,31,191,31,198,31,109,31,83,31,141,31,140,31,140,30,140,29,140,28,204,31,81,31,184,31,94,31,83,31,83,30,191,31,86,31,241,31,78,31,2,31,237,31,201,31,127,31,252,31,120,31,195,31,54,31,226,31,138,31,138,30,147,31,147,30,206,31,33,31,68,31,157,31,80,31,110,31,110,30,53,31,53,30,148,31,148,30,186,31,187,31,5,31,146,31,65,31,245,31,218,31,186,31,68,31,153,31,38,31,246,31,246,30,57,31,119,31,73,31,40,31,65,31,65,30,45,31,50,31,50,30,32,31,50,31,50,30,27,31,236,31,131,31,103,31,21,31,1,31,1,30,50,31,150,31,76,31,176,31,176,30,187,31,200,31,2,31,197,31,196,31,19,31,179,31,64,31,64,30,207,31,135,31,1,31,154,31,166,31,132,31,5,31,99,31,188,31,170,31,98,31,101,31,181,31,57,31,2,31,107,31,185,31,185,30,196,31,86,31,230,31,61,31,147,31,214,31,228,31,136,31,76,31,195,31,135,31,132,31,132,30,67,31,204,31,204,30,121,31,121,30,252,31,111,31,209,31,204,31,204,30,204,29,120,31,60,31,54,31,255,31,77,31,77,30,168,31,42,31,21,31,112,31,112,30,228,31,232,31,77,31,27,31,72,31,72,30,69,31,32,31,217,31,217,30,217,29,5,31,137,31,117,31,117,30,29,31,216,31,24,31,33,31,113,31,97,31,215,31,186,31,113,31,239,31,30,31,233,31,120,31,120,30,165,31,89,31,223,31,168,31,101,31,23,31,195,31,180,31,5,31,157,31,5,31,36,31,229,31,40,31,125,31,118,31,118,30,118,29,216,31,216,30,222,31,123,31,139,31,162,31,162,30,45,31,45,30,144,31,138,31,165,31,120,31,20,31,195,31,86,31,78,31,72,31,77,31,59,31,243,31,89,31,247,31,36,31,36,30,41,31,141,31,57,31,152,31,139,31,139,30,107,31,107,30,87,31,69,31,27,31,101,31,101,30,101,29,255,31,151,31,255,31,255,30,231,31,231,30,93,31,154,31,118,31,118,30,106,31,106,30,168,31,150,31,114,31,207,31,207,30,22,31,22,30,22,29,107,31,233,31,170,31,170,30,23,31,116,31,219,31,201,31,33,31,22,31,22,30,126,31,25,31,103,31,54,31,54,30,60,31,77,31,77,30,13,31,128,31,112,31,152,31,136,31,139,31,201,31,219,31,219,30,157,31,75,31,133,31,54,31,54,30,179,31,207,31,59,31,12,31,12,30,93,31,93,30,93,29,93,28,28,31,26,31,26,30,104,31,10,31,149,31,8,31,50,31,170,31,36,31,183,31,29,31,29,30,162,31,19,31,96,31,33,31,170,31,170,30,195,31,249,31,249,30,19,31,19,30,152,31,152,30,152,29,63,31,195,31,195,30,87,31,194,31,170,31,240,31,240,30,147,31,147,30,147,29,193,31,83,31,33,31,91,31,91,30,206,31,26,31,4,31,117,31,4,31,153,31,153,30,26,31,48,31,7,31,7,30,162,31,162,30,213,31,206,31,238,31,27,31,150,31,17,31,212,31,238,31,143,31,143,30,215,31,185,31,148,31,239,31,19,31,92,31,57,31,148,31,125,31,33,31,168,31,1,31,156,31,255,31,177,31,43,31,190,31,190,30,96,31,103,31,102,31,182,31,88,31,151,31,169,31,45,31,108,31,9,31,9,30,183,31,70,31,107,31,12,31,241,31,81,31,81,30,20,31,253,31,196,31,143,31,143,30,117,31,56,31,56,30,191,31,123,31,130,31,248,31,59,31,253,31,253,30,195,31,19,31,216,31,216,30,95,31,95,30,95,29,235,31,3,31,62,31,130,31,130,30,85,31,230,31,32,31,220,31,50,31,156,31,190,31,172,31,47,31,47,30,47,29,151,31,151,30,148,31,199,31,67,31,131,31,114,31,114,30,57,31,243,31,243,30,243,29,50,31,50,30,99,31,159,31,233,31,42,31,42,30,109,31,109,30,218,31,149,31,150,31,191,31,66,31,91,31,139,31,78,31,26,31,12,31,48,31,79,31,79,30,79,29,185,31,185,30,185,29,185,28,155,31,179,31,179,30,16,31,16,30,236,31,221,31,27,31,44,31,44,30,252,31,56,31,67,31,41,31,226,31,217,31,30,31,245,31,105,31,152,31,152,30,152,29,197,31,192,31,165,31,143,31,82,31,82,30,94,31,144,31,207,31,207,30,131,31,164,31,164,30,164,29,234,31,146,31,168,31,168,30,222,31,235,31,185,31,237,31,237,30,229,31,104,31,187,31,62,31,155,31,155,30,47,31,60,31,43,31,43,30,83,31,89,31,2,31,95,31,1,31,18,31,224,31,108,31,108,30,190,31,160,31,220,31,244,31,244,30,33,31,33,30,225,31,221,31,216,31,86,31,211,31,211,30,54,31,54,30,157,31,125,31,17,31,22,31,22,30,72,31,227,31,211,31,239,31,185,31,185,30,170,31,170,30,170,29,174,31,120,31,48,31,119,31,132,31,113,31,163,31,85,31,85,30,85,29,143,31,246,31,82,31,29,31,58,31,58,30,171,31,67,31,148,31,187,31,124,31,124,30,157,31,157,30,157,29,56,31,215,31,28,31,229,31,229,30,229,29,142,31,142,30,252,31,83,31,133,31,21,31,170,31,116,31,64,31,32,31,68,31,161,31,142,31,84,31,254,31,213,31,9,31,132,31,132,30,70,31,37,31,9,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
