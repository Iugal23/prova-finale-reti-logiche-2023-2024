-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_51 is
end project_tb_51;

architecture project_tb_arch_51 of project_tb_51 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 995;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (173,0,20,0,65,0,0,0,33,0,103,0,47,0,0,0,0,0,165,0,11,0,33,0,0,0,69,0,0,0,217,0,3,0,0,0,153,0,97,0,221,0,0,0,65,0,0,0,21,0,38,0,64,0,131,0,102,0,0,0,244,0,78,0,178,0,107,0,209,0,9,0,0,0,0,0,169,0,176,0,0,0,15,0,253,0,78,0,201,0,78,0,133,0,0,0,59,0,0,0,118,0,55,0,51,0,16,0,129,0,41,0,18,0,0,0,66,0,15,0,60,0,144,0,165,0,92,0,26,0,0,0,142,0,98,0,163,0,4,0,52,0,26,0,0,0,118,0,231,0,209,0,75,0,198,0,155,0,4,0,14,0,119,0,127,0,252,0,167,0,137,0,115,0,0,0,0,0,165,0,178,0,41,0,42,0,49,0,45,0,0,0,128,0,213,0,39,0,199,0,40,0,65,0,0,0,235,0,137,0,117,0,247,0,197,0,79,0,237,0,236,0,203,0,201,0,92,0,122,0,88,0,242,0,91,0,162,0,23,0,138,0,93,0,255,0,141,0,196,0,0,0,127,0,0,0,166,0,221,0,0,0,218,0,0,0,0,0,0,0,42,0,195,0,80,0,0,0,100,0,0,0,126,0,7,0,0,0,74,0,36,0,95,0,0,0,210,0,11,0,12,0,166,0,192,0,0,0,238,0,30,0,209,0,219,0,235,0,7,0,20,0,159,0,241,0,172,0,17,0,189,0,120,0,46,0,0,0,0,0,0,0,0,0,13,0,16,0,144,0,0,0,7,0,181,0,241,0,53,0,121,0,17,0,90,0,80,0,0,0,61,0,180,0,82,0,78,0,108,0,99,0,0,0,0,0,157,0,26,0,94,0,0,0,0,0,71,0,59,0,46,0,112,0,56,0,70,0,181,0,243,0,17,0,147,0,252,0,241,0,0,0,132,0,161,0,226,0,202,0,199,0,40,0,158,0,65,0,163,0,0,0,0,0,28,0,116,0,0,0,252,0,76,0,210,0,68,0,200,0,0,0,130,0,199,0,252,0,46,0,189,0,137,0,124,0,163,0,49,0,143,0,29,0,34,0,101,0,149,0,129,0,40,0,73,0,110,0,93,0,220,0,0,0,233,0,28,0,50,0,67,0,183,0,0,0,13,0,0,0,74,0,253,0,8,0,213,0,142,0,149,0,242,0,194,0,0,0,184,0,0,0,0,0,0,0,0,0,190,0,26,0,32,0,0,0,74,0,115,0,172,0,234,0,167,0,63,0,0,0,66,0,177,0,51,0,170,0,249,0,77,0,194,0,125,0,199,0,226,0,73,0,191,0,12,0,0,0,10,0,171,0,88,0,30,0,37,0,179,0,221,0,82,0,12,0,29,0,171,0,73,0,0,0,190,0,225,0,74,0,251,0,138,0,0,0,64,0,0,0,132,0,0,0,240,0,23,0,74,0,52,0,120,0,217,0,64,0,61,0,155,0,242,0,243,0,0,0,16,0,134,0,108,0,132,0,87,0,95,0,92,0,19,0,217,0,109,0,0,0,181,0,74,0,0,0,39,0,2,0,53,0,9,0,16,0,254,0,79,0,133,0,102,0,244,0,46,0,189,0,32,0,147,0,161,0,86,0,16,0,78,0,69,0,46,0,0,0,32,0,79,0,191,0,0,0,36,0,133,0,0,0,140,0,245,0,0,0,0,0,0,0,111,0,154,0,10,0,129,0,0,0,241,0,164,0,22,0,70,0,95,0,152,0,0,0,0,0,153,0,175,0,142,0,0,0,231,0,239,0,0,0,0,0,0,0,78,0,0,0,48,0,159,0,71,0,99,0,95,0,0,0,0,0,29,0,118,0,84,0,210,0,160,0,50,0,62,0,45,0,132,0,0,0,236,0,135,0,182,0,105,0,0,0,113,0,81,0,165,0,0,0,213,0,209,0,234,0,231,0,244,0,46,0,192,0,13,0,204,0,29,0,203,0,160,0,0,0,0,0,0,0,57,0,192,0,221,0,133,0,201,0,0,0,26,0,140,0,0,0,0,0,128,0,59,0,118,0,110,0,0,0,16,0,158,0,0,0,0,0,2,0,212,0,151,0,178,0,0,0,87,0,158,0,32,0,146,0,191,0,166,0,76,0,236,0,21,0,1,0,53,0,2,0,184,0,107,0,206,0,235,0,8,0,68,0,146,0,4,0,0,0,0,0,40,0,51,0,253,0,80,0,246,0,212,0,149,0,46,0,0,0,109,0,225,0,0,0,0,0,3,0,73,0,122,0,214,0,32,0,168,0,0,0,26,0,59,0,0,0,174,0,1,0,0,0,207,0,174,0,35,0,206,0,175,0,38,0,13,0,13,0,11,0,202,0,187,0,168,0,218,0,108,0,165,0,34,0,208,0,0,0,100,0,229,0,87,0,91,0,106,0,233,0,193,0,0,0,105,0,145,0,95,0,150,0,234,0,137,0,0,0,0,0,71,0,164,0,186,0,193,0,245,0,11,0,138,0,44,0,246,0,186,0,111,0,48,0,8,0,0,0,177,0,244,0,82,0,212,0,94,0,22,0,127,0,110,0,133,0,167,0,144,0,9,0,153,0,0,0,101,0,2,0,26,0,58,0,82,0,123,0,236,0,171,0,142,0,51,0,46,0,74,0,163,0,71,0,85,0,64,0,102,0,96,0,134,0,80,0,182,0,123,0,87,0,241,0,189,0,170,0,84,0,226,0,154,0,182,0,92,0,238,0,0,0,174,0,78,0,208,0,0,0,19,0,0,0,0,0,55,0,147,0,0,0,166,0,97,0,112,0,97,0,148,0,184,0,52,0,0,0,219,0,0,0,159,0,128,0,122,0,29,0,95,0,5,0,228,0,16,0,204,0,29,0,203,0,99,0,255,0,72,0,226,0,198,0,189,0,42,0,198,0,72,0,150,0,73,0,208,0,216,0,27,0,167,0,120,0,228,0,241,0,233,0,62,0,162,0,0,0,99,0,105,0,0,0,219,0,95,0,65,0,0,0,104,0,213,0,95,0,0,0,111,0,0,0,30,0,149,0,0,0,81,0,26,0,0,0,0,0,93,0,0,0,0,0,78,0,215,0,177,0,0,0,249,0,225,0,254,0,0,0,167,0,0,0,107,0,130,0,182,0,60,0,94,0,0,0,62,0,73,0,0,0,167,0,144,0,208,0,143,0,81,0,19,0,74,0,252,0,0,0,124,0,175,0,175,0,190,0,145,0,226,0,110,0,0,0,0,0,207,0,64,0,102,0,133,0,172,0,0,0,212,0,0,0,250,0,18,0,0,0,0,0,0,0,126,0,16,0,153,0,245,0,150,0,145,0,194,0,17,0,243,0,0,0,106,0,142,0,0,0,120,0,236,0,58,0,105,0,210,0,185,0,0,0,146,0,0,0,247,0,156,0,214,0,0,0,0,0,237,0,93,0,0,0,211,0,174,0,97,0,0,0,0,0,97,0,216,0,46,0,28,0,252,0,0,0,0,0,0,0,0,0,46,0,0,0,143,0,124,0,0,0,61,0,0,0,185,0,64,0,195,0,181,0,251,0,75,0,0,0,0,0,0,0,119,0,221,0,91,0,234,0,22,0,198,0,213,0,20,0,37,0,0,0,0,0,64,0,178,0,107,0,144,0,116,0,20,0,104,0,53,0,152,0,0,0,54,0,177,0,219,0,185,0,24,0,166,0,43,0,154,0,127,0,0,0,0,0,219,0,255,0,0,0,246,0,128,0,237,0,91,0,118,0,0,0,97,0,178,0,14,0,66,0,241,0,39,0,21,0,7,0,26,0,202,0,46,0,21,0,53,0,0,0,228,0,106,0,65,0,57,0,133,0,71,0,112,0,73,0,219,0,143,0,85,0,111,0,202,0,196,0,246,0,126,0,17,0,111,0,208,0,25,0,199,0,187,0,62,0,148,0,198,0,161,0,234,0,246,0,32,0,0,0,224,0,0,0,197,0,0,0,0,0,0,0,239,0,0,0,7,0,5,0,183,0,0,0,240,0,34,0,189,0,242,0,104,0,126,0,221,0,171,0,203,0,146,0,23,0,10,0,180,0,0,0,245,0,0,0,65,0,0,0,7,0,0,0,0,0,51,0,0,0,0,0,129,0,236,0,205,0,0,0,202,0,0,0,24,0,0,0,107,0,26,0,55,0,129,0,0,0,14,0,128,0,71,0,0,0,71,0,29,0,63,0,123,0,242,0,121,0,45,0,29,0,188,0,59,0,138,0,0,0,87,0,15,0,4,0,252,0,82,0,29,0,249,0,228,0,0,0,210,0,49,0,241,0,20,0,66,0,219,0,0,0,67,0,245,0,0,0,99,0,226,0,0,0,171,0,242,0,40,0,92,0,3,0,207,0,136,0,148,0,68,0,164,0,105,0,16,0,78,0,85,0,161,0,0,0,186,0,195,0,25,0,32,0,135,0,248,0,0,0,103,0);
signal scenario_full  : scenario_type := (173,31,20,31,65,31,65,30,33,31,103,31,47,31,47,30,47,29,165,31,11,31,33,31,33,30,69,31,69,30,217,31,3,31,3,30,153,31,97,31,221,31,221,30,65,31,65,30,21,31,38,31,64,31,131,31,102,31,102,30,244,31,78,31,178,31,107,31,209,31,9,31,9,30,9,29,169,31,176,31,176,30,15,31,253,31,78,31,201,31,78,31,133,31,133,30,59,31,59,30,118,31,55,31,51,31,16,31,129,31,41,31,18,31,18,30,66,31,15,31,60,31,144,31,165,31,92,31,26,31,26,30,142,31,98,31,163,31,4,31,52,31,26,31,26,30,118,31,231,31,209,31,75,31,198,31,155,31,4,31,14,31,119,31,127,31,252,31,167,31,137,31,115,31,115,30,115,29,165,31,178,31,41,31,42,31,49,31,45,31,45,30,128,31,213,31,39,31,199,31,40,31,65,31,65,30,235,31,137,31,117,31,247,31,197,31,79,31,237,31,236,31,203,31,201,31,92,31,122,31,88,31,242,31,91,31,162,31,23,31,138,31,93,31,255,31,141,31,196,31,196,30,127,31,127,30,166,31,221,31,221,30,218,31,218,30,218,29,218,28,42,31,195,31,80,31,80,30,100,31,100,30,126,31,7,31,7,30,74,31,36,31,95,31,95,30,210,31,11,31,12,31,166,31,192,31,192,30,238,31,30,31,209,31,219,31,235,31,7,31,20,31,159,31,241,31,172,31,17,31,189,31,120,31,46,31,46,30,46,29,46,28,46,27,13,31,16,31,144,31,144,30,7,31,181,31,241,31,53,31,121,31,17,31,90,31,80,31,80,30,61,31,180,31,82,31,78,31,108,31,99,31,99,30,99,29,157,31,26,31,94,31,94,30,94,29,71,31,59,31,46,31,112,31,56,31,70,31,181,31,243,31,17,31,147,31,252,31,241,31,241,30,132,31,161,31,226,31,202,31,199,31,40,31,158,31,65,31,163,31,163,30,163,29,28,31,116,31,116,30,252,31,76,31,210,31,68,31,200,31,200,30,130,31,199,31,252,31,46,31,189,31,137,31,124,31,163,31,49,31,143,31,29,31,34,31,101,31,149,31,129,31,40,31,73,31,110,31,93,31,220,31,220,30,233,31,28,31,50,31,67,31,183,31,183,30,13,31,13,30,74,31,253,31,8,31,213,31,142,31,149,31,242,31,194,31,194,30,184,31,184,30,184,29,184,28,184,27,190,31,26,31,32,31,32,30,74,31,115,31,172,31,234,31,167,31,63,31,63,30,66,31,177,31,51,31,170,31,249,31,77,31,194,31,125,31,199,31,226,31,73,31,191,31,12,31,12,30,10,31,171,31,88,31,30,31,37,31,179,31,221,31,82,31,12,31,29,31,171,31,73,31,73,30,190,31,225,31,74,31,251,31,138,31,138,30,64,31,64,30,132,31,132,30,240,31,23,31,74,31,52,31,120,31,217,31,64,31,61,31,155,31,242,31,243,31,243,30,16,31,134,31,108,31,132,31,87,31,95,31,92,31,19,31,217,31,109,31,109,30,181,31,74,31,74,30,39,31,2,31,53,31,9,31,16,31,254,31,79,31,133,31,102,31,244,31,46,31,189,31,32,31,147,31,161,31,86,31,16,31,78,31,69,31,46,31,46,30,32,31,79,31,191,31,191,30,36,31,133,31,133,30,140,31,245,31,245,30,245,29,245,28,111,31,154,31,10,31,129,31,129,30,241,31,164,31,22,31,70,31,95,31,152,31,152,30,152,29,153,31,175,31,142,31,142,30,231,31,239,31,239,30,239,29,239,28,78,31,78,30,48,31,159,31,71,31,99,31,95,31,95,30,95,29,29,31,118,31,84,31,210,31,160,31,50,31,62,31,45,31,132,31,132,30,236,31,135,31,182,31,105,31,105,30,113,31,81,31,165,31,165,30,213,31,209,31,234,31,231,31,244,31,46,31,192,31,13,31,204,31,29,31,203,31,160,31,160,30,160,29,160,28,57,31,192,31,221,31,133,31,201,31,201,30,26,31,140,31,140,30,140,29,128,31,59,31,118,31,110,31,110,30,16,31,158,31,158,30,158,29,2,31,212,31,151,31,178,31,178,30,87,31,158,31,32,31,146,31,191,31,166,31,76,31,236,31,21,31,1,31,53,31,2,31,184,31,107,31,206,31,235,31,8,31,68,31,146,31,4,31,4,30,4,29,40,31,51,31,253,31,80,31,246,31,212,31,149,31,46,31,46,30,109,31,225,31,225,30,225,29,3,31,73,31,122,31,214,31,32,31,168,31,168,30,26,31,59,31,59,30,174,31,1,31,1,30,207,31,174,31,35,31,206,31,175,31,38,31,13,31,13,31,11,31,202,31,187,31,168,31,218,31,108,31,165,31,34,31,208,31,208,30,100,31,229,31,87,31,91,31,106,31,233,31,193,31,193,30,105,31,145,31,95,31,150,31,234,31,137,31,137,30,137,29,71,31,164,31,186,31,193,31,245,31,11,31,138,31,44,31,246,31,186,31,111,31,48,31,8,31,8,30,177,31,244,31,82,31,212,31,94,31,22,31,127,31,110,31,133,31,167,31,144,31,9,31,153,31,153,30,101,31,2,31,26,31,58,31,82,31,123,31,236,31,171,31,142,31,51,31,46,31,74,31,163,31,71,31,85,31,64,31,102,31,96,31,134,31,80,31,182,31,123,31,87,31,241,31,189,31,170,31,84,31,226,31,154,31,182,31,92,31,238,31,238,30,174,31,78,31,208,31,208,30,19,31,19,30,19,29,55,31,147,31,147,30,166,31,97,31,112,31,97,31,148,31,184,31,52,31,52,30,219,31,219,30,159,31,128,31,122,31,29,31,95,31,5,31,228,31,16,31,204,31,29,31,203,31,99,31,255,31,72,31,226,31,198,31,189,31,42,31,198,31,72,31,150,31,73,31,208,31,216,31,27,31,167,31,120,31,228,31,241,31,233,31,62,31,162,31,162,30,99,31,105,31,105,30,219,31,95,31,65,31,65,30,104,31,213,31,95,31,95,30,111,31,111,30,30,31,149,31,149,30,81,31,26,31,26,30,26,29,93,31,93,30,93,29,78,31,215,31,177,31,177,30,249,31,225,31,254,31,254,30,167,31,167,30,107,31,130,31,182,31,60,31,94,31,94,30,62,31,73,31,73,30,167,31,144,31,208,31,143,31,81,31,19,31,74,31,252,31,252,30,124,31,175,31,175,31,190,31,145,31,226,31,110,31,110,30,110,29,207,31,64,31,102,31,133,31,172,31,172,30,212,31,212,30,250,31,18,31,18,30,18,29,18,28,126,31,16,31,153,31,245,31,150,31,145,31,194,31,17,31,243,31,243,30,106,31,142,31,142,30,120,31,236,31,58,31,105,31,210,31,185,31,185,30,146,31,146,30,247,31,156,31,214,31,214,30,214,29,237,31,93,31,93,30,211,31,174,31,97,31,97,30,97,29,97,31,216,31,46,31,28,31,252,31,252,30,252,29,252,28,252,27,46,31,46,30,143,31,124,31,124,30,61,31,61,30,185,31,64,31,195,31,181,31,251,31,75,31,75,30,75,29,75,28,119,31,221,31,91,31,234,31,22,31,198,31,213,31,20,31,37,31,37,30,37,29,64,31,178,31,107,31,144,31,116,31,20,31,104,31,53,31,152,31,152,30,54,31,177,31,219,31,185,31,24,31,166,31,43,31,154,31,127,31,127,30,127,29,219,31,255,31,255,30,246,31,128,31,237,31,91,31,118,31,118,30,97,31,178,31,14,31,66,31,241,31,39,31,21,31,7,31,26,31,202,31,46,31,21,31,53,31,53,30,228,31,106,31,65,31,57,31,133,31,71,31,112,31,73,31,219,31,143,31,85,31,111,31,202,31,196,31,246,31,126,31,17,31,111,31,208,31,25,31,199,31,187,31,62,31,148,31,198,31,161,31,234,31,246,31,32,31,32,30,224,31,224,30,197,31,197,30,197,29,197,28,239,31,239,30,7,31,5,31,183,31,183,30,240,31,34,31,189,31,242,31,104,31,126,31,221,31,171,31,203,31,146,31,23,31,10,31,180,31,180,30,245,31,245,30,65,31,65,30,7,31,7,30,7,29,51,31,51,30,51,29,129,31,236,31,205,31,205,30,202,31,202,30,24,31,24,30,107,31,26,31,55,31,129,31,129,30,14,31,128,31,71,31,71,30,71,31,29,31,63,31,123,31,242,31,121,31,45,31,29,31,188,31,59,31,138,31,138,30,87,31,15,31,4,31,252,31,82,31,29,31,249,31,228,31,228,30,210,31,49,31,241,31,20,31,66,31,219,31,219,30,67,31,245,31,245,30,99,31,226,31,226,30,171,31,242,31,40,31,92,31,3,31,207,31,136,31,148,31,68,31,164,31,105,31,16,31,78,31,85,31,161,31,161,30,186,31,195,31,25,31,32,31,135,31,248,31,248,30,103,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
