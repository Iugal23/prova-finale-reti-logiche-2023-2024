-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_335 is
end project_tb_335;

architecture project_tb_arch_335 of project_tb_335 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 978;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (136,0,180,0,0,0,96,0,10,0,66,0,0,0,0,0,0,0,81,0,39,0,171,0,5,0,207,0,0,0,61,0,125,0,225,0,33,0,207,0,27,0,2,0,210,0,19,0,141,0,0,0,229,0,0,0,12,0,138,0,49,0,142,0,12,0,40,0,35,0,0,0,210,0,211,0,0,0,148,0,158,0,121,0,59,0,239,0,142,0,179,0,198,0,121,0,0,0,0,0,116,0,0,0,0,0,0,0,64,0,63,0,244,0,65,0,43,0,0,0,53,0,208,0,0,0,33,0,0,0,0,0,26,0,128,0,108,0,135,0,40,0,40,0,144,0,63,0,175,0,88,0,136,0,0,0,0,0,171,0,146,0,0,0,249,0,253,0,173,0,139,0,233,0,107,0,122,0,36,0,130,0,210,0,121,0,93,0,128,0,11,0,0,0,22,0,41,0,233,0,60,0,218,0,199,0,0,0,210,0,140,0,135,0,0,0,0,0,0,0,38,0,65,0,0,0,0,0,188,0,0,0,142,0,236,0,109,0,64,0,176,0,0,0,220,0,0,0,0,0,0,0,211,0,185,0,0,0,245,0,133,0,104,0,225,0,117,0,163,0,228,0,248,0,145,0,105,0,179,0,40,0,0,0,207,0,49,0,175,0,157,0,0,0,10,0,156,0,172,0,182,0,0,0,106,0,224,0,49,0,48,0,0,0,207,0,234,0,211,0,222,0,220,0,235,0,57,0,1,0,146,0,106,0,2,0,9,0,0,0,164,0,40,0,212,0,70,0,0,0,20,0,208,0,33,0,148,0,252,0,182,0,236,0,42,0,185,0,178,0,207,0,23,0,98,0,98,0,78,0,21,0,0,0,0,0,144,0,131,0,66,0,145,0,191,0,107,0,0,0,0,0,253,0,193,0,80,0,64,0,251,0,16,0,130,0,127,0,110,0,60,0,222,0,2,0,73,0,67,0,2,0,241,0,51,0,183,0,0,0,0,0,0,0,37,0,184,0,134,0,187,0,113,0,67,0,129,0,0,0,240,0,96,0,205,0,229,0,77,0,255,0,51,0,91,0,0,0,0,0,158,0,204,0,160,0,174,0,0,0,214,0,118,0,0,0,200,0,238,0,221,0,0,0,210,0,0,0,135,0,99,0,119,0,101,0,241,0,211,0,5,0,131,0,76,0,125,0,251,0,208,0,136,0,13,0,30,0,64,0,93,0,1,0,63,0,33,0,121,0,50,0,158,0,74,0,161,0,0,0,0,0,110,0,136,0,240,0,0,0,0,0,53,0,111,0,216,0,235,0,0,0,66,0,241,0,164,0,118,0,0,0,134,0,0,0,46,0,42,0,0,0,224,0,0,0,0,0,204,0,180,0,153,0,222,0,149,0,223,0,0,0,62,0,77,0,100,0,0,0,247,0,252,0,0,0,0,0,0,0,82,0,0,0,0,0,228,0,6,0,41,0,84,0,155,0,76,0,21,0,92,0,83,0,103,0,0,0,0,0,0,0,149,0,234,0,130,0,167,0,39,0,127,0,174,0,241,0,31,0,229,0,26,0,197,0,196,0,26,0,0,0,213,0,0,0,23,0,0,0,222,0,247,0,26,0,96,0,192,0,10,0,174,0,67,0,16,0,0,0,3,0,21,0,142,0,0,0,136,0,48,0,0,0,166,0,188,0,73,0,58,0,78,0,243,0,216,0,170,0,174,0,233,0,107,0,170,0,0,0,0,0,111,0,39,0,177,0,254,0,44,0,93,0,0,0,54,0,20,0,113,0,190,0,129,0,31,0,0,0,202,0,233,0,160,0,118,0,2,0,0,0,32,0,247,0,59,0,161,0,200,0,169,0,209,0,232,0,187,0,155,0,36,0,0,0,27,0,137,0,208,0,255,0,13,0,95,0,6,0,143,0,239,0,219,0,202,0,63,0,90,0,109,0,0,0,220,0,101,0,0,0,235,0,0,0,152,0,0,0,141,0,180,0,137,0,141,0,133,0,91,0,169,0,87,0,175,0,0,0,170,0,168,0,0,0,116,0,180,0,135,0,34,0,208,0,42,0,146,0,119,0,56,0,75,0,250,0,0,0,0,0,204,0,8,0,241,0,201,0,201,0,231,0,139,0,249,0,57,0,254,0,0,0,232,0,51,0,144,0,197,0,143,0,0,0,0,0,62,0,0,0,121,0,131,0,0,0,83,0,0,0,70,0,151,0,0,0,152,0,186,0,181,0,245,0,0,0,76,0,195,0,93,0,191,0,162,0,86,0,0,0,0,0,103,0,140,0,183,0,235,0,111,0,18,0,7,0,118,0,251,0,0,0,178,0,0,0,127,0,57,0,88,0,0,0,20,0,86,0,127,0,192,0,131,0,45,0,0,0,62,0,217,0,221,0,0,0,0,0,180,0,214,0,125,0,176,0,56,0,203,0,152,0,183,0,129,0,10,0,234,0,186,0,113,0,0,0,91,0,0,0,0,0,0,0,0,0,79,0,0,0,238,0,0,0,254,0,68,0,242,0,164,0,0,0,187,0,254,0,113,0,0,0,0,0,205,0,0,0,60,0,145,0,110,0,131,0,253,0,105,0,0,0,36,0,78,0,90,0,213,0,111,0,98,0,203,0,12,0,4,0,67,0,173,0,232,0,0,0,0,0,0,0,0,0,36,0,125,0,0,0,0,0,68,0,0,0,157,0,0,0,131,0,246,0,176,0,0,0,0,0,74,0,246,0,220,0,134,0,183,0,112,0,118,0,61,0,138,0,0,0,0,0,15,0,89,0,0,0,223,0,66,0,228,0,86,0,0,0,131,0,227,0,11,0,141,0,253,0,212,0,47,0,247,0,163,0,39,0,229,0,59,0,0,0,254,0,203,0,165,0,0,0,165,0,160,0,119,0,0,0,211,0,252,0,55,0,153,0,91,0,44,0,7,0,20,0,196,0,97,0,0,0,31,0,45,0,0,0,132,0,232,0,68,0,150,0,0,0,28,0,91,0,251,0,0,0,46,0,86,0,94,0,52,0,20,0,0,0,241,0,177,0,0,0,98,0,161,0,113,0,99,0,208,0,156,0,135,0,22,0,73,0,166,0,130,0,0,0,50,0,213,0,201,0,211,0,97,0,0,0,110,0,207,0,111,0,0,0,68,0,4,0,0,0,24,0,130,0,129,0,1,0,17,0,192,0,133,0,116,0,5,0,210,0,102,0,0,0,228,0,35,0,0,0,175,0,61,0,73,0,96,0,147,0,0,0,0,0,52,0,0,0,206,0,97,0,227,0,4,0,91,0,175,0,2,0,117,0,170,0,0,0,153,0,190,0,33,0,72,0,125,0,88,0,182,0,233,0,0,0,251,0,17,0,113,0,246,0,106,0,122,0,174,0,248,0,158,0,88,0,172,0,158,0,172,0,182,0,167,0,160,0,97,0,201,0,194,0,218,0,37,0,185,0,176,0,160,0,0,0,173,0,214,0,132,0,7,0,158,0,8,0,163,0,148,0,96,0,215,0,97,0,0,0,106,0,0,0,0,0,42,0,215,0,104,0,218,0,239,0,91,0,190,0,184,0,90,0,75,0,73,0,79,0,182,0,91,0,24,0,153,0,147,0,253,0,0,0,229,0,0,0,0,0,113,0,151,0,0,0,105,0,135,0,0,0,150,0,151,0,0,0,0,0,241,0,0,0,25,0,230,0,212,0,248,0,233,0,26,0,101,0,141,0,237,0,178,0,198,0,5,0,244,0,120,0,0,0,82,0,0,0,233,0,137,0,175,0,135,0,108,0,59,0,71,0,99,0,0,0,0,0,157,0,71,0,99,0,0,0,204,0,0,0,0,0,98,0,50,0,20,0,171,0,109,0,0,0,204,0,238,0,85,0,130,0,52,0,10,0,0,0,93,0,119,0,6,0,44,0,172,0,71,0,0,0,30,0,132,0,18,0,16,0,44,0,1,0,198,0,0,0,146,0,74,0,0,0,21,0,0,0,167,0,40,0,95,0,0,0,250,0,165,0,147,0,39,0,59,0,203,0,0,0,235,0,229,0,208,0,136,0,169,0,0,0,0,0,93,0,246,0,72,0,185,0,93,0,88,0,222,0,18,0,103,0,22,0,244,0,99,0,2,0,0,0,0,0,162,0,149,0,130,0,111,0,0,0,145,0,142,0,0,0,22,0,106,0,112,0,187,0,51,0,22,0,151,0,88,0,0,0,137,0,231,0,0,0,153,0,186,0,30,0,0,0,0,0,137,0,221,0,0,0,13,0,154,0,138,0,113,0,68,0,224,0,77,0,208,0,58,0,97,0,73,0,0,0,0,0,173,0,250,0,176,0,250,0,159,0,192,0,117,0,144,0,20,0,246,0,149,0,0,0,0,0,201,0,0,0,0,0,5,0);
signal scenario_full  : scenario_type := (136,31,180,31,180,30,96,31,10,31,66,31,66,30,66,29,66,28,81,31,39,31,171,31,5,31,207,31,207,30,61,31,125,31,225,31,33,31,207,31,27,31,2,31,210,31,19,31,141,31,141,30,229,31,229,30,12,31,138,31,49,31,142,31,12,31,40,31,35,31,35,30,210,31,211,31,211,30,148,31,158,31,121,31,59,31,239,31,142,31,179,31,198,31,121,31,121,30,121,29,116,31,116,30,116,29,116,28,64,31,63,31,244,31,65,31,43,31,43,30,53,31,208,31,208,30,33,31,33,30,33,29,26,31,128,31,108,31,135,31,40,31,40,31,144,31,63,31,175,31,88,31,136,31,136,30,136,29,171,31,146,31,146,30,249,31,253,31,173,31,139,31,233,31,107,31,122,31,36,31,130,31,210,31,121,31,93,31,128,31,11,31,11,30,22,31,41,31,233,31,60,31,218,31,199,31,199,30,210,31,140,31,135,31,135,30,135,29,135,28,38,31,65,31,65,30,65,29,188,31,188,30,142,31,236,31,109,31,64,31,176,31,176,30,220,31,220,30,220,29,220,28,211,31,185,31,185,30,245,31,133,31,104,31,225,31,117,31,163,31,228,31,248,31,145,31,105,31,179,31,40,31,40,30,207,31,49,31,175,31,157,31,157,30,10,31,156,31,172,31,182,31,182,30,106,31,224,31,49,31,48,31,48,30,207,31,234,31,211,31,222,31,220,31,235,31,57,31,1,31,146,31,106,31,2,31,9,31,9,30,164,31,40,31,212,31,70,31,70,30,20,31,208,31,33,31,148,31,252,31,182,31,236,31,42,31,185,31,178,31,207,31,23,31,98,31,98,31,78,31,21,31,21,30,21,29,144,31,131,31,66,31,145,31,191,31,107,31,107,30,107,29,253,31,193,31,80,31,64,31,251,31,16,31,130,31,127,31,110,31,60,31,222,31,2,31,73,31,67,31,2,31,241,31,51,31,183,31,183,30,183,29,183,28,37,31,184,31,134,31,187,31,113,31,67,31,129,31,129,30,240,31,96,31,205,31,229,31,77,31,255,31,51,31,91,31,91,30,91,29,158,31,204,31,160,31,174,31,174,30,214,31,118,31,118,30,200,31,238,31,221,31,221,30,210,31,210,30,135,31,99,31,119,31,101,31,241,31,211,31,5,31,131,31,76,31,125,31,251,31,208,31,136,31,13,31,30,31,64,31,93,31,1,31,63,31,33,31,121,31,50,31,158,31,74,31,161,31,161,30,161,29,110,31,136,31,240,31,240,30,240,29,53,31,111,31,216,31,235,31,235,30,66,31,241,31,164,31,118,31,118,30,134,31,134,30,46,31,42,31,42,30,224,31,224,30,224,29,204,31,180,31,153,31,222,31,149,31,223,31,223,30,62,31,77,31,100,31,100,30,247,31,252,31,252,30,252,29,252,28,82,31,82,30,82,29,228,31,6,31,41,31,84,31,155,31,76,31,21,31,92,31,83,31,103,31,103,30,103,29,103,28,149,31,234,31,130,31,167,31,39,31,127,31,174,31,241,31,31,31,229,31,26,31,197,31,196,31,26,31,26,30,213,31,213,30,23,31,23,30,222,31,247,31,26,31,96,31,192,31,10,31,174,31,67,31,16,31,16,30,3,31,21,31,142,31,142,30,136,31,48,31,48,30,166,31,188,31,73,31,58,31,78,31,243,31,216,31,170,31,174,31,233,31,107,31,170,31,170,30,170,29,111,31,39,31,177,31,254,31,44,31,93,31,93,30,54,31,20,31,113,31,190,31,129,31,31,31,31,30,202,31,233,31,160,31,118,31,2,31,2,30,32,31,247,31,59,31,161,31,200,31,169,31,209,31,232,31,187,31,155,31,36,31,36,30,27,31,137,31,208,31,255,31,13,31,95,31,6,31,143,31,239,31,219,31,202,31,63,31,90,31,109,31,109,30,220,31,101,31,101,30,235,31,235,30,152,31,152,30,141,31,180,31,137,31,141,31,133,31,91,31,169,31,87,31,175,31,175,30,170,31,168,31,168,30,116,31,180,31,135,31,34,31,208,31,42,31,146,31,119,31,56,31,75,31,250,31,250,30,250,29,204,31,8,31,241,31,201,31,201,31,231,31,139,31,249,31,57,31,254,31,254,30,232,31,51,31,144,31,197,31,143,31,143,30,143,29,62,31,62,30,121,31,131,31,131,30,83,31,83,30,70,31,151,31,151,30,152,31,186,31,181,31,245,31,245,30,76,31,195,31,93,31,191,31,162,31,86,31,86,30,86,29,103,31,140,31,183,31,235,31,111,31,18,31,7,31,118,31,251,31,251,30,178,31,178,30,127,31,57,31,88,31,88,30,20,31,86,31,127,31,192,31,131,31,45,31,45,30,62,31,217,31,221,31,221,30,221,29,180,31,214,31,125,31,176,31,56,31,203,31,152,31,183,31,129,31,10,31,234,31,186,31,113,31,113,30,91,31,91,30,91,29,91,28,91,27,79,31,79,30,238,31,238,30,254,31,68,31,242,31,164,31,164,30,187,31,254,31,113,31,113,30,113,29,205,31,205,30,60,31,145,31,110,31,131,31,253,31,105,31,105,30,36,31,78,31,90,31,213,31,111,31,98,31,203,31,12,31,4,31,67,31,173,31,232,31,232,30,232,29,232,28,232,27,36,31,125,31,125,30,125,29,68,31,68,30,157,31,157,30,131,31,246,31,176,31,176,30,176,29,74,31,246,31,220,31,134,31,183,31,112,31,118,31,61,31,138,31,138,30,138,29,15,31,89,31,89,30,223,31,66,31,228,31,86,31,86,30,131,31,227,31,11,31,141,31,253,31,212,31,47,31,247,31,163,31,39,31,229,31,59,31,59,30,254,31,203,31,165,31,165,30,165,31,160,31,119,31,119,30,211,31,252,31,55,31,153,31,91,31,44,31,7,31,20,31,196,31,97,31,97,30,31,31,45,31,45,30,132,31,232,31,68,31,150,31,150,30,28,31,91,31,251,31,251,30,46,31,86,31,94,31,52,31,20,31,20,30,241,31,177,31,177,30,98,31,161,31,113,31,99,31,208,31,156,31,135,31,22,31,73,31,166,31,130,31,130,30,50,31,213,31,201,31,211,31,97,31,97,30,110,31,207,31,111,31,111,30,68,31,4,31,4,30,24,31,130,31,129,31,1,31,17,31,192,31,133,31,116,31,5,31,210,31,102,31,102,30,228,31,35,31,35,30,175,31,61,31,73,31,96,31,147,31,147,30,147,29,52,31,52,30,206,31,97,31,227,31,4,31,91,31,175,31,2,31,117,31,170,31,170,30,153,31,190,31,33,31,72,31,125,31,88,31,182,31,233,31,233,30,251,31,17,31,113,31,246,31,106,31,122,31,174,31,248,31,158,31,88,31,172,31,158,31,172,31,182,31,167,31,160,31,97,31,201,31,194,31,218,31,37,31,185,31,176,31,160,31,160,30,173,31,214,31,132,31,7,31,158,31,8,31,163,31,148,31,96,31,215,31,97,31,97,30,106,31,106,30,106,29,42,31,215,31,104,31,218,31,239,31,91,31,190,31,184,31,90,31,75,31,73,31,79,31,182,31,91,31,24,31,153,31,147,31,253,31,253,30,229,31,229,30,229,29,113,31,151,31,151,30,105,31,135,31,135,30,150,31,151,31,151,30,151,29,241,31,241,30,25,31,230,31,212,31,248,31,233,31,26,31,101,31,141,31,237,31,178,31,198,31,5,31,244,31,120,31,120,30,82,31,82,30,233,31,137,31,175,31,135,31,108,31,59,31,71,31,99,31,99,30,99,29,157,31,71,31,99,31,99,30,204,31,204,30,204,29,98,31,50,31,20,31,171,31,109,31,109,30,204,31,238,31,85,31,130,31,52,31,10,31,10,30,93,31,119,31,6,31,44,31,172,31,71,31,71,30,30,31,132,31,18,31,16,31,44,31,1,31,198,31,198,30,146,31,74,31,74,30,21,31,21,30,167,31,40,31,95,31,95,30,250,31,165,31,147,31,39,31,59,31,203,31,203,30,235,31,229,31,208,31,136,31,169,31,169,30,169,29,93,31,246,31,72,31,185,31,93,31,88,31,222,31,18,31,103,31,22,31,244,31,99,31,2,31,2,30,2,29,162,31,149,31,130,31,111,31,111,30,145,31,142,31,142,30,22,31,106,31,112,31,187,31,51,31,22,31,151,31,88,31,88,30,137,31,231,31,231,30,153,31,186,31,30,31,30,30,30,29,137,31,221,31,221,30,13,31,154,31,138,31,113,31,68,31,224,31,77,31,208,31,58,31,97,31,73,31,73,30,73,29,173,31,250,31,176,31,250,31,159,31,192,31,117,31,144,31,20,31,246,31,149,31,149,30,149,29,201,31,201,30,201,29,5,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
