-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_526 is
end project_tb_526;

architecture project_tb_arch_526 of project_tb_526 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 441;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (21,0,0,0,37,0,44,0,225,0,231,0,95,0,0,0,163,0,131,0,133,0,0,0,228,0,63,0,0,0,19,0,0,0,0,0,30,0,0,0,244,0,83,0,198,0,33,0,201,0,13,0,184,0,62,0,110,0,56,0,0,0,147,0,180,0,62,0,0,0,206,0,87,0,121,0,246,0,247,0,123,0,253,0,181,0,126,0,70,0,162,0,241,0,142,0,55,0,11,0,69,0,0,0,0,0,210,0,0,0,255,0,47,0,0,0,4,0,0,0,19,0,172,0,73,0,116,0,30,0,153,0,67,0,120,0,219,0,252,0,12,0,0,0,171,0,0,0,180,0,81,0,193,0,58,0,177,0,145,0,142,0,0,0,48,0,112,0,220,0,0,0,45,0,252,0,0,0,66,0,0,0,82,0,104,0,168,0,216,0,0,0,23,0,84,0,0,0,110,0,0,0,233,0,133,0,208,0,0,0,177,0,180,0,82,0,205,0,111,0,0,0,94,0,160,0,176,0,0,0,140,0,68,0,74,0,255,0,51,0,0,0,21,0,28,0,80,0,0,0,75,0,169,0,0,0,91,0,175,0,242,0,35,0,129,0,0,0,48,0,0,0,0,0,189,0,28,0,41,0,32,0,76,0,130,0,86,0,160,0,28,0,152,0,242,0,221,0,252,0,0,0,128,0,0,0,0,0,136,0,60,0,202,0,183,0,58,0,57,0,110,0,101,0,66,0,37,0,165,0,125,0,177,0,247,0,84,0,63,0,22,0,63,0,248,0,166,0,18,0,211,0,18,0,1,0,0,0,141,0,0,0,0,0,149,0,178,0,110,0,68,0,101,0,102,0,55,0,251,0,0,0,174,0,206,0,0,0,0,0,180,0,38,0,7,0,0,0,143,0,83,0,255,0,66,0,75,0,98,0,182,0,50,0,2,0,0,0,210,0,88,0,183,0,254,0,0,0,0,0,137,0,1,0,231,0,38,0,51,0,0,0,146,0,171,0,216,0,83,0,0,0,157,0,24,0,127,0,99,0,0,0,6,0,52,0,219,0,178,0,51,0,0,0,129,0,38,0,255,0,96,0,146,0,0,0,0,0,117,0,0,0,0,0,245,0,197,0,0,0,5,0,19,0,0,0,126,0,0,0,25,0,154,0,0,0,26,0,72,0,208,0,0,0,23,0,0,0,7,0,13,0,14,0,3,0,0,0,136,0,212,0,155,0,61,0,0,0,0,0,100,0,0,0,16,0,160,0,120,0,110,0,204,0,0,0,111,0,168,0,31,0,35,0,0,0,229,0,0,0,219,0,0,0,132,0,0,0,238,0,0,0,115,0,0,0,231,0,202,0,0,0,40,0,212,0,84,0,228,0,60,0,155,0,218,0,0,0,124,0,0,0,0,0,156,0,168,0,0,0,19,0,122,0,83,0,241,0,181,0,115,0,135,0,229,0,121,0,239,0,64,0,0,0,127,0,154,0,126,0,0,0,0,0,202,0,74,0,93,0,224,0,127,0,12,0,235,0,96,0,86,0,149,0,0,0,133,0,216,0,86,0,22,0,87,0,151,0,163,0,56,0,0,0,68,0,81,0,239,0,154,0,217,0,234,0,82,0,130,0,147,0,91,0,160,0,0,0,135,0,157,0,230,0,0,0,185,0,57,0,70,0,0,0,173,0,3,0,131,0,78,0,0,0,100,0,80,0,118,0,120,0,26,0,80,0,11,0,208,0,182,0,0,0,143,0,0,0,75,0,15,0,214,0,134,0,0,0,144,0,144,0,0,0,156,0,145,0,108,0,242,0,148,0,0,0,47,0,0,0,0,0,245,0,0,0,134,0,210,0,211,0,95,0,247,0,86,0,52,0,61,0,100,0,11,0,65,0,131,0,126,0,116,0,0,0,52,0,0,0,159,0,0,0,102,0,76,0,136,0,253,0,15,0,4,0,156,0,8,0,0,0,0,0,238,0,145,0,174,0,181,0);
signal scenario_full  : scenario_type := (21,31,21,30,37,31,44,31,225,31,231,31,95,31,95,30,163,31,131,31,133,31,133,30,228,31,63,31,63,30,19,31,19,30,19,29,30,31,30,30,244,31,83,31,198,31,33,31,201,31,13,31,184,31,62,31,110,31,56,31,56,30,147,31,180,31,62,31,62,30,206,31,87,31,121,31,246,31,247,31,123,31,253,31,181,31,126,31,70,31,162,31,241,31,142,31,55,31,11,31,69,31,69,30,69,29,210,31,210,30,255,31,47,31,47,30,4,31,4,30,19,31,172,31,73,31,116,31,30,31,153,31,67,31,120,31,219,31,252,31,12,31,12,30,171,31,171,30,180,31,81,31,193,31,58,31,177,31,145,31,142,31,142,30,48,31,112,31,220,31,220,30,45,31,252,31,252,30,66,31,66,30,82,31,104,31,168,31,216,31,216,30,23,31,84,31,84,30,110,31,110,30,233,31,133,31,208,31,208,30,177,31,180,31,82,31,205,31,111,31,111,30,94,31,160,31,176,31,176,30,140,31,68,31,74,31,255,31,51,31,51,30,21,31,28,31,80,31,80,30,75,31,169,31,169,30,91,31,175,31,242,31,35,31,129,31,129,30,48,31,48,30,48,29,189,31,28,31,41,31,32,31,76,31,130,31,86,31,160,31,28,31,152,31,242,31,221,31,252,31,252,30,128,31,128,30,128,29,136,31,60,31,202,31,183,31,58,31,57,31,110,31,101,31,66,31,37,31,165,31,125,31,177,31,247,31,84,31,63,31,22,31,63,31,248,31,166,31,18,31,211,31,18,31,1,31,1,30,141,31,141,30,141,29,149,31,178,31,110,31,68,31,101,31,102,31,55,31,251,31,251,30,174,31,206,31,206,30,206,29,180,31,38,31,7,31,7,30,143,31,83,31,255,31,66,31,75,31,98,31,182,31,50,31,2,31,2,30,210,31,88,31,183,31,254,31,254,30,254,29,137,31,1,31,231,31,38,31,51,31,51,30,146,31,171,31,216,31,83,31,83,30,157,31,24,31,127,31,99,31,99,30,6,31,52,31,219,31,178,31,51,31,51,30,129,31,38,31,255,31,96,31,146,31,146,30,146,29,117,31,117,30,117,29,245,31,197,31,197,30,5,31,19,31,19,30,126,31,126,30,25,31,154,31,154,30,26,31,72,31,208,31,208,30,23,31,23,30,7,31,13,31,14,31,3,31,3,30,136,31,212,31,155,31,61,31,61,30,61,29,100,31,100,30,16,31,160,31,120,31,110,31,204,31,204,30,111,31,168,31,31,31,35,31,35,30,229,31,229,30,219,31,219,30,132,31,132,30,238,31,238,30,115,31,115,30,231,31,202,31,202,30,40,31,212,31,84,31,228,31,60,31,155,31,218,31,218,30,124,31,124,30,124,29,156,31,168,31,168,30,19,31,122,31,83,31,241,31,181,31,115,31,135,31,229,31,121,31,239,31,64,31,64,30,127,31,154,31,126,31,126,30,126,29,202,31,74,31,93,31,224,31,127,31,12,31,235,31,96,31,86,31,149,31,149,30,133,31,216,31,86,31,22,31,87,31,151,31,163,31,56,31,56,30,68,31,81,31,239,31,154,31,217,31,234,31,82,31,130,31,147,31,91,31,160,31,160,30,135,31,157,31,230,31,230,30,185,31,57,31,70,31,70,30,173,31,3,31,131,31,78,31,78,30,100,31,80,31,118,31,120,31,26,31,80,31,11,31,208,31,182,31,182,30,143,31,143,30,75,31,15,31,214,31,134,31,134,30,144,31,144,31,144,30,156,31,145,31,108,31,242,31,148,31,148,30,47,31,47,30,47,29,245,31,245,30,134,31,210,31,211,31,95,31,247,31,86,31,52,31,61,31,100,31,11,31,65,31,131,31,126,31,116,31,116,30,52,31,52,30,159,31,159,30,102,31,76,31,136,31,253,31,15,31,4,31,156,31,8,31,8,30,8,29,238,31,145,31,174,31,181,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
