-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_349 is
end project_tb_349;

architecture project_tb_arch_349 of project_tb_349 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 302;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (187,0,184,0,224,0,94,0,83,0,18,0,56,0,152,0,254,0,22,0,0,0,44,0,52,0,119,0,240,0,98,0,110,0,143,0,0,0,252,0,240,0,123,0,210,0,0,0,149,0,0,0,0,0,58,0,112,0,67,0,147,0,212,0,0,0,0,0,213,0,0,0,176,0,229,0,115,0,0,0,111,0,158,0,0,0,131,0,34,0,171,0,106,0,56,0,0,0,0,0,0,0,22,0,0,0,122,0,47,0,148,0,150,0,0,0,49,0,0,0,209,0,19,0,110,0,39,0,186,0,42,0,137,0,108,0,0,0,62,0,0,0,0,0,0,0,163,0,0,0,0,0,111,0,95,0,0,0,199,0,0,0,62,0,77,0,123,0,0,0,172,0,190,0,42,0,182,0,21,0,0,0,160,0,158,0,0,0,0,0,241,0,196,0,189,0,142,0,177,0,181,0,16,0,166,0,32,0,94,0,0,0,207,0,73,0,225,0,0,0,206,0,178,0,0,0,179,0,194,0,6,0,97,0,0,0,130,0,45,0,201,0,0,0,0,0,166,0,213,0,200,0,185,0,0,0,224,0,136,0,175,0,37,0,18,0,51,0,85,0,35,0,146,0,250,0,27,0,98,0,58,0,0,0,95,0,152,0,190,0,113,0,226,0,148,0,0,0,1,0,235,0,0,0,193,0,116,0,185,0,94,0,122,0,119,0,117,0,215,0,0,0,185,0,0,0,218,0,135,0,211,0,253,0,199,0,67,0,187,0,208,0,0,0,142,0,83,0,121,0,41,0,79,0,0,0,112,0,135,0,167,0,110,0,106,0,0,0,0,0,128,0,90,0,0,0,75,0,0,0,39,0,200,0,225,0,0,0,0,0,155,0,164,0,16,0,254,0,25,0,0,0,196,0,108,0,76,0,0,0,178,0,169,0,42,0,3,0,0,0,218,0,205,0,125,0,127,0,12,0,59,0,127,0,189,0,243,0,0,0,0,0,62,0,76,0,38,0,231,0,10,0,166,0,196,0,72,0,112,0,141,0,0,0,16,0,175,0,97,0,0,0,96,0,203,0,227,0,123,0,0,0,136,0,86,0,131,0,0,0,109,0,239,0,195,0,152,0,4,0,195,0,148,0,157,0,131,0,243,0,0,0,116,0,0,0,0,0,157,0,136,0,178,0,0,0,9,0,91,0,77,0,85,0,18,0,211,0,5,0,0,0,133,0,0,0,211,0,110,0,82,0,252,0,105,0,0,0,120,0,62,0,0,0,201,0,181,0,109,0,0,0,0,0,128,0,36,0,70,0,178,0,64,0,214,0,67,0,165,0,206,0,0,0,88,0,237,0,122,0,77,0,0,0);
signal scenario_full  : scenario_type := (187,31,184,31,224,31,94,31,83,31,18,31,56,31,152,31,254,31,22,31,22,30,44,31,52,31,119,31,240,31,98,31,110,31,143,31,143,30,252,31,240,31,123,31,210,31,210,30,149,31,149,30,149,29,58,31,112,31,67,31,147,31,212,31,212,30,212,29,213,31,213,30,176,31,229,31,115,31,115,30,111,31,158,31,158,30,131,31,34,31,171,31,106,31,56,31,56,30,56,29,56,28,22,31,22,30,122,31,47,31,148,31,150,31,150,30,49,31,49,30,209,31,19,31,110,31,39,31,186,31,42,31,137,31,108,31,108,30,62,31,62,30,62,29,62,28,163,31,163,30,163,29,111,31,95,31,95,30,199,31,199,30,62,31,77,31,123,31,123,30,172,31,190,31,42,31,182,31,21,31,21,30,160,31,158,31,158,30,158,29,241,31,196,31,189,31,142,31,177,31,181,31,16,31,166,31,32,31,94,31,94,30,207,31,73,31,225,31,225,30,206,31,178,31,178,30,179,31,194,31,6,31,97,31,97,30,130,31,45,31,201,31,201,30,201,29,166,31,213,31,200,31,185,31,185,30,224,31,136,31,175,31,37,31,18,31,51,31,85,31,35,31,146,31,250,31,27,31,98,31,58,31,58,30,95,31,152,31,190,31,113,31,226,31,148,31,148,30,1,31,235,31,235,30,193,31,116,31,185,31,94,31,122,31,119,31,117,31,215,31,215,30,185,31,185,30,218,31,135,31,211,31,253,31,199,31,67,31,187,31,208,31,208,30,142,31,83,31,121,31,41,31,79,31,79,30,112,31,135,31,167,31,110,31,106,31,106,30,106,29,128,31,90,31,90,30,75,31,75,30,39,31,200,31,225,31,225,30,225,29,155,31,164,31,16,31,254,31,25,31,25,30,196,31,108,31,76,31,76,30,178,31,169,31,42,31,3,31,3,30,218,31,205,31,125,31,127,31,12,31,59,31,127,31,189,31,243,31,243,30,243,29,62,31,76,31,38,31,231,31,10,31,166,31,196,31,72,31,112,31,141,31,141,30,16,31,175,31,97,31,97,30,96,31,203,31,227,31,123,31,123,30,136,31,86,31,131,31,131,30,109,31,239,31,195,31,152,31,4,31,195,31,148,31,157,31,131,31,243,31,243,30,116,31,116,30,116,29,157,31,136,31,178,31,178,30,9,31,91,31,77,31,85,31,18,31,211,31,5,31,5,30,133,31,133,30,211,31,110,31,82,31,252,31,105,31,105,30,120,31,62,31,62,30,201,31,181,31,109,31,109,30,109,29,128,31,36,31,70,31,178,31,64,31,214,31,67,31,165,31,206,31,206,30,88,31,237,31,122,31,77,31,77,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
