-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1003;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (133,0,202,0,0,0,232,0,77,0,145,0,65,0,250,0,221,0,221,0,34,0,0,0,194,0,226,0,106,0,181,0,43,0,0,0,0,0,65,0,52,0,159,0,0,0,18,0,40,0,0,0,9,0,0,0,0,0,35,0,81,0,0,0,199,0,0,0,132,0,218,0,0,0,247,0,182,0,93,0,38,0,202,0,0,0,159,0,111,0,175,0,45,0,22,0,253,0,3,0,0,0,0,0,237,0,222,0,90,0,0,0,223,0,13,0,7,0,188,0,30,0,98,0,0,0,123,0,89,0,219,0,17,0,196,0,99,0,88,0,102,0,166,0,111,0,0,0,36,0,97,0,0,0,215,0,152,0,132,0,69,0,240,0,215,0,74,0,24,0,105,0,0,0,221,0,173,0,4,0,0,0,196,0,68,0,50,0,0,0,173,0,57,0,57,0,172,0,44,0,56,0,223,0,49,0,11,0,105,0,162,0,0,0,136,0,220,0,28,0,96,0,15,0,162,0,0,0,121,0,174,0,88,0,151,0,127,0,236,0,0,0,43,0,240,0,246,0,120,0,181,0,92,0,190,0,43,0,218,0,223,0,36,0,92,0,54,0,88,0,88,0,0,0,147,0,65,0,33,0,219,0,175,0,8,0,64,0,79,0,216,0,0,0,188,0,243,0,206,0,0,0,84,0,112,0,45,0,85,0,0,0,158,0,33,0,0,0,91,0,178,0,20,0,154,0,0,0,235,0,0,0,6,0,57,0,120,0,211,0,199,0,189,0,32,0,108,0,4,0,0,0,181,0,72,0,143,0,82,0,2,0,9,0,198,0,93,0,233,0,168,0,240,0,241,0,69,0,75,0,170,0,140,0,232,0,30,0,64,0,124,0,0,0,145,0,28,0,57,0,209,0,0,0,0,0,134,0,0,0,137,0,59,0,28,0,74,0,171,0,131,0,26,0,204,0,241,0,62,0,248,0,202,0,132,0,143,0,241,0,231,0,182,0,251,0,189,0,107,0,14,0,111,0,143,0,173,0,0,0,0,0,249,0,146,0,166,0,134,0,6,0,93,0,99,0,75,0,75,0,221,0,6,0,45,0,17,0,0,0,178,0,98,0,0,0,103,0,0,0,63,0,126,0,77,0,186,0,118,0,0,0,0,0,78,0,0,0,0,0,151,0,57,0,242,0,178,0,125,0,0,0,78,0,21,0,0,0,0,0,65,0,142,0,0,0,57,0,121,0,0,0,244,0,188,0,32,0,41,0,246,0,182,0,34,0,216,0,0,0,239,0,146,0,0,0,75,0,190,0,90,0,151,0,137,0,0,0,0,0,111,0,0,0,255,0,247,0,27,0,20,0,227,0,31,0,159,0,201,0,0,0,59,0,25,0,89,0,149,0,9,0,225,0,127,0,31,0,171,0,70,0,20,0,0,0,150,0,155,0,255,0,0,0,126,0,0,0,162,0,238,0,105,0,0,0,81,0,178,0,67,0,175,0,220,0,105,0,182,0,79,0,144,0,0,0,198,0,20,0,81,0,206,0,71,0,1,0,88,0,221,0,187,0,0,0,0,0,121,0,0,0,89,0,201,0,20,0,84,0,105,0,28,0,198,0,0,0,133,0,0,0,0,0,0,0,49,0,216,0,212,0,248,0,126,0,1,0,177,0,226,0,6,0,0,0,235,0,237,0,0,0,35,0,0,0,0,0,56,0,0,0,175,0,136,0,173,0,175,0,254,0,42,0,42,0,167,0,0,0,6,0,0,0,76,0,101,0,33,0,110,0,238,0,93,0,47,0,199,0,236,0,78,0,96,0,123,0,243,0,0,0,91,0,182,0,0,0,143,0,56,0,208,0,11,0,0,0,126,0,159,0,0,0,187,0,0,0,0,0,40,0,227,0,1,0,16,0,183,0,198,0,73,0,183,0,0,0,234,0,150,0,0,0,51,0,50,0,128,0,0,0,163,0,71,0,211,0,103,0,88,0,35,0,71,0,65,0,54,0,115,0,204,0,97,0,177,0,70,0,118,0,143,0,227,0,132,0,242,0,226,0,244,0,37,0,172,0,48,0,125,0,113,0,243,0,69,0,235,0,0,0,0,0,0,0,27,0,51,0,57,0,75,0,0,0,19,0,176,0,85,0,0,0,119,0,0,0,40,0,87,0,0,0,107,0,0,0,146,0,0,0,234,0,198,0,64,0,243,0,0,0,0,0,219,0,52,0,0,0,89,0,248,0,0,0,23,0,49,0,51,0,36,0,252,0,135,0,129,0,104,0,0,0,20,0,251,0,242,0,27,0,194,0,56,0,110,0,32,0,133,0,0,0,113,0,149,0,0,0,14,0,119,0,36,0,62,0,147,0,220,0,109,0,32,0,148,0,169,0,129,0,158,0,0,0,0,0,249,0,134,0,0,0,72,0,0,0,244,0,13,0,41,0,215,0,43,0,0,0,239,0,213,0,64,0,149,0,0,0,40,0,196,0,185,0,45,0,166,0,175,0,120,0,245,0,167,0,241,0,128,0,49,0,50,0,131,0,0,0,17,0,202,0,53,0,182,0,200,0,189,0,31,0,176,0,123,0,0,0,156,0,123,0,235,0,243,0,227,0,230,0,98,0,253,0,0,0,219,0,0,0,68,0,64,0,36,0,189,0,20,0,140,0,39,0,90,0,191,0,16,0,0,0,213,0,21,0,79,0,59,0,228,0,193,0,244,0,114,0,108,0,177,0,33,0,200,0,0,0,214,0,0,0,0,0,102,0,0,0,242,0,58,0,0,0,48,0,76,0,235,0,138,0,180,0,0,0,97,0,79,0,110,0,9,0,89,0,184,0,61,0,226,0,156,0,0,0,157,0,174,0,26,0,26,0,190,0,46,0,52,0,102,0,0,0,111,0,156,0,115,0,100,0,162,0,3,0,189,0,82,0,76,0,219,0,31,0,134,0,0,0,98,0,0,0,94,0,70,0,0,0,199,0,0,0,47,0,13,0,210,0,0,0,99,0,50,0,109,0,67,0,0,0,183,0,0,0,186,0,178,0,216,0,0,0,63,0,89,0,0,0,186,0,0,0,54,0,245,0,0,0,162,0,156,0,121,0,187,0,0,0,148,0,194,0,0,0,247,0,27,0,40,0,132,0,0,0,0,0,176,0,61,0,158,0,15,0,164,0,221,0,152,0,161,0,6,0,83,0,132,0,5,0,0,0,224,0,36,0,0,0,54,0,0,0,8,0,6,0,67,0,0,0,153,0,0,0,164,0,189,0,0,0,250,0,45,0,87,0,219,0,167,0,209,0,34,0,0,0,132,0,135,0,0,0,49,0,115,0,249,0,58,0,0,0,50,0,55,0,152,0,0,0,130,0,54,0,17,0,0,0,171,0,62,0,162,0,0,0,165,0,0,0,49,0,249,0,148,0,234,0,155,0,67,0,113,0,201,0,0,0,160,0,0,0,0,0,0,0,186,0,186,0,34,0,115,0,133,0,214,0,38,0,0,0,248,0,0,0,197,0,51,0,137,0,67,0,250,0,249,0,28,0,61,0,71,0,0,0,230,0,52,0,82,0,0,0,123,0,26,0,170,0,0,0,228,0,147,0,71,0,122,0,176,0,142,0,251,0,160,0,72,0,83,0,204,0,119,0,0,0,0,0,61,0,102,0,43,0,250,0,181,0,125,0,0,0,221,0,80,0,0,0,178,0,0,0,210,0,134,0,0,0,27,0,251,0,42,0,231,0,0,0,7,0,112,0,228,0,59,0,116,0,118,0,52,0,83,0,195,0,13,0,0,0,88,0,15,0,157,0,57,0,0,0,101,0,179,0,0,0,134,0,253,0,105,0,0,0,145,0,9,0,115,0,121,0,221,0,155,0,0,0,145,0,214,0,8,0,210,0,0,0,201,0,213,0,107,0,0,0,88,0,244,0,181,0,109,0,80,0,190,0,217,0,0,0,97,0,0,0,155,0,224,0,0,0,0,0,0,0,169,0,172,0,0,0,220,0,0,0,0,0,16,0,0,0,166,0,140,0,20,0,0,0,88,0,0,0,163,0,52,0,0,0,0,0,0,0,41,0,18,0,129,0,90,0,0,0,0,0,162,0,205,0,239,0,174,0,0,0,175,0,0,0,45,0,125,0,83,0,0,0,51,0,166,0,0,0,224,0,143,0,23,0,0,0,3,0,0,0,0,0,36,0,226,0,0,0,220,0,61,0,225,0,173,0,0,0,202,0,92,0,0,0,10,0,175,0,246,0,156,0,0,0,0,0,85,0,175,0,0,0,154,0,20,0,117,0,236,0,248,0,157,0,0,0,202,0,233,0,94,0,85,0,250,0,0,0,131,0,59,0,140,0,69,0,240,0,32,0,150,0,66,0,254,0,0,0,11,0,6,0,238,0,104,0,183,0,138,0,52,0,0,0,0,0,0,0,4,0,54,0,0,0,2,0,120,0,249,0,215,0,0,0,15,0,136,0,152,0,79,0,227,0,237,0,136,0,0,0,1,0,226,0);
signal scenario_full  : scenario_type := (133,31,202,31,202,30,232,31,77,31,145,31,65,31,250,31,221,31,221,31,34,31,34,30,194,31,226,31,106,31,181,31,43,31,43,30,43,29,65,31,52,31,159,31,159,30,18,31,40,31,40,30,9,31,9,30,9,29,35,31,81,31,81,30,199,31,199,30,132,31,218,31,218,30,247,31,182,31,93,31,38,31,202,31,202,30,159,31,111,31,175,31,45,31,22,31,253,31,3,31,3,30,3,29,237,31,222,31,90,31,90,30,223,31,13,31,7,31,188,31,30,31,98,31,98,30,123,31,89,31,219,31,17,31,196,31,99,31,88,31,102,31,166,31,111,31,111,30,36,31,97,31,97,30,215,31,152,31,132,31,69,31,240,31,215,31,74,31,24,31,105,31,105,30,221,31,173,31,4,31,4,30,196,31,68,31,50,31,50,30,173,31,57,31,57,31,172,31,44,31,56,31,223,31,49,31,11,31,105,31,162,31,162,30,136,31,220,31,28,31,96,31,15,31,162,31,162,30,121,31,174,31,88,31,151,31,127,31,236,31,236,30,43,31,240,31,246,31,120,31,181,31,92,31,190,31,43,31,218,31,223,31,36,31,92,31,54,31,88,31,88,31,88,30,147,31,65,31,33,31,219,31,175,31,8,31,64,31,79,31,216,31,216,30,188,31,243,31,206,31,206,30,84,31,112,31,45,31,85,31,85,30,158,31,33,31,33,30,91,31,178,31,20,31,154,31,154,30,235,31,235,30,6,31,57,31,120,31,211,31,199,31,189,31,32,31,108,31,4,31,4,30,181,31,72,31,143,31,82,31,2,31,9,31,198,31,93,31,233,31,168,31,240,31,241,31,69,31,75,31,170,31,140,31,232,31,30,31,64,31,124,31,124,30,145,31,28,31,57,31,209,31,209,30,209,29,134,31,134,30,137,31,59,31,28,31,74,31,171,31,131,31,26,31,204,31,241,31,62,31,248,31,202,31,132,31,143,31,241,31,231,31,182,31,251,31,189,31,107,31,14,31,111,31,143,31,173,31,173,30,173,29,249,31,146,31,166,31,134,31,6,31,93,31,99,31,75,31,75,31,221,31,6,31,45,31,17,31,17,30,178,31,98,31,98,30,103,31,103,30,63,31,126,31,77,31,186,31,118,31,118,30,118,29,78,31,78,30,78,29,151,31,57,31,242,31,178,31,125,31,125,30,78,31,21,31,21,30,21,29,65,31,142,31,142,30,57,31,121,31,121,30,244,31,188,31,32,31,41,31,246,31,182,31,34,31,216,31,216,30,239,31,146,31,146,30,75,31,190,31,90,31,151,31,137,31,137,30,137,29,111,31,111,30,255,31,247,31,27,31,20,31,227,31,31,31,159,31,201,31,201,30,59,31,25,31,89,31,149,31,9,31,225,31,127,31,31,31,171,31,70,31,20,31,20,30,150,31,155,31,255,31,255,30,126,31,126,30,162,31,238,31,105,31,105,30,81,31,178,31,67,31,175,31,220,31,105,31,182,31,79,31,144,31,144,30,198,31,20,31,81,31,206,31,71,31,1,31,88,31,221,31,187,31,187,30,187,29,121,31,121,30,89,31,201,31,20,31,84,31,105,31,28,31,198,31,198,30,133,31,133,30,133,29,133,28,49,31,216,31,212,31,248,31,126,31,1,31,177,31,226,31,6,31,6,30,235,31,237,31,237,30,35,31,35,30,35,29,56,31,56,30,175,31,136,31,173,31,175,31,254,31,42,31,42,31,167,31,167,30,6,31,6,30,76,31,101,31,33,31,110,31,238,31,93,31,47,31,199,31,236,31,78,31,96,31,123,31,243,31,243,30,91,31,182,31,182,30,143,31,56,31,208,31,11,31,11,30,126,31,159,31,159,30,187,31,187,30,187,29,40,31,227,31,1,31,16,31,183,31,198,31,73,31,183,31,183,30,234,31,150,31,150,30,51,31,50,31,128,31,128,30,163,31,71,31,211,31,103,31,88,31,35,31,71,31,65,31,54,31,115,31,204,31,97,31,177,31,70,31,118,31,143,31,227,31,132,31,242,31,226,31,244,31,37,31,172,31,48,31,125,31,113,31,243,31,69,31,235,31,235,30,235,29,235,28,27,31,51,31,57,31,75,31,75,30,19,31,176,31,85,31,85,30,119,31,119,30,40,31,87,31,87,30,107,31,107,30,146,31,146,30,234,31,198,31,64,31,243,31,243,30,243,29,219,31,52,31,52,30,89,31,248,31,248,30,23,31,49,31,51,31,36,31,252,31,135,31,129,31,104,31,104,30,20,31,251,31,242,31,27,31,194,31,56,31,110,31,32,31,133,31,133,30,113,31,149,31,149,30,14,31,119,31,36,31,62,31,147,31,220,31,109,31,32,31,148,31,169,31,129,31,158,31,158,30,158,29,249,31,134,31,134,30,72,31,72,30,244,31,13,31,41,31,215,31,43,31,43,30,239,31,213,31,64,31,149,31,149,30,40,31,196,31,185,31,45,31,166,31,175,31,120,31,245,31,167,31,241,31,128,31,49,31,50,31,131,31,131,30,17,31,202,31,53,31,182,31,200,31,189,31,31,31,176,31,123,31,123,30,156,31,123,31,235,31,243,31,227,31,230,31,98,31,253,31,253,30,219,31,219,30,68,31,64,31,36,31,189,31,20,31,140,31,39,31,90,31,191,31,16,31,16,30,213,31,21,31,79,31,59,31,228,31,193,31,244,31,114,31,108,31,177,31,33,31,200,31,200,30,214,31,214,30,214,29,102,31,102,30,242,31,58,31,58,30,48,31,76,31,235,31,138,31,180,31,180,30,97,31,79,31,110,31,9,31,89,31,184,31,61,31,226,31,156,31,156,30,157,31,174,31,26,31,26,31,190,31,46,31,52,31,102,31,102,30,111,31,156,31,115,31,100,31,162,31,3,31,189,31,82,31,76,31,219,31,31,31,134,31,134,30,98,31,98,30,94,31,70,31,70,30,199,31,199,30,47,31,13,31,210,31,210,30,99,31,50,31,109,31,67,31,67,30,183,31,183,30,186,31,178,31,216,31,216,30,63,31,89,31,89,30,186,31,186,30,54,31,245,31,245,30,162,31,156,31,121,31,187,31,187,30,148,31,194,31,194,30,247,31,27,31,40,31,132,31,132,30,132,29,176,31,61,31,158,31,15,31,164,31,221,31,152,31,161,31,6,31,83,31,132,31,5,31,5,30,224,31,36,31,36,30,54,31,54,30,8,31,6,31,67,31,67,30,153,31,153,30,164,31,189,31,189,30,250,31,45,31,87,31,219,31,167,31,209,31,34,31,34,30,132,31,135,31,135,30,49,31,115,31,249,31,58,31,58,30,50,31,55,31,152,31,152,30,130,31,54,31,17,31,17,30,171,31,62,31,162,31,162,30,165,31,165,30,49,31,249,31,148,31,234,31,155,31,67,31,113,31,201,31,201,30,160,31,160,30,160,29,160,28,186,31,186,31,34,31,115,31,133,31,214,31,38,31,38,30,248,31,248,30,197,31,51,31,137,31,67,31,250,31,249,31,28,31,61,31,71,31,71,30,230,31,52,31,82,31,82,30,123,31,26,31,170,31,170,30,228,31,147,31,71,31,122,31,176,31,142,31,251,31,160,31,72,31,83,31,204,31,119,31,119,30,119,29,61,31,102,31,43,31,250,31,181,31,125,31,125,30,221,31,80,31,80,30,178,31,178,30,210,31,134,31,134,30,27,31,251,31,42,31,231,31,231,30,7,31,112,31,228,31,59,31,116,31,118,31,52,31,83,31,195,31,13,31,13,30,88,31,15,31,157,31,57,31,57,30,101,31,179,31,179,30,134,31,253,31,105,31,105,30,145,31,9,31,115,31,121,31,221,31,155,31,155,30,145,31,214,31,8,31,210,31,210,30,201,31,213,31,107,31,107,30,88,31,244,31,181,31,109,31,80,31,190,31,217,31,217,30,97,31,97,30,155,31,224,31,224,30,224,29,224,28,169,31,172,31,172,30,220,31,220,30,220,29,16,31,16,30,166,31,140,31,20,31,20,30,88,31,88,30,163,31,52,31,52,30,52,29,52,28,41,31,18,31,129,31,90,31,90,30,90,29,162,31,205,31,239,31,174,31,174,30,175,31,175,30,45,31,125,31,83,31,83,30,51,31,166,31,166,30,224,31,143,31,23,31,23,30,3,31,3,30,3,29,36,31,226,31,226,30,220,31,61,31,225,31,173,31,173,30,202,31,92,31,92,30,10,31,175,31,246,31,156,31,156,30,156,29,85,31,175,31,175,30,154,31,20,31,117,31,236,31,248,31,157,31,157,30,202,31,233,31,94,31,85,31,250,31,250,30,131,31,59,31,140,31,69,31,240,31,32,31,150,31,66,31,254,31,254,30,11,31,6,31,238,31,104,31,183,31,138,31,52,31,52,30,52,29,52,28,4,31,54,31,54,30,2,31,120,31,249,31,215,31,215,30,15,31,136,31,152,31,79,31,227,31,237,31,136,31,136,30,1,31,226,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
