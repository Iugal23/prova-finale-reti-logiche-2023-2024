-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 402;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,113,0,1,0,215,0,85,0,84,0,35,0,46,0,0,0,238,0,12,0,40,0,0,0,109,0,161,0,0,0,152,0,0,0,193,0,137,0,22,0,0,0,0,0,28,0,64,0,227,0,117,0,199,0,47,0,235,0,219,0,20,0,45,0,166,0,0,0,0,0,106,0,193,0,9,0,172,0,103,0,250,0,255,0,52,0,0,0,19,0,186,0,23,0,221,0,0,0,161,0,252,0,188,0,0,0,196,0,0,0,0,0,8,0,247,0,16,0,168,0,170,0,155,0,20,0,135,0,147,0,17,0,0,0,190,0,251,0,137,0,119,0,128,0,0,0,0,0,173,0,205,0,0,0,206,0,145,0,99,0,0,0,131,0,11,0,74,0,219,0,44,0,229,0,231,0,198,0,166,0,0,0,0,0,119,0,79,0,228,0,0,0,59,0,30,0,158,0,114,0,165,0,1,0,50,0,48,0,164,0,83,0,89,0,58,0,0,0,148,0,0,0,120,0,0,0,206,0,235,0,220,0,0,0,0,0,70,0,148,0,0,0,0,0,190,0,58,0,245,0,237,0,0,0,33,0,126,0,160,0,0,0,235,0,10,0,114,0,0,0,160,0,6,0,87,0,78,0,226,0,115,0,111,0,39,0,51,0,61,0,0,0,38,0,204,0,23,0,135,0,132,0,205,0,58,0,138,0,0,0,55,0,244,0,73,0,134,0,157,0,175,0,154,0,0,0,33,0,98,0,247,0,0,0,145,0,160,0,71,0,68,0,120,0,55,0,0,0,212,0,69,0,127,0,106,0,0,0,0,0,253,0,0,0,242,0,51,0,56,0,163,0,94,0,86,0,9,0,4,0,219,0,177,0,160,0,0,0,174,0,0,0,181,0,164,0,131,0,0,0,90,0,42,0,101,0,133,0,214,0,0,0,115,0,60,0,107,0,0,0,141,0,161,0,251,0,63,0,0,0,219,0,0,0,0,0,135,0,0,0,119,0,232,0,100,0,8,0,50,0,31,0,208,0,78,0,0,0,205,0,8,0,88,0,0,0,123,0,39,0,229,0,243,0,31,0,20,0,0,0,203,0,46,0,151,0,49,0,188,0,88,0,9,0,9,0,113,0,156,0,233,0,105,0,0,0,208,0,217,0,45,0,113,0,50,0,11,0,250,0,199,0,91,0,201,0,242,0,235,0,0,0,8,0,231,0,249,0,0,0,0,0,0,0,0,0,119,0,0,0,211,0,0,0,189,0,10,0,92,0,174,0,0,0,60,0,117,0,253,0,150,0,132,0,16,0,72,0,69,0,0,0,89,0,43,0,0,0,114,0,94,0,16,0,26,0,160,0,162,0,122,0,65,0,143,0,248,0,191,0,17,0,166,0,8,0,0,0,0,0,172,0,114,0,0,0,211,0,209,0,0,0,4,0,0,0,51,0,28,0,114,0,222,0,250,0,9,0,123,0,229,0,130,0,81,0,90,0,118,0,67,0,0,0,250,0,135,0,22,0,104,0,98,0,76,0,40,0,184,0,0,0,98,0,121,0,106,0,0,0,3,0,119,0,114,0,0,0,5,0,231,0,121,0,138,0,125,0,6,0,0,0,107,0,224,0,18,0,0,0,102,0,0,0,94,0,163,0,251,0,28,0,233,0,143,0,86,0,135,0,246,0,220,0,197,0,36,0,0,0,211,0,153,0,0,0,129,0,112,0,0,0,208,0,0,0,188,0,46,0,23,0,0,0,68,0,0,0,0,0,172,0,159,0,0,0,0,0,0,0,251,0,0,0,192,0,12,0,246,0,182,0);
signal scenario_full  : scenario_type := (0,0,113,31,1,31,215,31,85,31,84,31,35,31,46,31,46,30,238,31,12,31,40,31,40,30,109,31,161,31,161,30,152,31,152,30,193,31,137,31,22,31,22,30,22,29,28,31,64,31,227,31,117,31,199,31,47,31,235,31,219,31,20,31,45,31,166,31,166,30,166,29,106,31,193,31,9,31,172,31,103,31,250,31,255,31,52,31,52,30,19,31,186,31,23,31,221,31,221,30,161,31,252,31,188,31,188,30,196,31,196,30,196,29,8,31,247,31,16,31,168,31,170,31,155,31,20,31,135,31,147,31,17,31,17,30,190,31,251,31,137,31,119,31,128,31,128,30,128,29,173,31,205,31,205,30,206,31,145,31,99,31,99,30,131,31,11,31,74,31,219,31,44,31,229,31,231,31,198,31,166,31,166,30,166,29,119,31,79,31,228,31,228,30,59,31,30,31,158,31,114,31,165,31,1,31,50,31,48,31,164,31,83,31,89,31,58,31,58,30,148,31,148,30,120,31,120,30,206,31,235,31,220,31,220,30,220,29,70,31,148,31,148,30,148,29,190,31,58,31,245,31,237,31,237,30,33,31,126,31,160,31,160,30,235,31,10,31,114,31,114,30,160,31,6,31,87,31,78,31,226,31,115,31,111,31,39,31,51,31,61,31,61,30,38,31,204,31,23,31,135,31,132,31,205,31,58,31,138,31,138,30,55,31,244,31,73,31,134,31,157,31,175,31,154,31,154,30,33,31,98,31,247,31,247,30,145,31,160,31,71,31,68,31,120,31,55,31,55,30,212,31,69,31,127,31,106,31,106,30,106,29,253,31,253,30,242,31,51,31,56,31,163,31,94,31,86,31,9,31,4,31,219,31,177,31,160,31,160,30,174,31,174,30,181,31,164,31,131,31,131,30,90,31,42,31,101,31,133,31,214,31,214,30,115,31,60,31,107,31,107,30,141,31,161,31,251,31,63,31,63,30,219,31,219,30,219,29,135,31,135,30,119,31,232,31,100,31,8,31,50,31,31,31,208,31,78,31,78,30,205,31,8,31,88,31,88,30,123,31,39,31,229,31,243,31,31,31,20,31,20,30,203,31,46,31,151,31,49,31,188,31,88,31,9,31,9,31,113,31,156,31,233,31,105,31,105,30,208,31,217,31,45,31,113,31,50,31,11,31,250,31,199,31,91,31,201,31,242,31,235,31,235,30,8,31,231,31,249,31,249,30,249,29,249,28,249,27,119,31,119,30,211,31,211,30,189,31,10,31,92,31,174,31,174,30,60,31,117,31,253,31,150,31,132,31,16,31,72,31,69,31,69,30,89,31,43,31,43,30,114,31,94,31,16,31,26,31,160,31,162,31,122,31,65,31,143,31,248,31,191,31,17,31,166,31,8,31,8,30,8,29,172,31,114,31,114,30,211,31,209,31,209,30,4,31,4,30,51,31,28,31,114,31,222,31,250,31,9,31,123,31,229,31,130,31,81,31,90,31,118,31,67,31,67,30,250,31,135,31,22,31,104,31,98,31,76,31,40,31,184,31,184,30,98,31,121,31,106,31,106,30,3,31,119,31,114,31,114,30,5,31,231,31,121,31,138,31,125,31,6,31,6,30,107,31,224,31,18,31,18,30,102,31,102,30,94,31,163,31,251,31,28,31,233,31,143,31,86,31,135,31,246,31,220,31,197,31,36,31,36,30,211,31,153,31,153,30,129,31,112,31,112,30,208,31,208,30,188,31,46,31,23,31,23,30,68,31,68,30,68,29,172,31,159,31,159,30,159,29,159,28,251,31,251,30,192,31,12,31,246,31,182,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
