-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_940 is
end project_tb_940;

architecture project_tb_arch_940 of project_tb_940 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 487;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,222,0,0,0,0,0,182,0,18,0,0,0,1,0,162,0,249,0,108,0,137,0,0,0,0,0,0,0,156,0,102,0,213,0,50,0,0,0,191,0,20,0,96,0,213,0,155,0,17,0,0,0,97,0,161,0,9,0,20,0,0,0,19,0,159,0,0,0,249,0,81,0,119,0,247,0,241,0,31,0,37,0,0,0,231,0,201,0,0,0,25,0,135,0,228,0,84,0,221,0,0,0,5,0,163,0,104,0,148,0,142,0,79,0,219,0,18,0,0,0,229,0,82,0,0,0,91,0,0,0,0,0,0,0,0,0,17,0,0,0,23,0,57,0,0,0,0,0,38,0,193,0,1,0,0,0,173,0,192,0,142,0,0,0,65,0,104,0,176,0,63,0,202,0,215,0,66,0,6,0,115,0,211,0,215,0,247,0,48,0,0,0,225,0,39,0,204,0,88,0,0,0,167,0,191,0,0,0,0,0,158,0,170,0,0,0,70,0,127,0,122,0,216,0,0,0,8,0,73,0,0,0,85,0,178,0,51,0,85,0,149,0,113,0,0,0,93,0,0,0,167,0,230,0,0,0,0,0,248,0,207,0,180,0,96,0,132,0,38,0,71,0,112,0,148,0,115,0,211,0,13,0,166,0,25,0,207,0,211,0,62,0,33,0,158,0,98,0,144,0,72,0,151,0,254,0,209,0,234,0,114,0,215,0,175,0,0,0,238,0,61,0,203,0,240,0,159,0,195,0,198,0,212,0,220,0,235,0,149,0,45,0,0,0,0,0,0,0,248,0,0,0,0,0,235,0,0,0,131,0,90,0,18,0,0,0,107,0,125,0,27,0,186,0,118,0,37,0,0,0,0,0,221,0,10,0,55,0,0,0,228,0,225,0,171,0,123,0,105,0,38,0,249,0,173,0,54,0,193,0,85,0,125,0,47,0,146,0,160,0,150,0,28,0,235,0,18,0,250,0,217,0,0,0,101,0,109,0,41,0,79,0,5,0,41,0,128,0,169,0,12,0,13,0,92,0,0,0,43,0,0,0,170,0,0,0,0,0,37,0,38,0,247,0,236,0,77,0,78,0,0,0,2,0,0,0,75,0,0,0,158,0,187,0,82,0,37,0,19,0,32,0,0,0,28,0,0,0,0,0,159,0,54,0,0,0,199,0,105,0,247,0,205,0,228,0,0,0,45,0,182,0,75,0,0,0,39,0,49,0,0,0,0,0,209,0,42,0,236,0,254,0,93,0,43,0,226,0,197,0,0,0,135,0,239,0,173,0,137,0,154,0,0,0,198,0,40,0,67,0,233,0,67,0,52,0,185,0,114,0,132,0,180,0,146,0,0,0,59,0,151,0,180,0,70,0,0,0,103,0,110,0,189,0,186,0,12,0,74,0,0,0,40,0,43,0,215,0,207,0,94,0,236,0,207,0,219,0,236,0,161,0,31,0,82,0,86,0,0,0,215,0,203,0,31,0,0,0,231,0,0,0,35,0,153,0,111,0,241,0,102,0,0,0,0,0,150,0,0,0,102,0,141,0,177,0,0,0,77,0,193,0,112,0,168,0,14,0,2,0,104,0,127,0,0,0,248,0,119,0,216,0,15,0,147,0,218,0,24,0,0,0,253,0,0,0,213,0,207,0,205,0,81,0,109,0,182,0,0,0,0,0,115,0,17,0,233,0,91,0,0,0,132,0,0,0,113,0,244,0,176,0,100,0,147,0,42,0,166,0,145,0,7,0,253,0,241,0,0,0,50,0,144,0,143,0,94,0,68,0,232,0,0,0,0,0,110,0,31,0,0,0,0,0,252,0,206,0,149,0,125,0,15,0,58,0,13,0,186,0,0,0,57,0,222,0,103,0,223,0,0,0,48,0,0,0,175,0,215,0,0,0,176,0,101,0,252,0,231,0,160,0,0,0,33,0,92,0,0,0,152,0,110,0,32,0,57,0,26,0,120,0,252,0,201,0,0,0,173,0,214,0,111,0,0,0,55,0,82,0,148,0,133,0,8,0,53,0,0,0,179,0,237,0,215,0,98,0,227,0,169,0,0,0,71,0,186,0,0,0,37,0,0,0,0,0,38,0,100,0,240,0,135,0,153,0,3,0,12,0,12,0,0,0,48,0,232,0,6,0,0,0,175,0,246,0,92,0,17,0,103,0,19,0,159,0,99,0,92,0,207,0);
signal scenario_full  : scenario_type := (0,0,222,31,222,30,222,29,182,31,18,31,18,30,1,31,162,31,249,31,108,31,137,31,137,30,137,29,137,28,156,31,102,31,213,31,50,31,50,30,191,31,20,31,96,31,213,31,155,31,17,31,17,30,97,31,161,31,9,31,20,31,20,30,19,31,159,31,159,30,249,31,81,31,119,31,247,31,241,31,31,31,37,31,37,30,231,31,201,31,201,30,25,31,135,31,228,31,84,31,221,31,221,30,5,31,163,31,104,31,148,31,142,31,79,31,219,31,18,31,18,30,229,31,82,31,82,30,91,31,91,30,91,29,91,28,91,27,17,31,17,30,23,31,57,31,57,30,57,29,38,31,193,31,1,31,1,30,173,31,192,31,142,31,142,30,65,31,104,31,176,31,63,31,202,31,215,31,66,31,6,31,115,31,211,31,215,31,247,31,48,31,48,30,225,31,39,31,204,31,88,31,88,30,167,31,191,31,191,30,191,29,158,31,170,31,170,30,70,31,127,31,122,31,216,31,216,30,8,31,73,31,73,30,85,31,178,31,51,31,85,31,149,31,113,31,113,30,93,31,93,30,167,31,230,31,230,30,230,29,248,31,207,31,180,31,96,31,132,31,38,31,71,31,112,31,148,31,115,31,211,31,13,31,166,31,25,31,207,31,211,31,62,31,33,31,158,31,98,31,144,31,72,31,151,31,254,31,209,31,234,31,114,31,215,31,175,31,175,30,238,31,61,31,203,31,240,31,159,31,195,31,198,31,212,31,220,31,235,31,149,31,45,31,45,30,45,29,45,28,248,31,248,30,248,29,235,31,235,30,131,31,90,31,18,31,18,30,107,31,125,31,27,31,186,31,118,31,37,31,37,30,37,29,221,31,10,31,55,31,55,30,228,31,225,31,171,31,123,31,105,31,38,31,249,31,173,31,54,31,193,31,85,31,125,31,47,31,146,31,160,31,150,31,28,31,235,31,18,31,250,31,217,31,217,30,101,31,109,31,41,31,79,31,5,31,41,31,128,31,169,31,12,31,13,31,92,31,92,30,43,31,43,30,170,31,170,30,170,29,37,31,38,31,247,31,236,31,77,31,78,31,78,30,2,31,2,30,75,31,75,30,158,31,187,31,82,31,37,31,19,31,32,31,32,30,28,31,28,30,28,29,159,31,54,31,54,30,199,31,105,31,247,31,205,31,228,31,228,30,45,31,182,31,75,31,75,30,39,31,49,31,49,30,49,29,209,31,42,31,236,31,254,31,93,31,43,31,226,31,197,31,197,30,135,31,239,31,173,31,137,31,154,31,154,30,198,31,40,31,67,31,233,31,67,31,52,31,185,31,114,31,132,31,180,31,146,31,146,30,59,31,151,31,180,31,70,31,70,30,103,31,110,31,189,31,186,31,12,31,74,31,74,30,40,31,43,31,215,31,207,31,94,31,236,31,207,31,219,31,236,31,161,31,31,31,82,31,86,31,86,30,215,31,203,31,31,31,31,30,231,31,231,30,35,31,153,31,111,31,241,31,102,31,102,30,102,29,150,31,150,30,102,31,141,31,177,31,177,30,77,31,193,31,112,31,168,31,14,31,2,31,104,31,127,31,127,30,248,31,119,31,216,31,15,31,147,31,218,31,24,31,24,30,253,31,253,30,213,31,207,31,205,31,81,31,109,31,182,31,182,30,182,29,115,31,17,31,233,31,91,31,91,30,132,31,132,30,113,31,244,31,176,31,100,31,147,31,42,31,166,31,145,31,7,31,253,31,241,31,241,30,50,31,144,31,143,31,94,31,68,31,232,31,232,30,232,29,110,31,31,31,31,30,31,29,252,31,206,31,149,31,125,31,15,31,58,31,13,31,186,31,186,30,57,31,222,31,103,31,223,31,223,30,48,31,48,30,175,31,215,31,215,30,176,31,101,31,252,31,231,31,160,31,160,30,33,31,92,31,92,30,152,31,110,31,32,31,57,31,26,31,120,31,252,31,201,31,201,30,173,31,214,31,111,31,111,30,55,31,82,31,148,31,133,31,8,31,53,31,53,30,179,31,237,31,215,31,98,31,227,31,169,31,169,30,71,31,186,31,186,30,37,31,37,30,37,29,38,31,100,31,240,31,135,31,153,31,3,31,12,31,12,31,12,30,48,31,232,31,6,31,6,30,175,31,246,31,92,31,17,31,103,31,19,31,159,31,99,31,92,31,207,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
