-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 930;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (165,0,17,0,22,0,35,0,174,0,0,0,185,0,141,0,136,0,247,0,100,0,122,0,0,0,128,0,238,0,225,0,227,0,5,0,235,0,0,0,80,0,0,0,202,0,248,0,7,0,0,0,158,0,148,0,251,0,49,0,242,0,123,0,116,0,0,0,147,0,60,0,173,0,17,0,0,0,0,0,145,0,76,0,0,0,60,0,253,0,0,0,29,0,108,0,0,0,0,0,209,0,1,0,233,0,222,0,202,0,37,0,208,0,70,0,0,0,247,0,233,0,207,0,0,0,87,0,138,0,221,0,0,0,39,0,195,0,252,0,129,0,189,0,0,0,191,0,80,0,212,0,136,0,171,0,156,0,225,0,167,0,8,0,4,0,209,0,248,0,113,0,0,0,159,0,119,0,98,0,160,0,101,0,38,0,131,0,0,0,5,0,178,0,24,0,37,0,175,0,37,0,116,0,2,0,0,0,2,0,86,0,131,0,245,0,236,0,65,0,235,0,25,0,0,0,100,0,26,0,111,0,210,0,79,0,49,0,0,0,0,0,0,0,75,0,0,0,0,0,188,0,137,0,175,0,124,0,124,0,147,0,137,0,221,0,0,0,246,0,30,0,175,0,34,0,17,0,174,0,0,0,59,0,199,0,168,0,226,0,0,0,207,0,184,0,0,0,138,0,20,0,61,0,170,0,208,0,165,0,251,0,93,0,64,0,241,0,229,0,219,0,72,0,89,0,0,0,0,0,157,0,223,0,39,0,193,0,234,0,0,0,118,0,52,0,238,0,20,0,222,0,207,0,0,0,67,0,242,0,25,0,233,0,191,0,199,0,0,0,67,0,164,0,150,0,168,0,53,0,144,0,211,0,149,0,170,0,199,0,54,0,108,0,39,0,0,0,201,0,227,0,25,0,0,0,25,0,237,0,167,0,135,0,57,0,166,0,167,0,173,0,68,0,4,0,156,0,221,0,92,0,199,0,0,0,194,0,212,0,250,0,243,0,28,0,43,0,118,0,0,0,205,0,249,0,23,0,0,0,9,0,140,0,129,0,78,0,155,0,242,0,108,0,14,0,240,0,128,0,154,0,116,0,161,0,189,0,142,0,217,0,99,0,0,0,242,0,104,0,54,0,194,0,211,0,143,0,201,0,0,0,220,0,96,0,0,0,2,0,214,0,1,0,46,0,181,0,196,0,27,0,237,0,54,0,26,0,121,0,0,0,164,0,145,0,193,0,212,0,109,0,128,0,106,0,1,0,184,0,0,0,67,0,34,0,185,0,0,0,0,0,0,0,0,0,109,0,193,0,234,0,0,0,61,0,176,0,254,0,46,0,216,0,63,0,26,0,0,0,186,0,239,0,215,0,183,0,91,0,0,0,243,0,246,0,170,0,195,0,46,0,0,0,82,0,63,0,96,0,246,0,99,0,244,0,0,0,9,0,158,0,34,0,237,0,70,0,123,0,0,0,25,0,112,0,0,0,5,0,251,0,0,0,147,0,0,0,0,0,107,0,243,0,123,0,26,0,32,0,0,0,97,0,144,0,255,0,200,0,193,0,71,0,22,0,216,0,215,0,241,0,0,0,209,0,244,0,245,0,84,0,132,0,0,0,0,0,206,0,224,0,206,0,182,0,249,0,0,0,0,0,0,0,126,0,121,0,0,0,225,0,172,0,124,0,0,0,222,0,208,0,72,0,159,0,0,0,169,0,253,0,201,0,228,0,170,0,0,0,190,0,0,0,242,0,247,0,222,0,202,0,171,0,231,0,39,0,57,0,97,0,64,0,0,0,193,0,189,0,139,0,114,0,106,0,126,0,82,0,0,0,221,0,154,0,247,0,117,0,160,0,137,0,185,0,167,0,127,0,58,0,102,0,219,0,203,0,0,0,212,0,122,0,221,0,68,0,0,0,160,0,121,0,122,0,116,0,167,0,131,0,6,0,7,0,0,0,0,0,220,0,106,0,48,0,0,0,0,0,0,0,206,0,163,0,136,0,249,0,0,0,148,0,0,0,28,0,183,0,241,0,25,0,0,0,90,0,137,0,237,0,111,0,236,0,42,0,175,0,230,0,0,0,253,0,219,0,160,0,200,0,75,0,163,0,102,0,114,0,186,0,183,0,52,0,0,0,0,0,182,0,72,0,0,0,22,0,156,0,185,0,237,0,47,0,219,0,10,0,0,0,0,0,98,0,0,0,142,0,152,0,215,0,249,0,44,0,0,0,198,0,0,0,0,0,103,0,0,0,13,0,249,0,105,0,248,0,0,0,126,0,95,0,230,0,146,0,0,0,62,0,187,0,79,0,163,0,0,0,186,0,152,0,199,0,60,0,154,0,251,0,0,0,162,0,60,0,0,0,37,0,211,0,226,0,148,0,87,0,47,0,136,0,218,0,221,0,141,0,0,0,0,0,87,0,195,0,207,0,0,0,55,0,194,0,179,0,227,0,18,0,65,0,29,0,122,0,0,0,85,0,116,0,99,0,0,0,159,0,16,0,180,0,174,0,170,0,78,0,51,0,218,0,0,0,27,0,0,0,161,0,176,0,133,0,156,0,124,0,98,0,139,0,108,0,72,0,29,0,5,0,1,0,1,0,0,0,138,0,0,0,0,0,0,0,252,0,127,0,88,0,0,0,40,0,0,0,222,0,200,0,37,0,157,0,54,0,140,0,171,0,214,0,231,0,110,0,57,0,0,0,177,0,171,0,0,0,138,0,103,0,0,0,189,0,13,0,117,0,195,0,137,0,98,0,0,0,101,0,185,0,60,0,177,0,81,0,184,0,208,0,139,0,109,0,228,0,219,0,0,0,184,0,0,0,205,0,110,0,99,0,215,0,240,0,152,0,89,0,234,0,0,0,160,0,132,0,0,0,0,0,133,0,137,0,90,0,51,0,208,0,204,0,254,0,141,0,227,0,164,0,157,0,219,0,172,0,234,0,0,0,239,0,174,0,0,0,0,0,93,0,0,0,239,0,204,0,78,0,254,0,29,0,211,0,111,0,0,0,207,0,89,0,167,0,255,0,0,0,0,0,230,0,111,0,114,0,21,0,175,0,237,0,211,0,97,0,84,0,156,0,0,0,0,0,99,0,0,0,104,0,38,0,210,0,19,0,17,0,226,0,0,0,0,0,248,0,218,0,0,0,224,0,23,0,143,0,230,0,236,0,49,0,131,0,42,0,90,0,98,0,93,0,58,0,242,0,0,0,54,0,210,0,247,0,93,0,147,0,154,0,83,0,0,0,168,0,105,0,131,0,151,0,76,0,247,0,0,0,156,0,0,0,148,0,0,0,70,0,157,0,71,0,14,0,143,0,34,0,0,0,199,0,202,0,186,0,252,0,59,0,0,0,208,0,14,0,39,0,98,0,236,0,211,0,23,0,38,0,172,0,14,0,195,0,58,0,130,0,78,0,221,0,0,0,0,0,86,0,237,0,13,0,150,0,95,0,0,0,255,0,134,0,37,0,229,0,106,0,0,0,6,0,0,0,103,0,0,0,55,0,0,0,0,0,31,0,0,0,113,0,0,0,93,0,0,0,243,0,75,0,241,0,0,0,189,0,93,0,109,0,0,0,189,0,255,0,145,0,65,0,186,0,0,0,159,0,228,0,145,0,87,0,26,0,173,0,0,0,86,0,104,0,175,0,0,0,20,0,213,0,251,0,0,0,216,0,0,0,175,0,26,0,30,0,146,0,143,0,216,0,114,0,75,0,112,0,198,0,189,0,5,0,180,0,244,0,23,0,7,0,102,0,0,0,69,0,158,0,83,0,205,0,0,0,0,0,101,0,247,0,227,0,197,0,174,0,0,0,28,0,62,0,79,0,202,0,0,0,23,0,218,0,0,0,55,0,121,0,0,0,163,0,68,0,0,0,163,0,0,0,154,0,97,0,117,0,0,0,41,0,199,0,184,0,88,0,139,0,210,0,192,0,90,0,14,0,222,0,233,0,82,0,183,0,0,0,152,0,191,0,0,0,68,0,226,0,240,0,0,0,95,0,141,0,0,0,0,0,175,0,8,0,247,0,27,0,110,0,224,0,152,0,73,0,250,0,0,0,0,0,65,0,212,0,233,0,33,0,48,0,244,0,17,0,0,0,0,0,29,0,0,0,117,0,243,0,193,0,84,0,160,0,56,0,138,0,11,0,57,0,218,0,152,0,113,0,0,0);
signal scenario_full  : scenario_type := (165,31,17,31,22,31,35,31,174,31,174,30,185,31,141,31,136,31,247,31,100,31,122,31,122,30,128,31,238,31,225,31,227,31,5,31,235,31,235,30,80,31,80,30,202,31,248,31,7,31,7,30,158,31,148,31,251,31,49,31,242,31,123,31,116,31,116,30,147,31,60,31,173,31,17,31,17,30,17,29,145,31,76,31,76,30,60,31,253,31,253,30,29,31,108,31,108,30,108,29,209,31,1,31,233,31,222,31,202,31,37,31,208,31,70,31,70,30,247,31,233,31,207,31,207,30,87,31,138,31,221,31,221,30,39,31,195,31,252,31,129,31,189,31,189,30,191,31,80,31,212,31,136,31,171,31,156,31,225,31,167,31,8,31,4,31,209,31,248,31,113,31,113,30,159,31,119,31,98,31,160,31,101,31,38,31,131,31,131,30,5,31,178,31,24,31,37,31,175,31,37,31,116,31,2,31,2,30,2,31,86,31,131,31,245,31,236,31,65,31,235,31,25,31,25,30,100,31,26,31,111,31,210,31,79,31,49,31,49,30,49,29,49,28,75,31,75,30,75,29,188,31,137,31,175,31,124,31,124,31,147,31,137,31,221,31,221,30,246,31,30,31,175,31,34,31,17,31,174,31,174,30,59,31,199,31,168,31,226,31,226,30,207,31,184,31,184,30,138,31,20,31,61,31,170,31,208,31,165,31,251,31,93,31,64,31,241,31,229,31,219,31,72,31,89,31,89,30,89,29,157,31,223,31,39,31,193,31,234,31,234,30,118,31,52,31,238,31,20,31,222,31,207,31,207,30,67,31,242,31,25,31,233,31,191,31,199,31,199,30,67,31,164,31,150,31,168,31,53,31,144,31,211,31,149,31,170,31,199,31,54,31,108,31,39,31,39,30,201,31,227,31,25,31,25,30,25,31,237,31,167,31,135,31,57,31,166,31,167,31,173,31,68,31,4,31,156,31,221,31,92,31,199,31,199,30,194,31,212,31,250,31,243,31,28,31,43,31,118,31,118,30,205,31,249,31,23,31,23,30,9,31,140,31,129,31,78,31,155,31,242,31,108,31,14,31,240,31,128,31,154,31,116,31,161,31,189,31,142,31,217,31,99,31,99,30,242,31,104,31,54,31,194,31,211,31,143,31,201,31,201,30,220,31,96,31,96,30,2,31,214,31,1,31,46,31,181,31,196,31,27,31,237,31,54,31,26,31,121,31,121,30,164,31,145,31,193,31,212,31,109,31,128,31,106,31,1,31,184,31,184,30,67,31,34,31,185,31,185,30,185,29,185,28,185,27,109,31,193,31,234,31,234,30,61,31,176,31,254,31,46,31,216,31,63,31,26,31,26,30,186,31,239,31,215,31,183,31,91,31,91,30,243,31,246,31,170,31,195,31,46,31,46,30,82,31,63,31,96,31,246,31,99,31,244,31,244,30,9,31,158,31,34,31,237,31,70,31,123,31,123,30,25,31,112,31,112,30,5,31,251,31,251,30,147,31,147,30,147,29,107,31,243,31,123,31,26,31,32,31,32,30,97,31,144,31,255,31,200,31,193,31,71,31,22,31,216,31,215,31,241,31,241,30,209,31,244,31,245,31,84,31,132,31,132,30,132,29,206,31,224,31,206,31,182,31,249,31,249,30,249,29,249,28,126,31,121,31,121,30,225,31,172,31,124,31,124,30,222,31,208,31,72,31,159,31,159,30,169,31,253,31,201,31,228,31,170,31,170,30,190,31,190,30,242,31,247,31,222,31,202,31,171,31,231,31,39,31,57,31,97,31,64,31,64,30,193,31,189,31,139,31,114,31,106,31,126,31,82,31,82,30,221,31,154,31,247,31,117,31,160,31,137,31,185,31,167,31,127,31,58,31,102,31,219,31,203,31,203,30,212,31,122,31,221,31,68,31,68,30,160,31,121,31,122,31,116,31,167,31,131,31,6,31,7,31,7,30,7,29,220,31,106,31,48,31,48,30,48,29,48,28,206,31,163,31,136,31,249,31,249,30,148,31,148,30,28,31,183,31,241,31,25,31,25,30,90,31,137,31,237,31,111,31,236,31,42,31,175,31,230,31,230,30,253,31,219,31,160,31,200,31,75,31,163,31,102,31,114,31,186,31,183,31,52,31,52,30,52,29,182,31,72,31,72,30,22,31,156,31,185,31,237,31,47,31,219,31,10,31,10,30,10,29,98,31,98,30,142,31,152,31,215,31,249,31,44,31,44,30,198,31,198,30,198,29,103,31,103,30,13,31,249,31,105,31,248,31,248,30,126,31,95,31,230,31,146,31,146,30,62,31,187,31,79,31,163,31,163,30,186,31,152,31,199,31,60,31,154,31,251,31,251,30,162,31,60,31,60,30,37,31,211,31,226,31,148,31,87,31,47,31,136,31,218,31,221,31,141,31,141,30,141,29,87,31,195,31,207,31,207,30,55,31,194,31,179,31,227,31,18,31,65,31,29,31,122,31,122,30,85,31,116,31,99,31,99,30,159,31,16,31,180,31,174,31,170,31,78,31,51,31,218,31,218,30,27,31,27,30,161,31,176,31,133,31,156,31,124,31,98,31,139,31,108,31,72,31,29,31,5,31,1,31,1,31,1,30,138,31,138,30,138,29,138,28,252,31,127,31,88,31,88,30,40,31,40,30,222,31,200,31,37,31,157,31,54,31,140,31,171,31,214,31,231,31,110,31,57,31,57,30,177,31,171,31,171,30,138,31,103,31,103,30,189,31,13,31,117,31,195,31,137,31,98,31,98,30,101,31,185,31,60,31,177,31,81,31,184,31,208,31,139,31,109,31,228,31,219,31,219,30,184,31,184,30,205,31,110,31,99,31,215,31,240,31,152,31,89,31,234,31,234,30,160,31,132,31,132,30,132,29,133,31,137,31,90,31,51,31,208,31,204,31,254,31,141,31,227,31,164,31,157,31,219,31,172,31,234,31,234,30,239,31,174,31,174,30,174,29,93,31,93,30,239,31,204,31,78,31,254,31,29,31,211,31,111,31,111,30,207,31,89,31,167,31,255,31,255,30,255,29,230,31,111,31,114,31,21,31,175,31,237,31,211,31,97,31,84,31,156,31,156,30,156,29,99,31,99,30,104,31,38,31,210,31,19,31,17,31,226,31,226,30,226,29,248,31,218,31,218,30,224,31,23,31,143,31,230,31,236,31,49,31,131,31,42,31,90,31,98,31,93,31,58,31,242,31,242,30,54,31,210,31,247,31,93,31,147,31,154,31,83,31,83,30,168,31,105,31,131,31,151,31,76,31,247,31,247,30,156,31,156,30,148,31,148,30,70,31,157,31,71,31,14,31,143,31,34,31,34,30,199,31,202,31,186,31,252,31,59,31,59,30,208,31,14,31,39,31,98,31,236,31,211,31,23,31,38,31,172,31,14,31,195,31,58,31,130,31,78,31,221,31,221,30,221,29,86,31,237,31,13,31,150,31,95,31,95,30,255,31,134,31,37,31,229,31,106,31,106,30,6,31,6,30,103,31,103,30,55,31,55,30,55,29,31,31,31,30,113,31,113,30,93,31,93,30,243,31,75,31,241,31,241,30,189,31,93,31,109,31,109,30,189,31,255,31,145,31,65,31,186,31,186,30,159,31,228,31,145,31,87,31,26,31,173,31,173,30,86,31,104,31,175,31,175,30,20,31,213,31,251,31,251,30,216,31,216,30,175,31,26,31,30,31,146,31,143,31,216,31,114,31,75,31,112,31,198,31,189,31,5,31,180,31,244,31,23,31,7,31,102,31,102,30,69,31,158,31,83,31,205,31,205,30,205,29,101,31,247,31,227,31,197,31,174,31,174,30,28,31,62,31,79,31,202,31,202,30,23,31,218,31,218,30,55,31,121,31,121,30,163,31,68,31,68,30,163,31,163,30,154,31,97,31,117,31,117,30,41,31,199,31,184,31,88,31,139,31,210,31,192,31,90,31,14,31,222,31,233,31,82,31,183,31,183,30,152,31,191,31,191,30,68,31,226,31,240,31,240,30,95,31,141,31,141,30,141,29,175,31,8,31,247,31,27,31,110,31,224,31,152,31,73,31,250,31,250,30,250,29,65,31,212,31,233,31,33,31,48,31,244,31,17,31,17,30,17,29,29,31,29,30,117,31,243,31,193,31,84,31,160,31,56,31,138,31,11,31,57,31,218,31,152,31,113,31,113,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
