-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 856;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,40,0,249,0,162,0,0,0,27,0,218,0,0,0,0,0,206,0,0,0,0,0,89,0,71,0,0,0,206,0,101,0,0,0,0,0,60,0,173,0,103,0,108,0,117,0,214,0,0,0,102,0,142,0,13,0,32,0,87,0,0,0,0,0,197,0,174,0,98,0,80,0,139,0,0,0,0,0,199,0,158,0,106,0,222,0,182,0,21,0,0,0,0,0,118,0,58,0,169,0,253,0,201,0,131,0,19,0,102,0,14,0,166,0,0,0,56,0,218,0,67,0,0,0,0,0,120,0,0,0,236,0,0,0,92,0,74,0,242,0,0,0,157,0,57,0,0,0,0,0,99,0,170,0,149,0,135,0,21,0,199,0,97,0,0,0,217,0,251,0,140,0,108,0,136,0,91,0,78,0,162,0,0,0,9,0,109,0,210,0,0,0,18,0,241,0,0,0,69,0,21,0,36,0,111,0,212,0,50,0,0,0,79,0,142,0,0,0,156,0,112,0,92,0,102,0,166,0,0,0,41,0,0,0,224,0,20,0,0,0,195,0,181,0,35,0,240,0,0,0,135,0,179,0,3,0,0,0,80,0,0,0,0,0,114,0,238,0,135,0,163,0,245,0,0,0,170,0,89,0,41,0,20,0,149,0,203,0,0,0,6,0,207,0,221,0,97,0,133,0,33,0,161,0,131,0,0,0,225,0,121,0,74,0,102,0,190,0,216,0,226,0,160,0,227,0,7,0,0,0,109,0,6,0,148,0,0,0,192,0,182,0,170,0,164,0,157,0,236,0,86,0,179,0,170,0,173,0,217,0,88,0,51,0,25,0,201,0,43,0,225,0,246,0,21,0,27,0,0,0,105,0,177,0,29,0,90,0,218,0,0,0,19,0,100,0,214,0,163,0,0,0,0,0,189,0,20,0,0,0,213,0,27,0,42,0,139,0,244,0,43,0,0,0,165,0,72,0,0,0,255,0,20,0,133,0,145,0,157,0,146,0,0,0,211,0,155,0,39,0,179,0,0,0,148,0,122,0,96,0,198,0,15,0,106,0,181,0,95,0,0,0,200,0,226,0,0,0,228,0,149,0,215,0,118,0,39,0,167,0,0,0,11,0,113,0,154,0,63,0,0,0,161,0,9,0,70,0,232,0,0,0,203,0,38,0,129,0,0,0,129,0,0,0,24,0,8,0,17,0,82,0,73,0,212,0,27,0,0,0,124,0,17,0,34,0,0,0,205,0,0,0,71,0,229,0,146,0,72,0,208,0,205,0,220,0,238,0,249,0,188,0,14,0,109,0,250,0,0,0,0,0,197,0,51,0,145,0,2,0,0,0,0,0,16,0,210,0,91,0,0,0,204,0,213,0,97,0,175,0,0,0,0,0,123,0,16,0,0,0,53,0,174,0,0,0,0,0,221,0,3,0,237,0,166,0,53,0,75,0,20,0,243,0,28,0,32,0,213,0,80,0,69,0,99,0,195,0,241,0,178,0,55,0,37,0,121,0,208,0,203,0,0,0,98,0,0,0,231,0,0,0,71,0,247,0,0,0,206,0,46,0,0,0,0,0,55,0,130,0,132,0,91,0,0,0,73,0,0,0,89,0,0,0,107,0,0,0,62,0,247,0,221,0,67,0,70,0,105,0,0,0,133,0,104,0,141,0,106,0,246,0,134,0,150,0,121,0,229,0,0,0,127,0,6,0,56,0,15,0,69,0,21,0,131,0,0,0,160,0,66,0,206,0,0,0,11,0,145,0,198,0,101,0,0,0,0,0,224,0,141,0,43,0,215,0,0,0,57,0,0,0,121,0,233,0,24,0,165,0,126,0,83,0,238,0,64,0,0,0,141,0,15,0,8,0,95,0,182,0,0,0,71,0,0,0,46,0,109,0,43,0,0,0,250,0,229,0,0,0,70,0,28,0,166,0,56,0,32,0,104,0,183,0,164,0,152,0,0,0,8,0,61,0,0,0,0,0,0,0,36,0,177,0,17,0,159,0,8,0,65,0,0,0,0,0,119,0,142,0,0,0,6,0,37,0,245,0,226,0,58,0,66,0,0,0,145,0,15,0,63,0,206,0,0,0,51,0,51,0,126,0,238,0,195,0,94,0,143,0,0,0,56,0,217,0,16,0,217,0,121,0,41,0,61,0,0,0,23,0,228,0,203,0,52,0,168,0,70,0,192,0,77,0,99,0,229,0,0,0,0,0,137,0,89,0,61,0,21,0,115,0,168,0,0,0,0,0,20,0,231,0,183,0,2,0,64,0,34,0,212,0,197,0,77,0,202,0,201,0,0,0,135,0,120,0,91,0,191,0,123,0,0,0,86,0,0,0,197,0,14,0,84,0,0,0,81,0,0,0,0,0,109,0,0,0,207,0,174,0,200,0,0,0,97,0,78,0,210,0,0,0,252,0,170,0,119,0,118,0,0,0,168,0,130,0,104,0,101,0,13,0,36,0,151,0,212,0,0,0,140,0,199,0,224,0,161,0,0,0,139,0,69,0,0,0,0,0,0,0,240,0,5,0,227,0,0,0,173,0,0,0,228,0,178,0,0,0,133,0,0,0,58,0,29,0,130,0,178,0,15,0,0,0,18,0,97,0,96,0,14,0,212,0,67,0,50,0,116,0,127,0,171,0,57,0,0,0,122,0,111,0,56,0,184,0,0,0,0,0,0,0,251,0,142,0,16,0,140,0,0,0,243,0,106,0,37,0,0,0,241,0,11,0,60,0,0,0,122,0,66,0,27,0,244,0,0,0,7,0,46,0,184,0,0,0,126,0,51,0,152,0,0,0,41,0,218,0,0,0,154,0,0,0,142,0,37,0,58,0,238,0,0,0,82,0,7,0,136,0,0,0,97,0,188,0,212,0,0,0,51,0,26,0,228,0,163,0,46,0,97,0,39,0,123,0,83,0,121,0,244,0,69,0,235,0,156,0,42,0,134,0,172,0,227,0,204,0,224,0,138,0,75,0,130,0,164,0,0,0,197,0,3,0,0,0,26,0,166,0,158,0,0,0,253,0,11,0,0,0,193,0,0,0,0,0,25,0,82,0,91,0,193,0,0,0,145,0,80,0,0,0,38,0,71,0,47,0,159,0,90,0,203,0,139,0,114,0,82,0,216,0,35,0,87,0,44,0,92,0,26,0,0,0,0,0,194,0,0,0,0,0,78,0,0,0,50,0,39,0,107,0,67,0,247,0,201,0,55,0,0,0,92,0,109,0,119,0,54,0,253,0,243,0,0,0,207,0,89,0,0,0,41,0,169,0,33,0,10,0,82,0,63,0,100,0,77,0,43,0,0,0,86,0,0,0,63,0,165,0,190,0,7,0,60,0,209,0,0,0,253,0,194,0,227,0,0,0,123,0,95,0,0,0,255,0,2,0,232,0,172,0,248,0,161,0,0,0,0,0,245,0,178,0,216,0,245,0,0,0,238,0,228,0,38,0,91,0,241,0,4,0,179,0,85,0,64,0,252,0,246,0,0,0,206,0,194,0,232,0,0,0,0,0,129,0,147,0,129,0,194,0,213,0,0,0,29,0,0,0,45,0,92,0,238,0,239,0,1,0,218,0,143,0,15,0,227,0,13,0,127,0,157,0,0,0,142,0,41,0,210,0,223,0,205,0,42,0,10,0,20,0,0,0,236,0,50,0,0,0,144,0,167,0,0,0,209,0,102,0,0,0,234,0,183,0,198,0,32,0,10,0,0,0,152,0,7,0,197,0,217,0,101,0,0,0,218,0,149,0,0,0,195,0,48,0,84,0,242,0,239,0,122,0,251,0,139,0,16,0,196,0,70,0,0,0,39,0,0,0,216,0,239,0,0,0,104,0,254,0);
signal scenario_full  : scenario_type := (0,0,40,31,249,31,162,31,162,30,27,31,218,31,218,30,218,29,206,31,206,30,206,29,89,31,71,31,71,30,206,31,101,31,101,30,101,29,60,31,173,31,103,31,108,31,117,31,214,31,214,30,102,31,142,31,13,31,32,31,87,31,87,30,87,29,197,31,174,31,98,31,80,31,139,31,139,30,139,29,199,31,158,31,106,31,222,31,182,31,21,31,21,30,21,29,118,31,58,31,169,31,253,31,201,31,131,31,19,31,102,31,14,31,166,31,166,30,56,31,218,31,67,31,67,30,67,29,120,31,120,30,236,31,236,30,92,31,74,31,242,31,242,30,157,31,57,31,57,30,57,29,99,31,170,31,149,31,135,31,21,31,199,31,97,31,97,30,217,31,251,31,140,31,108,31,136,31,91,31,78,31,162,31,162,30,9,31,109,31,210,31,210,30,18,31,241,31,241,30,69,31,21,31,36,31,111,31,212,31,50,31,50,30,79,31,142,31,142,30,156,31,112,31,92,31,102,31,166,31,166,30,41,31,41,30,224,31,20,31,20,30,195,31,181,31,35,31,240,31,240,30,135,31,179,31,3,31,3,30,80,31,80,30,80,29,114,31,238,31,135,31,163,31,245,31,245,30,170,31,89,31,41,31,20,31,149,31,203,31,203,30,6,31,207,31,221,31,97,31,133,31,33,31,161,31,131,31,131,30,225,31,121,31,74,31,102,31,190,31,216,31,226,31,160,31,227,31,7,31,7,30,109,31,6,31,148,31,148,30,192,31,182,31,170,31,164,31,157,31,236,31,86,31,179,31,170,31,173,31,217,31,88,31,51,31,25,31,201,31,43,31,225,31,246,31,21,31,27,31,27,30,105,31,177,31,29,31,90,31,218,31,218,30,19,31,100,31,214,31,163,31,163,30,163,29,189,31,20,31,20,30,213,31,27,31,42,31,139,31,244,31,43,31,43,30,165,31,72,31,72,30,255,31,20,31,133,31,145,31,157,31,146,31,146,30,211,31,155,31,39,31,179,31,179,30,148,31,122,31,96,31,198,31,15,31,106,31,181,31,95,31,95,30,200,31,226,31,226,30,228,31,149,31,215,31,118,31,39,31,167,31,167,30,11,31,113,31,154,31,63,31,63,30,161,31,9,31,70,31,232,31,232,30,203,31,38,31,129,31,129,30,129,31,129,30,24,31,8,31,17,31,82,31,73,31,212,31,27,31,27,30,124,31,17,31,34,31,34,30,205,31,205,30,71,31,229,31,146,31,72,31,208,31,205,31,220,31,238,31,249,31,188,31,14,31,109,31,250,31,250,30,250,29,197,31,51,31,145,31,2,31,2,30,2,29,16,31,210,31,91,31,91,30,204,31,213,31,97,31,175,31,175,30,175,29,123,31,16,31,16,30,53,31,174,31,174,30,174,29,221,31,3,31,237,31,166,31,53,31,75,31,20,31,243,31,28,31,32,31,213,31,80,31,69,31,99,31,195,31,241,31,178,31,55,31,37,31,121,31,208,31,203,31,203,30,98,31,98,30,231,31,231,30,71,31,247,31,247,30,206,31,46,31,46,30,46,29,55,31,130,31,132,31,91,31,91,30,73,31,73,30,89,31,89,30,107,31,107,30,62,31,247,31,221,31,67,31,70,31,105,31,105,30,133,31,104,31,141,31,106,31,246,31,134,31,150,31,121,31,229,31,229,30,127,31,6,31,56,31,15,31,69,31,21,31,131,31,131,30,160,31,66,31,206,31,206,30,11,31,145,31,198,31,101,31,101,30,101,29,224,31,141,31,43,31,215,31,215,30,57,31,57,30,121,31,233,31,24,31,165,31,126,31,83,31,238,31,64,31,64,30,141,31,15,31,8,31,95,31,182,31,182,30,71,31,71,30,46,31,109,31,43,31,43,30,250,31,229,31,229,30,70,31,28,31,166,31,56,31,32,31,104,31,183,31,164,31,152,31,152,30,8,31,61,31,61,30,61,29,61,28,36,31,177,31,17,31,159,31,8,31,65,31,65,30,65,29,119,31,142,31,142,30,6,31,37,31,245,31,226,31,58,31,66,31,66,30,145,31,15,31,63,31,206,31,206,30,51,31,51,31,126,31,238,31,195,31,94,31,143,31,143,30,56,31,217,31,16,31,217,31,121,31,41,31,61,31,61,30,23,31,228,31,203,31,52,31,168,31,70,31,192,31,77,31,99,31,229,31,229,30,229,29,137,31,89,31,61,31,21,31,115,31,168,31,168,30,168,29,20,31,231,31,183,31,2,31,64,31,34,31,212,31,197,31,77,31,202,31,201,31,201,30,135,31,120,31,91,31,191,31,123,31,123,30,86,31,86,30,197,31,14,31,84,31,84,30,81,31,81,30,81,29,109,31,109,30,207,31,174,31,200,31,200,30,97,31,78,31,210,31,210,30,252,31,170,31,119,31,118,31,118,30,168,31,130,31,104,31,101,31,13,31,36,31,151,31,212,31,212,30,140,31,199,31,224,31,161,31,161,30,139,31,69,31,69,30,69,29,69,28,240,31,5,31,227,31,227,30,173,31,173,30,228,31,178,31,178,30,133,31,133,30,58,31,29,31,130,31,178,31,15,31,15,30,18,31,97,31,96,31,14,31,212,31,67,31,50,31,116,31,127,31,171,31,57,31,57,30,122,31,111,31,56,31,184,31,184,30,184,29,184,28,251,31,142,31,16,31,140,31,140,30,243,31,106,31,37,31,37,30,241,31,11,31,60,31,60,30,122,31,66,31,27,31,244,31,244,30,7,31,46,31,184,31,184,30,126,31,51,31,152,31,152,30,41,31,218,31,218,30,154,31,154,30,142,31,37,31,58,31,238,31,238,30,82,31,7,31,136,31,136,30,97,31,188,31,212,31,212,30,51,31,26,31,228,31,163,31,46,31,97,31,39,31,123,31,83,31,121,31,244,31,69,31,235,31,156,31,42,31,134,31,172,31,227,31,204,31,224,31,138,31,75,31,130,31,164,31,164,30,197,31,3,31,3,30,26,31,166,31,158,31,158,30,253,31,11,31,11,30,193,31,193,30,193,29,25,31,82,31,91,31,193,31,193,30,145,31,80,31,80,30,38,31,71,31,47,31,159,31,90,31,203,31,139,31,114,31,82,31,216,31,35,31,87,31,44,31,92,31,26,31,26,30,26,29,194,31,194,30,194,29,78,31,78,30,50,31,39,31,107,31,67,31,247,31,201,31,55,31,55,30,92,31,109,31,119,31,54,31,253,31,243,31,243,30,207,31,89,31,89,30,41,31,169,31,33,31,10,31,82,31,63,31,100,31,77,31,43,31,43,30,86,31,86,30,63,31,165,31,190,31,7,31,60,31,209,31,209,30,253,31,194,31,227,31,227,30,123,31,95,31,95,30,255,31,2,31,232,31,172,31,248,31,161,31,161,30,161,29,245,31,178,31,216,31,245,31,245,30,238,31,228,31,38,31,91,31,241,31,4,31,179,31,85,31,64,31,252,31,246,31,246,30,206,31,194,31,232,31,232,30,232,29,129,31,147,31,129,31,194,31,213,31,213,30,29,31,29,30,45,31,92,31,238,31,239,31,1,31,218,31,143,31,15,31,227,31,13,31,127,31,157,31,157,30,142,31,41,31,210,31,223,31,205,31,42,31,10,31,20,31,20,30,236,31,50,31,50,30,144,31,167,31,167,30,209,31,102,31,102,30,234,31,183,31,198,31,32,31,10,31,10,30,152,31,7,31,197,31,217,31,101,31,101,30,218,31,149,31,149,30,195,31,48,31,84,31,242,31,239,31,122,31,251,31,139,31,16,31,196,31,70,31,70,30,39,31,39,30,216,31,239,31,239,30,104,31,254,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
