-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_506 is
end project_tb_506;

architecture project_tb_arch_506 of project_tb_506 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 734;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (17,0,28,0,165,0,11,0,17,0,50,0,120,0,14,0,88,0,165,0,146,0,0,0,167,0,54,0,195,0,43,0,116,0,206,0,72,0,42,0,3,0,0,0,43,0,168,0,221,0,238,0,74,0,1,0,0,0,91,0,189,0,167,0,199,0,0,0,0,0,209,0,23,0,71,0,234,0,57,0,0,0,117,0,178,0,164,0,246,0,0,0,49,0,75,0,139,0,0,0,44,0,111,0,243,0,57,0,111,0,196,0,0,0,23,0,25,0,92,0,238,0,244,0,120,0,60,0,37,0,0,0,120,0,0,0,249,0,126,0,14,0,0,0,171,0,205,0,0,0,18,0,70,0,0,0,175,0,207,0,0,0,125,0,155,0,214,0,7,0,41,0,191,0,196,0,0,0,62,0,121,0,0,0,2,0,186,0,40,0,0,0,12,0,23,0,0,0,143,0,0,0,101,0,128,0,203,0,106,0,0,0,40,0,0,0,188,0,178,0,41,0,100,0,57,0,0,0,89,0,0,0,186,0,225,0,160,0,233,0,30,0,81,0,222,0,218,0,0,0,0,0,0,0,0,0,0,0,81,0,0,0,81,0,74,0,206,0,33,0,80,0,0,0,134,0,80,0,88,0,61,0,103,0,204,0,0,0,111,0,21,0,0,0,249,0,117,0,2,0,222,0,65,0,99,0,14,0,213,0,229,0,121,0,222,0,65,0,0,0,102,0,101,0,47,0,63,0,7,0,204,0,151,0,32,0,222,0,138,0,59,0,231,0,139,0,246,0,134,0,177,0,230,0,162,0,0,0,126,0,0,0,55,0,201,0,186,0,32,0,18,0,177,0,38,0,3,0,84,0,0,0,250,0,0,0,197,0,15,0,89,0,143,0,0,0,205,0,143,0,0,0,0,0,44,0,223,0,186,0,243,0,0,0,46,0,17,0,55,0,172,0,0,0,0,0,0,0,0,0,0,0,123,0,0,0,215,0,3,0,102,0,0,0,247,0,0,0,175,0,0,0,107,0,88,0,0,0,243,0,116,0,129,0,104,0,245,0,35,0,55,0,0,0,0,0,49,0,35,0,29,0,46,0,218,0,242,0,205,0,59,0,0,0,64,0,76,0,47,0,44,0,92,0,249,0,237,0,19,0,2,0,102,0,67,0,0,0,157,0,0,0,192,0,160,0,160,0,27,0,0,0,30,0,240,0,107,0,133,0,83,0,36,0,204,0,215,0,93,0,12,0,203,0,13,0,33,0,110,0,235,0,194,0,78,0,0,0,168,0,244,0,148,0,155,0,185,0,171,0,133,0,208,0,191,0,225,0,207,0,167,0,248,0,159,0,0,0,243,0,81,0,0,0,98,0,0,0,73,0,66,0,0,0,0,0,190,0,174,0,212,0,0,0,136,0,95,0,224,0,0,0,252,0,69,0,101,0,149,0,152,0,186,0,100,0,54,0,0,0,150,0,121,0,74,0,0,0,137,0,21,0,0,0,149,0,220,0,184,0,142,0,182,0,136,0,162,0,180,0,13,0,180,0,249,0,86,0,13,0,63,0,59,0,51,0,35,0,184,0,186,0,0,0,86,0,170,0,252,0,205,0,82,0,45,0,40,0,9,0,50,0,164,0,208,0,0,0,58,0,53,0,35,0,41,0,78,0,0,0,63,0,236,0,109,0,184,0,89,0,160,0,0,0,78,0,104,0,255,0,151,0,97,0,237,0,214,0,211,0,40,0,175,0,153,0,113,0,8,0,29,0,82,0,120,0,244,0,0,0,112,0,152,0,105,0,15,0,0,0,0,0,0,0,129,0,18,0,112,0,96,0,130,0,66,0,187,0,97,0,227,0,243,0,164,0,115,0,101,0,161,0,155,0,59,0,0,0,0,0,27,0,0,0,0,0,172,0,4,0,18,0,0,0,225,0,29,0,221,0,174,0,143,0,3,0,0,0,198,0,0,0,243,0,235,0,243,0,78,0,79,0,147,0,8,0,51,0,71,0,0,0,45,0,14,0,0,0,197,0,71,0,226,0,214,0,129,0,0,0,151,0,201,0,149,0,31,0,127,0,205,0,138,0,239,0,200,0,191,0,17,0,217,0,12,0,112,0,64,0,60,0,193,0,13,0,72,0,0,0,205,0,55,0,0,0,147,0,6,0,21,0,215,0,218,0,78,0,77,0,4,0,193,0,124,0,91,0,0,0,133,0,45,0,105,0,0,0,224,0,128,0,40,0,247,0,194,0,0,0,35,0,192,0,6,0,0,0,81,0,181,0,0,0,37,0,0,0,250,0,0,0,0,0,0,0,253,0,1,0,56,0,211,0,245,0,186,0,2,0,207,0,209,0,0,0,116,0,133,0,29,0,76,0,86,0,128,0,0,0,132,0,238,0,197,0,254,0,0,0,9,0,0,0,54,0,248,0,0,0,0,0,129,0,0,0,103,0,86,0,76,0,19,0,58,0,180,0,144,0,105,0,239,0,76,0,105,0,243,0,0,0,87,0,243,0,244,0,122,0,246,0,0,0,250,0,0,0,0,0,215,0,0,0,210,0,0,0,71,0,165,0,0,0,1,0,0,0,239,0,0,0,107,0,0,0,43,0,83,0,43,0,180,0,68,0,4,0,94,0,0,0,71,0,215,0,0,0,59,0,0,0,0,0,0,0,146,0,213,0,214,0,251,0,55,0,194,0,0,0,1,0,149,0,190,0,78,0,206,0,205,0,58,0,44,0,177,0,63,0,17,0,232,0,148,0,238,0,106,0,193,0,0,0,247,0,199,0,200,0,0,0,38,0,46,0,7,0,52,0,172,0,29,0,223,0,174,0,0,0,28,0,175,0,0,0,4,0,43,0,166,0,59,0,0,0,150,0,200,0,0,0,83,0,206,0,0,0,230,0,0,0,125,0,208,0,150,0,129,0,22,0,0,0,235,0,59,0,65,0,109,0,32,0,0,0,8,0,182,0,225,0,205,0,215,0,96,0,61,0,90,0,153,0,102,0,25,0,0,0,0,0,86,0,173,0,95,0,176,0,152,0,151,0,0,0,49,0,46,0,18,0,219,0,125,0,179,0,118,0,0,0,173,0,77,0,154,0,103,0,197,0,33,0,44,0,70,0,17,0,60,0,0,0,26,0,73,0,0,0,48,0,73,0,164,0,69,0,38,0,201,0,68,0,0,0,35,0,41,0,56,0,0,0,230,0,90,0,54,0,0,0,142,0,0,0,0,0,28,0,2,0,246,0,120,0,188,0,166,0,0,0,183,0,46,0,123,0,204,0,98,0,212,0,198,0,221,0);
signal scenario_full  : scenario_type := (17,31,28,31,165,31,11,31,17,31,50,31,120,31,14,31,88,31,165,31,146,31,146,30,167,31,54,31,195,31,43,31,116,31,206,31,72,31,42,31,3,31,3,30,43,31,168,31,221,31,238,31,74,31,1,31,1,30,91,31,189,31,167,31,199,31,199,30,199,29,209,31,23,31,71,31,234,31,57,31,57,30,117,31,178,31,164,31,246,31,246,30,49,31,75,31,139,31,139,30,44,31,111,31,243,31,57,31,111,31,196,31,196,30,23,31,25,31,92,31,238,31,244,31,120,31,60,31,37,31,37,30,120,31,120,30,249,31,126,31,14,31,14,30,171,31,205,31,205,30,18,31,70,31,70,30,175,31,207,31,207,30,125,31,155,31,214,31,7,31,41,31,191,31,196,31,196,30,62,31,121,31,121,30,2,31,186,31,40,31,40,30,12,31,23,31,23,30,143,31,143,30,101,31,128,31,203,31,106,31,106,30,40,31,40,30,188,31,178,31,41,31,100,31,57,31,57,30,89,31,89,30,186,31,225,31,160,31,233,31,30,31,81,31,222,31,218,31,218,30,218,29,218,28,218,27,218,26,81,31,81,30,81,31,74,31,206,31,33,31,80,31,80,30,134,31,80,31,88,31,61,31,103,31,204,31,204,30,111,31,21,31,21,30,249,31,117,31,2,31,222,31,65,31,99,31,14,31,213,31,229,31,121,31,222,31,65,31,65,30,102,31,101,31,47,31,63,31,7,31,204,31,151,31,32,31,222,31,138,31,59,31,231,31,139,31,246,31,134,31,177,31,230,31,162,31,162,30,126,31,126,30,55,31,201,31,186,31,32,31,18,31,177,31,38,31,3,31,84,31,84,30,250,31,250,30,197,31,15,31,89,31,143,31,143,30,205,31,143,31,143,30,143,29,44,31,223,31,186,31,243,31,243,30,46,31,17,31,55,31,172,31,172,30,172,29,172,28,172,27,172,26,123,31,123,30,215,31,3,31,102,31,102,30,247,31,247,30,175,31,175,30,107,31,88,31,88,30,243,31,116,31,129,31,104,31,245,31,35,31,55,31,55,30,55,29,49,31,35,31,29,31,46,31,218,31,242,31,205,31,59,31,59,30,64,31,76,31,47,31,44,31,92,31,249,31,237,31,19,31,2,31,102,31,67,31,67,30,157,31,157,30,192,31,160,31,160,31,27,31,27,30,30,31,240,31,107,31,133,31,83,31,36,31,204,31,215,31,93,31,12,31,203,31,13,31,33,31,110,31,235,31,194,31,78,31,78,30,168,31,244,31,148,31,155,31,185,31,171,31,133,31,208,31,191,31,225,31,207,31,167,31,248,31,159,31,159,30,243,31,81,31,81,30,98,31,98,30,73,31,66,31,66,30,66,29,190,31,174,31,212,31,212,30,136,31,95,31,224,31,224,30,252,31,69,31,101,31,149,31,152,31,186,31,100,31,54,31,54,30,150,31,121,31,74,31,74,30,137,31,21,31,21,30,149,31,220,31,184,31,142,31,182,31,136,31,162,31,180,31,13,31,180,31,249,31,86,31,13,31,63,31,59,31,51,31,35,31,184,31,186,31,186,30,86,31,170,31,252,31,205,31,82,31,45,31,40,31,9,31,50,31,164,31,208,31,208,30,58,31,53,31,35,31,41,31,78,31,78,30,63,31,236,31,109,31,184,31,89,31,160,31,160,30,78,31,104,31,255,31,151,31,97,31,237,31,214,31,211,31,40,31,175,31,153,31,113,31,8,31,29,31,82,31,120,31,244,31,244,30,112,31,152,31,105,31,15,31,15,30,15,29,15,28,129,31,18,31,112,31,96,31,130,31,66,31,187,31,97,31,227,31,243,31,164,31,115,31,101,31,161,31,155,31,59,31,59,30,59,29,27,31,27,30,27,29,172,31,4,31,18,31,18,30,225,31,29,31,221,31,174,31,143,31,3,31,3,30,198,31,198,30,243,31,235,31,243,31,78,31,79,31,147,31,8,31,51,31,71,31,71,30,45,31,14,31,14,30,197,31,71,31,226,31,214,31,129,31,129,30,151,31,201,31,149,31,31,31,127,31,205,31,138,31,239,31,200,31,191,31,17,31,217,31,12,31,112,31,64,31,60,31,193,31,13,31,72,31,72,30,205,31,55,31,55,30,147,31,6,31,21,31,215,31,218,31,78,31,77,31,4,31,193,31,124,31,91,31,91,30,133,31,45,31,105,31,105,30,224,31,128,31,40,31,247,31,194,31,194,30,35,31,192,31,6,31,6,30,81,31,181,31,181,30,37,31,37,30,250,31,250,30,250,29,250,28,253,31,1,31,56,31,211,31,245,31,186,31,2,31,207,31,209,31,209,30,116,31,133,31,29,31,76,31,86,31,128,31,128,30,132,31,238,31,197,31,254,31,254,30,9,31,9,30,54,31,248,31,248,30,248,29,129,31,129,30,103,31,86,31,76,31,19,31,58,31,180,31,144,31,105,31,239,31,76,31,105,31,243,31,243,30,87,31,243,31,244,31,122,31,246,31,246,30,250,31,250,30,250,29,215,31,215,30,210,31,210,30,71,31,165,31,165,30,1,31,1,30,239,31,239,30,107,31,107,30,43,31,83,31,43,31,180,31,68,31,4,31,94,31,94,30,71,31,215,31,215,30,59,31,59,30,59,29,59,28,146,31,213,31,214,31,251,31,55,31,194,31,194,30,1,31,149,31,190,31,78,31,206,31,205,31,58,31,44,31,177,31,63,31,17,31,232,31,148,31,238,31,106,31,193,31,193,30,247,31,199,31,200,31,200,30,38,31,46,31,7,31,52,31,172,31,29,31,223,31,174,31,174,30,28,31,175,31,175,30,4,31,43,31,166,31,59,31,59,30,150,31,200,31,200,30,83,31,206,31,206,30,230,31,230,30,125,31,208,31,150,31,129,31,22,31,22,30,235,31,59,31,65,31,109,31,32,31,32,30,8,31,182,31,225,31,205,31,215,31,96,31,61,31,90,31,153,31,102,31,25,31,25,30,25,29,86,31,173,31,95,31,176,31,152,31,151,31,151,30,49,31,46,31,18,31,219,31,125,31,179,31,118,31,118,30,173,31,77,31,154,31,103,31,197,31,33,31,44,31,70,31,17,31,60,31,60,30,26,31,73,31,73,30,48,31,73,31,164,31,69,31,38,31,201,31,68,31,68,30,35,31,41,31,56,31,56,30,230,31,90,31,54,31,54,30,142,31,142,30,142,29,28,31,2,31,246,31,120,31,188,31,166,31,166,30,183,31,46,31,123,31,204,31,98,31,212,31,198,31,221,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
