-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_906 is
end project_tb_906;

architecture project_tb_arch_906 of project_tb_906 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 228;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (63,0,146,0,193,0,0,0,184,0,60,0,33,0,241,0,67,0,81,0,0,0,203,0,220,0,0,0,11,0,241,0,106,0,87,0,225,0,0,0,160,0,96,0,216,0,41,0,164,0,0,0,194,0,103,0,3,0,48,0,156,0,0,0,213,0,244,0,251,0,61,0,217,0,124,0,0,0,52,0,114,0,0,0,222,0,112,0,237,0,143,0,148,0,0,0,0,0,236,0,117,0,197,0,209,0,0,0,125,0,0,0,187,0,215,0,158,0,0,0,38,0,24,0,0,0,146,0,142,0,125,0,98,0,22,0,175,0,0,0,87,0,240,0,26,0,97,0,255,0,94,0,248,0,228,0,33,0,0,0,0,0,0,0,132,0,56,0,163,0,0,0,213,0,20,0,82,0,84,0,230,0,78,0,214,0,56,0,0,0,29,0,217,0,75,0,0,0,11,0,52,0,222,0,238,0,136,0,16,0,176,0,154,0,59,0,254,0,167,0,0,0,34,0,124,0,216,0,0,0,149,0,58,0,115,0,0,0,227,0,197,0,0,0,0,0,37,0,0,0,89,0,160,0,113,0,139,0,147,0,51,0,164,0,192,0,56,0,74,0,0,0,0,0,0,0,44,0,213,0,136,0,61,0,120,0,9,0,180,0,168,0,72,0,254,0,70,0,96,0,204,0,0,0,173,0,235,0,60,0,0,0,0,0,0,0,0,0,31,0,0,0,244,0,0,0,92,0,207,0,111,0,168,0,0,0,122,0,205,0,93,0,0,0,66,0,67,0,0,0,185,0,24,0,22,0,0,0,223,0,204,0,0,0,16,0,52,0,78,0,9,0,53,0,81,0,1,0,146,0,44,0,0,0,40,0,144,0,146,0,61,0,37,0,56,0,161,0,121,0,207,0,161,0,177,0,0,0,159,0,0,0,94,0,249,0,35,0,59,0,0,0,15,0,14,0,0,0,0,0,156,0,59,0,80,0,17,0,0,0,0,0,29,0,69,0,40,0,0,0,105,0,99,0,104,0);
signal scenario_full  : scenario_type := (63,31,146,31,193,31,193,30,184,31,60,31,33,31,241,31,67,31,81,31,81,30,203,31,220,31,220,30,11,31,241,31,106,31,87,31,225,31,225,30,160,31,96,31,216,31,41,31,164,31,164,30,194,31,103,31,3,31,48,31,156,31,156,30,213,31,244,31,251,31,61,31,217,31,124,31,124,30,52,31,114,31,114,30,222,31,112,31,237,31,143,31,148,31,148,30,148,29,236,31,117,31,197,31,209,31,209,30,125,31,125,30,187,31,215,31,158,31,158,30,38,31,24,31,24,30,146,31,142,31,125,31,98,31,22,31,175,31,175,30,87,31,240,31,26,31,97,31,255,31,94,31,248,31,228,31,33,31,33,30,33,29,33,28,132,31,56,31,163,31,163,30,213,31,20,31,82,31,84,31,230,31,78,31,214,31,56,31,56,30,29,31,217,31,75,31,75,30,11,31,52,31,222,31,238,31,136,31,16,31,176,31,154,31,59,31,254,31,167,31,167,30,34,31,124,31,216,31,216,30,149,31,58,31,115,31,115,30,227,31,197,31,197,30,197,29,37,31,37,30,89,31,160,31,113,31,139,31,147,31,51,31,164,31,192,31,56,31,74,31,74,30,74,29,74,28,44,31,213,31,136,31,61,31,120,31,9,31,180,31,168,31,72,31,254,31,70,31,96,31,204,31,204,30,173,31,235,31,60,31,60,30,60,29,60,28,60,27,31,31,31,30,244,31,244,30,92,31,207,31,111,31,168,31,168,30,122,31,205,31,93,31,93,30,66,31,67,31,67,30,185,31,24,31,22,31,22,30,223,31,204,31,204,30,16,31,52,31,78,31,9,31,53,31,81,31,1,31,146,31,44,31,44,30,40,31,144,31,146,31,61,31,37,31,56,31,161,31,121,31,207,31,161,31,177,31,177,30,159,31,159,30,94,31,249,31,35,31,59,31,59,30,15,31,14,31,14,30,14,29,156,31,59,31,80,31,17,31,17,30,17,29,29,31,69,31,40,31,40,30,105,31,99,31,104,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
