-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_362 is
end project_tb_362;

architecture project_tb_arch_362 of project_tb_362 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 639;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,108,0,80,0,5,0,0,0,0,0,245,0,184,0,108,0,149,0,199,0,140,0,231,0,0,0,58,0,252,0,146,0,129,0,62,0,30,0,0,0,79,0,246,0,0,0,79,0,210,0,204,0,139,0,0,0,131,0,0,0,9,0,233,0,249,0,215,0,116,0,88,0,101,0,117,0,18,0,0,0,94,0,0,0,15,0,57,0,39,0,62,0,21,0,204,0,3,0,40,0,122,0,201,0,0,0,0,0,26,0,94,0,200,0,196,0,213,0,71,0,202,0,21,0,214,0,0,0,32,0,0,0,138,0,14,0,170,0,17,0,0,0,26,0,0,0,33,0,84,0,30,0,0,0,196,0,0,0,80,0,248,0,107,0,86,0,207,0,126,0,229,0,249,0,96,0,0,0,240,0,155,0,109,0,26,0,149,0,207,0,67,0,14,0,89,0,18,0,0,0,58,0,160,0,70,0,114,0,90,0,0,0,138,0,91,0,199,0,112,0,0,0,36,0,220,0,0,0,0,0,0,0,119,0,204,0,0,0,137,0,177,0,63,0,2,0,2,0,75,0,255,0,70,0,119,0,242,0,193,0,84,0,255,0,219,0,36,0,82,0,60,0,138,0,89,0,0,0,66,0,92,0,19,0,155,0,110,0,0,0,217,0,111,0,230,0,65,0,46,0,251,0,80,0,113,0,0,0,89,0,176,0,0,0,88,0,99,0,116,0,81,0,5,0,142,0,146,0,0,0,0,0,130,0,152,0,162,0,0,0,250,0,22,0,192,0,151,0,126,0,0,0,36,0,208,0,0,0,215,0,72,0,0,0,119,0,91,0,247,0,198,0,0,0,232,0,79,0,140,0,242,0,161,0,185,0,147,0,34,0,12,0,61,0,0,0,157,0,0,0,127,0,117,0,0,0,63,0,48,0,33,0,64,0,0,0,92,0,124,0,157,0,59,0,174,0,167,0,210,0,0,0,77,0,0,0,189,0,245,0,0,0,0,0,248,0,0,0,6,0,56,0,0,0,164,0,145,0,0,0,146,0,0,0,40,0,214,0,227,0,104,0,21,0,157,0,53,0,151,0,6,0,211,0,203,0,198,0,91,0,50,0,206,0,150,0,147,0,0,0,138,0,45,0,51,0,0,0,211,0,0,0,185,0,246,0,151,0,54,0,208,0,120,0,230,0,56,0,49,0,44,0,241,0,93,0,228,0,119,0,1,0,0,0,8,0,240,0,245,0,186,0,222,0,0,0,226,0,17,0,128,0,0,0,236,0,57,0,0,0,209,0,134,0,0,0,37,0,0,0,84,0,109,0,190,0,175,0,149,0,16,0,0,0,64,0,122,0,0,0,30,0,238,0,211,0,245,0,241,0,56,0,68,0,146,0,0,0,245,0,238,0,0,0,0,0,143,0,0,0,172,0,0,0,168,0,0,0,223,0,0,0,0,0,125,0,88,0,78,0,100,0,109,0,0,0,223,0,40,0,188,0,69,0,245,0,232,0,116,0,69,0,106,0,113,0,108,0,229,0,0,0,25,0,252,0,214,0,144,0,124,0,92,0,209,0,157,0,116,0,235,0,0,0,151,0,242,0,134,0,198,0,199,0,0,0,191,0,220,0,187,0,16,0,165,0,108,0,146,0,223,0,217,0,14,0,18,0,158,0,196,0,175,0,30,0,68,0,254,0,6,0,75,0,140,0,157,0,98,0,254,0,0,0,49,0,0,0,95,0,196,0,0,0,39,0,73,0,0,0,0,0,0,0,98,0,61,0,59,0,0,0,0,0,234,0,159,0,0,0,57,0,192,0,78,0,7,0,188,0,0,0,0,0,236,0,0,0,253,0,52,0,0,0,231,0,0,0,0,0,70,0,194,0,250,0,94,0,0,0,31,0,202,0,166,0,126,0,114,0,168,0,108,0,0,0,85,0,104,0,141,0,78,0,0,0,239,0,0,0,215,0,0,0,0,0,201,0,193,0,193,0,97,0,107,0,142,0,139,0,70,0,172,0,221,0,173,0,202,0,98,0,44,0,36,0,0,0,0,0,29,0,84,0,207,0,0,0,193,0,0,0,19,0,34,0,47,0,169,0,221,0,169,0,114,0,230,0,210,0,202,0,226,0,96,0,50,0,51,0,51,0,113,0,0,0,0,0,0,0,7,0,9,0,0,0,103,0,0,0,137,0,125,0,69,0,198,0,125,0,194,0,129,0,0,0,211,0,229,0,131,0,182,0,246,0,1,0,103,0,231,0,0,0,0,0,0,0,0,0,31,0,0,0,204,0,181,0,62,0,251,0,3,0,56,0,210,0,176,0,0,0,34,0,71,0,164,0,68,0,111,0,115,0,29,0,116,0,0,0,202,0,17,0,198,0,177,0,236,0,158,0,89,0,0,0,173,0,47,0,228,0,205,0,71,0,171,0,9,0,30,0,14,0,217,0,140,0,0,0,175,0,155,0,165,0,217,0,0,0,124,0,208,0,16,0,0,0,126,0,123,0,42,0,238,0,8,0,111,0,0,0,193,0,0,0,207,0,135,0,4,0,150,0,44,0,224,0,170,0,101,0,0,0,220,0,0,0,0,0,0,0,37,0,66,0,191,0,241,0,115,0,253,0,0,0,96,0,227,0,82,0,142,0,134,0,0,0,154,0,162,0,92,0,8,0,31,0,185,0,0,0,103,0,202,0,88,0,0,0,185,0,68,0,10,0,0,0,191,0,0,0,245,0,89,0,67,0,128,0,29,0,120,0,189,0,128,0,129,0,128,0,182,0,65,0,56,0,141,0,131,0,32,0,86,0,21,0,197,0,228,0,0,0,0,0,15,0,132,0,0,0,196,0,0,0,246,0,13,0,102,0,220,0,217,0);
signal scenario_full  : scenario_type := (0,0,108,31,80,31,5,31,5,30,5,29,245,31,184,31,108,31,149,31,199,31,140,31,231,31,231,30,58,31,252,31,146,31,129,31,62,31,30,31,30,30,79,31,246,31,246,30,79,31,210,31,204,31,139,31,139,30,131,31,131,30,9,31,233,31,249,31,215,31,116,31,88,31,101,31,117,31,18,31,18,30,94,31,94,30,15,31,57,31,39,31,62,31,21,31,204,31,3,31,40,31,122,31,201,31,201,30,201,29,26,31,94,31,200,31,196,31,213,31,71,31,202,31,21,31,214,31,214,30,32,31,32,30,138,31,14,31,170,31,17,31,17,30,26,31,26,30,33,31,84,31,30,31,30,30,196,31,196,30,80,31,248,31,107,31,86,31,207,31,126,31,229,31,249,31,96,31,96,30,240,31,155,31,109,31,26,31,149,31,207,31,67,31,14,31,89,31,18,31,18,30,58,31,160,31,70,31,114,31,90,31,90,30,138,31,91,31,199,31,112,31,112,30,36,31,220,31,220,30,220,29,220,28,119,31,204,31,204,30,137,31,177,31,63,31,2,31,2,31,75,31,255,31,70,31,119,31,242,31,193,31,84,31,255,31,219,31,36,31,82,31,60,31,138,31,89,31,89,30,66,31,92,31,19,31,155,31,110,31,110,30,217,31,111,31,230,31,65,31,46,31,251,31,80,31,113,31,113,30,89,31,176,31,176,30,88,31,99,31,116,31,81,31,5,31,142,31,146,31,146,30,146,29,130,31,152,31,162,31,162,30,250,31,22,31,192,31,151,31,126,31,126,30,36,31,208,31,208,30,215,31,72,31,72,30,119,31,91,31,247,31,198,31,198,30,232,31,79,31,140,31,242,31,161,31,185,31,147,31,34,31,12,31,61,31,61,30,157,31,157,30,127,31,117,31,117,30,63,31,48,31,33,31,64,31,64,30,92,31,124,31,157,31,59,31,174,31,167,31,210,31,210,30,77,31,77,30,189,31,245,31,245,30,245,29,248,31,248,30,6,31,56,31,56,30,164,31,145,31,145,30,146,31,146,30,40,31,214,31,227,31,104,31,21,31,157,31,53,31,151,31,6,31,211,31,203,31,198,31,91,31,50,31,206,31,150,31,147,31,147,30,138,31,45,31,51,31,51,30,211,31,211,30,185,31,246,31,151,31,54,31,208,31,120,31,230,31,56,31,49,31,44,31,241,31,93,31,228,31,119,31,1,31,1,30,8,31,240,31,245,31,186,31,222,31,222,30,226,31,17,31,128,31,128,30,236,31,57,31,57,30,209,31,134,31,134,30,37,31,37,30,84,31,109,31,190,31,175,31,149,31,16,31,16,30,64,31,122,31,122,30,30,31,238,31,211,31,245,31,241,31,56,31,68,31,146,31,146,30,245,31,238,31,238,30,238,29,143,31,143,30,172,31,172,30,168,31,168,30,223,31,223,30,223,29,125,31,88,31,78,31,100,31,109,31,109,30,223,31,40,31,188,31,69,31,245,31,232,31,116,31,69,31,106,31,113,31,108,31,229,31,229,30,25,31,252,31,214,31,144,31,124,31,92,31,209,31,157,31,116,31,235,31,235,30,151,31,242,31,134,31,198,31,199,31,199,30,191,31,220,31,187,31,16,31,165,31,108,31,146,31,223,31,217,31,14,31,18,31,158,31,196,31,175,31,30,31,68,31,254,31,6,31,75,31,140,31,157,31,98,31,254,31,254,30,49,31,49,30,95,31,196,31,196,30,39,31,73,31,73,30,73,29,73,28,98,31,61,31,59,31,59,30,59,29,234,31,159,31,159,30,57,31,192,31,78,31,7,31,188,31,188,30,188,29,236,31,236,30,253,31,52,31,52,30,231,31,231,30,231,29,70,31,194,31,250,31,94,31,94,30,31,31,202,31,166,31,126,31,114,31,168,31,108,31,108,30,85,31,104,31,141,31,78,31,78,30,239,31,239,30,215,31,215,30,215,29,201,31,193,31,193,31,97,31,107,31,142,31,139,31,70,31,172,31,221,31,173,31,202,31,98,31,44,31,36,31,36,30,36,29,29,31,84,31,207,31,207,30,193,31,193,30,19,31,34,31,47,31,169,31,221,31,169,31,114,31,230,31,210,31,202,31,226,31,96,31,50,31,51,31,51,31,113,31,113,30,113,29,113,28,7,31,9,31,9,30,103,31,103,30,137,31,125,31,69,31,198,31,125,31,194,31,129,31,129,30,211,31,229,31,131,31,182,31,246,31,1,31,103,31,231,31,231,30,231,29,231,28,231,27,31,31,31,30,204,31,181,31,62,31,251,31,3,31,56,31,210,31,176,31,176,30,34,31,71,31,164,31,68,31,111,31,115,31,29,31,116,31,116,30,202,31,17,31,198,31,177,31,236,31,158,31,89,31,89,30,173,31,47,31,228,31,205,31,71,31,171,31,9,31,30,31,14,31,217,31,140,31,140,30,175,31,155,31,165,31,217,31,217,30,124,31,208,31,16,31,16,30,126,31,123,31,42,31,238,31,8,31,111,31,111,30,193,31,193,30,207,31,135,31,4,31,150,31,44,31,224,31,170,31,101,31,101,30,220,31,220,30,220,29,220,28,37,31,66,31,191,31,241,31,115,31,253,31,253,30,96,31,227,31,82,31,142,31,134,31,134,30,154,31,162,31,92,31,8,31,31,31,185,31,185,30,103,31,202,31,88,31,88,30,185,31,68,31,10,31,10,30,191,31,191,30,245,31,89,31,67,31,128,31,29,31,120,31,189,31,128,31,129,31,128,31,182,31,65,31,56,31,141,31,131,31,32,31,86,31,21,31,197,31,228,31,228,30,228,29,15,31,132,31,132,30,196,31,196,30,246,31,13,31,102,31,220,31,217,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
