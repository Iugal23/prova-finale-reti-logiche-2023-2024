-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 931;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (23,0,0,0,108,0,0,0,10,0,217,0,95,0,243,0,83,0,0,0,236,0,158,0,187,0,169,0,105,0,71,0,126,0,207,0,198,0,247,0,47,0,127,0,129,0,0,0,28,0,210,0,206,0,7,0,222,0,0,0,25,0,62,0,40,0,161,0,135,0,190,0,130,0,159,0,250,0,47,0,197,0,171,0,34,0,0,0,235,0,69,0,25,0,0,0,75,0,216,0,147,0,16,0,0,0,3,0,174,0,133,0,72,0,22,0,157,0,174,0,0,0,31,0,140,0,225,0,0,0,159,0,18,0,219,0,87,0,0,0,0,0,0,0,18,0,0,0,0,0,110,0,0,0,112,0,22,0,191,0,137,0,98,0,213,0,90,0,0,0,231,0,244,0,154,0,0,0,138,0,162,0,125,0,179,0,57,0,235,0,0,0,90,0,219,0,200,0,139,0,6,0,162,0,41,0,0,0,67,0,0,0,0,0,247,0,148,0,0,0,20,0,33,0,46,0,0,0,155,0,134,0,231,0,177,0,24,0,63,0,8,0,0,0,247,0,68,0,53,0,206,0,16,0,0,0,69,0,154,0,38,0,245,0,36,0,229,0,66,0,193,0,240,0,108,0,0,0,0,0,49,0,0,0,30,0,29,0,215,0,179,0,193,0,107,0,0,0,78,0,123,0,244,0,92,0,167,0,132,0,85,0,85,0,24,0,229,0,166,0,144,0,176,0,3,0,27,0,61,0,136,0,36,0,221,0,242,0,106,0,118,0,45,0,185,0,0,0,121,0,0,0,0,0,0,0,17,0,34,0,27,0,0,0,112,0,114,0,6,0,168,0,249,0,68,0,0,0,16,0,36,0,0,0,248,0,124,0,46,0,0,0,170,0,189,0,204,0,167,0,77,0,0,0,149,0,203,0,22,0,135,0,67,0,13,0,84,0,87,0,99,0,12,0,161,0,123,0,249,0,235,0,232,0,12,0,0,0,25,0,0,0,153,0,0,0,108,0,0,0,160,0,101,0,242,0,189,0,122,0,0,0,40,0,16,0,158,0,0,0,0,0,149,0,55,0,0,0,242,0,88,0,98,0,24,0,149,0,0,0,176,0,118,0,200,0,19,0,60,0,146,0,36,0,215,0,242,0,120,0,24,0,92,0,81,0,131,0,156,0,79,0,147,0,173,0,66,0,185,0,0,0,121,0,231,0,133,0,0,0,145,0,25,0,101,0,0,0,175,0,0,0,222,0,52,0,139,0,242,0,45,0,49,0,0,0,189,0,17,0,0,0,53,0,136,0,0,0,0,0,0,0,87,0,0,0,203,0,60,0,246,0,184,0,149,0,0,0,0,0,195,0,106,0,94,0,62,0,42,0,225,0,81,0,0,0,16,0,137,0,124,0,0,0,160,0,222,0,0,0,0,0,179,0,20,0,62,0,115,0,191,0,9,0,64,0,0,0,79,0,248,0,231,0,137,0,108,0,145,0,0,0,201,0,104,0,0,0,7,0,169,0,222,0,29,0,0,0,92,0,132,0,107,0,158,0,12,0,0,0,12,0,65,0,163,0,21,0,16,0,226,0,147,0,0,0,242,0,0,0,77,0,92,0,127,0,200,0,36,0,0,0,54,0,212,0,0,0,0,0,0,0,204,0,0,0,232,0,62,0,118,0,204,0,245,0,0,0,124,0,45,0,113,0,41,0,171,0,100,0,132,0,227,0,0,0,138,0,0,0,242,0,91,0,96,0,85,0,241,0,144,0,70,0,75,0,76,0,177,0,106,0,0,0,92,0,180,0,193,0,70,0,87,0,0,0,154,0,88,0,0,0,0,0,243,0,0,0,10,0,117,0,0,0,175,0,243,0,205,0,233,0,197,0,4,0,56,0,195,0,90,0,208,0,166,0,10,0,32,0,128,0,9,0,170,0,0,0,161,0,211,0,146,0,0,0,221,0,0,0,208,0,163,0,208,0,76,0,172,0,125,0,0,0,101,0,75,0,0,0,0,0,207,0,216,0,227,0,183,0,0,0,0,0,244,0,159,0,166,0,30,0,148,0,13,0,229,0,141,0,55,0,72,0,119,0,10,0,100,0,27,0,77,0,113,0,0,0,100,0,0,0,54,0,2,0,0,0,250,0,0,0,0,0,253,0,144,0,4,0,223,0,0,0,23,0,63,0,0,0,253,0,177,0,103,0,231,0,0,0,113,0,10,0,91,0,48,0,227,0,214,0,243,0,30,0,246,0,84,0,203,0,250,0,101,0,0,0,0,0,43,0,205,0,0,0,76,0,107,0,227,0,17,0,8,0,0,0,232,0,12,0,198,0,0,0,24,0,108,0,229,0,225,0,0,0,0,0,240,0,251,0,0,0,0,0,248,0,237,0,111,0,133,0,0,0,177,0,0,0,217,0,157,0,35,0,246,0,213,0,0,0,161,0,27,0,141,0,180,0,106,0,197,0,130,0,16,0,88,0,132,0,208,0,0,0,171,0,51,0,152,0,225,0,49,0,0,0,20,0,213,0,16,0,55,0,242,0,225,0,175,0,8,0,0,0,247,0,0,0,0,0,104,0,45,0,26,0,2,0,155,0,11,0,44,0,41,0,116,0,0,0,206,0,0,0,79,0,164,0,201,0,174,0,64,0,145,0,222,0,248,0,216,0,207,0,28,0,0,0,0,0,245,0,214,0,57,0,243,0,11,0,0,0,89,0,206,0,62,0,0,0,0,0,251,0,0,0,227,0,0,0,0,0,78,0,53,0,129,0,184,0,91,0,64,0,92,0,0,0,0,0,164,0,142,0,0,0,0,0,0,0,72,0,166,0,0,0,21,0,171,0,20,0,0,0,226,0,61,0,167,0,18,0,0,0,250,0,0,0,144,0,0,0,14,0,130,0,188,0,205,0,86,0,109,0,0,0,0,0,94,0,0,0,70,0,75,0,75,0,200,0,42,0,151,0,207,0,166,0,2,0,0,0,13,0,44,0,176,0,74,0,123,0,111,0,218,0,0,0,141,0,10,0,33,0,0,0,0,0,175,0,47,0,0,0,0,0,0,0,212,0,0,0,70,0,254,0,0,0,16,0,229,0,0,0,248,0,57,0,248,0,32,0,53,0,29,0,30,0,107,0,13,0,81,0,105,0,91,0,171,0,194,0,60,0,142,0,159,0,0,0,143,0,0,0,22,0,48,0,56,0,137,0,151,0,1,0,191,0,10,0,209,0,50,0,145,0,212,0,107,0,53,0,0,0,2,0,234,0,126,0,0,0,0,0,134,0,24,0,99,0,229,0,235,0,221,0,176,0,124,0,2,0,15,0,45,0,17,0,168,0,169,0,189,0,64,0,108,0,25,0,210,0,234,0,33,0,30,0,45,0,132,0,93,0,101,0,235,0,186,0,245,0,38,0,216,0,192,0,97,0,204,0,0,0,0,0,35,0,207,0,26,0,192,0,39,0,46,0,50,0,0,0,120,0,186,0,116,0,124,0,64,0,76,0,28,0,61,0,54,0,174,0,111,0,0,0,41,0,111,0,235,0,75,0,231,0,32,0,0,0,17,0,192,0,181,0,142,0,100,0,0,0,0,0,76,0,39,0,49,0,156,0,102,0,0,0,185,0,28,0,150,0,0,0,224,0,0,0,32,0,0,0,23,0,0,0,68,0,0,0,7,0,223,0,189,0,107,0,70,0,220,0,0,0,93,0,0,0,98,0,23,0,183,0,133,0,52,0,254,0,40,0,227,0,13,0,44,0,0,0,80,0,2,0,207,0,11,0,20,0,204,0,32,0,158,0,175,0,111,0,141,0,179,0,231,0,0,0,71,0,36,0,182,0,0,0,0,0,233,0,155,0,87,0,0,0,203,0,101,0,133,0,42,0,129,0,24,0,32,0,186,0,245,0,0,0,144,0,178,0,21,0,0,0,159,0,230,0,60,0,0,0,219,0,229,0,10,0,210,0,241,0,69,0,204,0,81,0,255,0,0,0,83,0,0,0,148,0,218,0,0,0,221,0,0,0,0,0,0,0,144,0,40,0,22,0,216,0,110,0,179,0,134,0,199,0,0,0,0,0,216,0,105,0,143,0,105,0,153,0,193,0,51,0,17,0,100,0,150,0,132,0,51,0,54,0,156,0,0,0,189,0,197,0,0,0,65,0,0,0,234,0,0,0,0,0,0,0,174,0);
signal scenario_full  : scenario_type := (23,31,23,30,108,31,108,30,10,31,217,31,95,31,243,31,83,31,83,30,236,31,158,31,187,31,169,31,105,31,71,31,126,31,207,31,198,31,247,31,47,31,127,31,129,31,129,30,28,31,210,31,206,31,7,31,222,31,222,30,25,31,62,31,40,31,161,31,135,31,190,31,130,31,159,31,250,31,47,31,197,31,171,31,34,31,34,30,235,31,69,31,25,31,25,30,75,31,216,31,147,31,16,31,16,30,3,31,174,31,133,31,72,31,22,31,157,31,174,31,174,30,31,31,140,31,225,31,225,30,159,31,18,31,219,31,87,31,87,30,87,29,87,28,18,31,18,30,18,29,110,31,110,30,112,31,22,31,191,31,137,31,98,31,213,31,90,31,90,30,231,31,244,31,154,31,154,30,138,31,162,31,125,31,179,31,57,31,235,31,235,30,90,31,219,31,200,31,139,31,6,31,162,31,41,31,41,30,67,31,67,30,67,29,247,31,148,31,148,30,20,31,33,31,46,31,46,30,155,31,134,31,231,31,177,31,24,31,63,31,8,31,8,30,247,31,68,31,53,31,206,31,16,31,16,30,69,31,154,31,38,31,245,31,36,31,229,31,66,31,193,31,240,31,108,31,108,30,108,29,49,31,49,30,30,31,29,31,215,31,179,31,193,31,107,31,107,30,78,31,123,31,244,31,92,31,167,31,132,31,85,31,85,31,24,31,229,31,166,31,144,31,176,31,3,31,27,31,61,31,136,31,36,31,221,31,242,31,106,31,118,31,45,31,185,31,185,30,121,31,121,30,121,29,121,28,17,31,34,31,27,31,27,30,112,31,114,31,6,31,168,31,249,31,68,31,68,30,16,31,36,31,36,30,248,31,124,31,46,31,46,30,170,31,189,31,204,31,167,31,77,31,77,30,149,31,203,31,22,31,135,31,67,31,13,31,84,31,87,31,99,31,12,31,161,31,123,31,249,31,235,31,232,31,12,31,12,30,25,31,25,30,153,31,153,30,108,31,108,30,160,31,101,31,242,31,189,31,122,31,122,30,40,31,16,31,158,31,158,30,158,29,149,31,55,31,55,30,242,31,88,31,98,31,24,31,149,31,149,30,176,31,118,31,200,31,19,31,60,31,146,31,36,31,215,31,242,31,120,31,24,31,92,31,81,31,131,31,156,31,79,31,147,31,173,31,66,31,185,31,185,30,121,31,231,31,133,31,133,30,145,31,25,31,101,31,101,30,175,31,175,30,222,31,52,31,139,31,242,31,45,31,49,31,49,30,189,31,17,31,17,30,53,31,136,31,136,30,136,29,136,28,87,31,87,30,203,31,60,31,246,31,184,31,149,31,149,30,149,29,195,31,106,31,94,31,62,31,42,31,225,31,81,31,81,30,16,31,137,31,124,31,124,30,160,31,222,31,222,30,222,29,179,31,20,31,62,31,115,31,191,31,9,31,64,31,64,30,79,31,248,31,231,31,137,31,108,31,145,31,145,30,201,31,104,31,104,30,7,31,169,31,222,31,29,31,29,30,92,31,132,31,107,31,158,31,12,31,12,30,12,31,65,31,163,31,21,31,16,31,226,31,147,31,147,30,242,31,242,30,77,31,92,31,127,31,200,31,36,31,36,30,54,31,212,31,212,30,212,29,212,28,204,31,204,30,232,31,62,31,118,31,204,31,245,31,245,30,124,31,45,31,113,31,41,31,171,31,100,31,132,31,227,31,227,30,138,31,138,30,242,31,91,31,96,31,85,31,241,31,144,31,70,31,75,31,76,31,177,31,106,31,106,30,92,31,180,31,193,31,70,31,87,31,87,30,154,31,88,31,88,30,88,29,243,31,243,30,10,31,117,31,117,30,175,31,243,31,205,31,233,31,197,31,4,31,56,31,195,31,90,31,208,31,166,31,10,31,32,31,128,31,9,31,170,31,170,30,161,31,211,31,146,31,146,30,221,31,221,30,208,31,163,31,208,31,76,31,172,31,125,31,125,30,101,31,75,31,75,30,75,29,207,31,216,31,227,31,183,31,183,30,183,29,244,31,159,31,166,31,30,31,148,31,13,31,229,31,141,31,55,31,72,31,119,31,10,31,100,31,27,31,77,31,113,31,113,30,100,31,100,30,54,31,2,31,2,30,250,31,250,30,250,29,253,31,144,31,4,31,223,31,223,30,23,31,63,31,63,30,253,31,177,31,103,31,231,31,231,30,113,31,10,31,91,31,48,31,227,31,214,31,243,31,30,31,246,31,84,31,203,31,250,31,101,31,101,30,101,29,43,31,205,31,205,30,76,31,107,31,227,31,17,31,8,31,8,30,232,31,12,31,198,31,198,30,24,31,108,31,229,31,225,31,225,30,225,29,240,31,251,31,251,30,251,29,248,31,237,31,111,31,133,31,133,30,177,31,177,30,217,31,157,31,35,31,246,31,213,31,213,30,161,31,27,31,141,31,180,31,106,31,197,31,130,31,16,31,88,31,132,31,208,31,208,30,171,31,51,31,152,31,225,31,49,31,49,30,20,31,213,31,16,31,55,31,242,31,225,31,175,31,8,31,8,30,247,31,247,30,247,29,104,31,45,31,26,31,2,31,155,31,11,31,44,31,41,31,116,31,116,30,206,31,206,30,79,31,164,31,201,31,174,31,64,31,145,31,222,31,248,31,216,31,207,31,28,31,28,30,28,29,245,31,214,31,57,31,243,31,11,31,11,30,89,31,206,31,62,31,62,30,62,29,251,31,251,30,227,31,227,30,227,29,78,31,53,31,129,31,184,31,91,31,64,31,92,31,92,30,92,29,164,31,142,31,142,30,142,29,142,28,72,31,166,31,166,30,21,31,171,31,20,31,20,30,226,31,61,31,167,31,18,31,18,30,250,31,250,30,144,31,144,30,14,31,130,31,188,31,205,31,86,31,109,31,109,30,109,29,94,31,94,30,70,31,75,31,75,31,200,31,42,31,151,31,207,31,166,31,2,31,2,30,13,31,44,31,176,31,74,31,123,31,111,31,218,31,218,30,141,31,10,31,33,31,33,30,33,29,175,31,47,31,47,30,47,29,47,28,212,31,212,30,70,31,254,31,254,30,16,31,229,31,229,30,248,31,57,31,248,31,32,31,53,31,29,31,30,31,107,31,13,31,81,31,105,31,91,31,171,31,194,31,60,31,142,31,159,31,159,30,143,31,143,30,22,31,48,31,56,31,137,31,151,31,1,31,191,31,10,31,209,31,50,31,145,31,212,31,107,31,53,31,53,30,2,31,234,31,126,31,126,30,126,29,134,31,24,31,99,31,229,31,235,31,221,31,176,31,124,31,2,31,15,31,45,31,17,31,168,31,169,31,189,31,64,31,108,31,25,31,210,31,234,31,33,31,30,31,45,31,132,31,93,31,101,31,235,31,186,31,245,31,38,31,216,31,192,31,97,31,204,31,204,30,204,29,35,31,207,31,26,31,192,31,39,31,46,31,50,31,50,30,120,31,186,31,116,31,124,31,64,31,76,31,28,31,61,31,54,31,174,31,111,31,111,30,41,31,111,31,235,31,75,31,231,31,32,31,32,30,17,31,192,31,181,31,142,31,100,31,100,30,100,29,76,31,39,31,49,31,156,31,102,31,102,30,185,31,28,31,150,31,150,30,224,31,224,30,32,31,32,30,23,31,23,30,68,31,68,30,7,31,223,31,189,31,107,31,70,31,220,31,220,30,93,31,93,30,98,31,23,31,183,31,133,31,52,31,254,31,40,31,227,31,13,31,44,31,44,30,80,31,2,31,207,31,11,31,20,31,204,31,32,31,158,31,175,31,111,31,141,31,179,31,231,31,231,30,71,31,36,31,182,31,182,30,182,29,233,31,155,31,87,31,87,30,203,31,101,31,133,31,42,31,129,31,24,31,32,31,186,31,245,31,245,30,144,31,178,31,21,31,21,30,159,31,230,31,60,31,60,30,219,31,229,31,10,31,210,31,241,31,69,31,204,31,81,31,255,31,255,30,83,31,83,30,148,31,218,31,218,30,221,31,221,30,221,29,221,28,144,31,40,31,22,31,216,31,110,31,179,31,134,31,199,31,199,30,199,29,216,31,105,31,143,31,105,31,153,31,193,31,51,31,17,31,100,31,150,31,132,31,51,31,54,31,156,31,156,30,189,31,197,31,197,30,65,31,65,30,234,31,234,30,234,29,234,28,174,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
