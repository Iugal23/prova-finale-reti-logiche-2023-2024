-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_943 is
end project_tb_943;

architecture project_tb_arch_943 of project_tb_943 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 716;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (243,0,0,0,251,0,108,0,227,0,199,0,156,0,61,0,105,0,104,0,0,0,40,0,213,0,16,0,54,0,121,0,133,0,244,0,113,0,8,0,0,0,88,0,58,0,0,0,0,0,246,0,77,0,101,0,142,0,217,0,36,0,222,0,169,0,0,0,162,0,67,0,0,0,130,0,27,0,167,0,5,0,229,0,106,0,95,0,187,0,187,0,202,0,73,0,1,0,128,0,57,0,73,0,193,0,71,0,0,0,196,0,22,0,137,0,194,0,108,0,0,0,50,0,167,0,15,0,241,0,239,0,43,0,247,0,254,0,127,0,165,0,35,0,204,0,0,0,0,0,119,0,109,0,0,0,134,0,175,0,75,0,155,0,0,0,92,0,66,0,208,0,239,0,76,0,0,0,7,0,133,0,0,0,0,0,89,0,146,0,0,0,197,0,16,0,159,0,97,0,178,0,6,0,108,0,246,0,103,0,236,0,46,0,47,0,38,0,0,0,223,0,53,0,0,0,200,0,208,0,0,0,9,0,65,0,35,0,0,0,222,0,99,0,0,0,158,0,215,0,0,0,197,0,0,0,219,0,40,0,228,0,55,0,16,0,202,0,34,0,22,0,17,0,236,0,146,0,56,0,158,0,71,0,0,0,0,0,175,0,142,0,171,0,197,0,0,0,120,0,147,0,22,0,226,0,117,0,139,0,114,0,251,0,187,0,22,0,178,0,28,0,114,0,163,0,0,0,96,0,92,0,47,0,197,0,12,0,0,0,232,0,161,0,156,0,253,0,239,0,217,0,77,0,201,0,0,0,212,0,120,0,208,0,0,0,246,0,0,0,148,0,0,0,0,0,249,0,0,0,108,0,222,0,35,0,147,0,196,0,52,0,103,0,36,0,75,0,136,0,218,0,100,0,10,0,47,0,0,0,188,0,29,0,0,0,72,0,112,0,0,0,11,0,94,0,0,0,0,0,0,0,0,0,0,0,80,0,160,0,191,0,68,0,168,0,104,0,123,0,66,0,137,0,0,0,138,0,129,0,0,0,95,0,33,0,0,0,112,0,0,0,0,0,68,0,139,0,119,0,112,0,43,0,53,0,0,0,197,0,89,0,233,0,74,0,178,0,235,0,54,0,0,0,53,0,7,0,201,0,0,0,212,0,239,0,126,0,54,0,54,0,214,0,0,0,0,0,0,0,143,0,41,0,136,0,147,0,178,0,29,0,173,0,159,0,51,0,192,0,42,0,166,0,0,0,226,0,166,0,182,0,70,0,0,0,171,0,116,0,38,0,167,0,228,0,187,0,162,0,0,0,107,0,175,0,199,0,135,0,172,0,131,0,43,0,88,0,0,0,56,0,185,0,182,0,239,0,156,0,5,0,95,0,247,0,63,0,43,0,0,0,0,0,71,0,77,0,148,0,162,0,32,0,113,0,195,0,0,0,116,0,0,0,187,0,140,0,235,0,66,0,235,0,183,0,0,0,194,0,0,0,20,0,227,0,0,0,214,0,106,0,125,0,100,0,21,0,243,0,200,0,176,0,176,0,0,0,211,0,0,0,0,0,162,0,181,0,163,0,216,0,0,0,167,0,63,0,43,0,33,0,176,0,0,0,130,0,107,0,235,0,174,0,66,0,163,0,223,0,222,0,163,0,86,0,61,0,195,0,131,0,0,0,0,0,253,0,181,0,23,0,235,0,224,0,241,0,30,0,9,0,0,0,214,0,162,0,0,0,236,0,164,0,78,0,0,0,66,0,190,0,153,0,41,0,231,0,239,0,227,0,52,0,242,0,65,0,111,0,179,0,1,0,90,0,186,0,202,0,215,0,0,0,0,0,0,0,181,0,164,0,132,0,125,0,0,0,129,0,201,0,0,0,107,0,80,0,62,0,170,0,75,0,143,0,244,0,89,0,74,0,0,0,0,0,77,0,117,0,197,0,105,0,195,0,214,0,27,0,98,0,212,0,234,0,0,0,160,0,155,0,18,0,0,0,24,0,174,0,223,0,0,0,0,0,135,0,203,0,118,0,0,0,132,0,0,0,0,0,225,0,85,0,97,0,74,0,53,0,0,0,74,0,0,0,142,0,85,0,46,0,0,0,56,0,243,0,184,0,0,0,189,0,21,0,0,0,249,0,114,0,50,0,183,0,64,0,251,0,172,0,253,0,126,0,0,0,180,0,173,0,180,0,174,0,130,0,213,0,14,0,0,0,97,0,132,0,7,0,0,0,0,0,214,0,185,0,44,0,0,0,101,0,148,0,118,0,110,0,0,0,0,0,160,0,215,0,190,0,237,0,194,0,3,0,127,0,239,0,219,0,0,0,78,0,0,0,166,0,214,0,150,0,136,0,25,0,215,0,0,0,9,0,175,0,54,0,248,0,78,0,177,0,213,0,15,0,155,0,194,0,0,0,221,0,163,0,131,0,126,0,63,0,240,0,86,0,0,0,15,0,249,0,227,0,245,0,235,0,140,0,118,0,0,0,213,0,59,0,234,0,0,0,61,0,244,0,0,0,200,0,213,0,32,0,196,0,0,0,0,0,231,0,45,0,178,0,127,0,87,0,88,0,0,0,192,0,0,0,13,0,147,0,169,0,0,0,66,0,138,0,16,0,175,0,205,0,94,0,138,0,54,0,61,0,50,0,97,0,199,0,0,0,0,0,20,0,0,0,65,0,0,0,217,0,180,0,31,0,0,0,236,0,77,0,172,0,0,0,0,0,197,0,81,0,195,0,189,0,85,0,214,0,105,0,88,0,119,0,156,0,119,0,206,0,185,0,68,0,0,0,92,0,26,0,0,0,127,0,0,0,68,0,161,0,72,0,89,0,241,0,114,0,254,0,243,0,115,0,133,0,42,0,44,0,178,0,0,0,0,0,90,0,0,0,205,0,215,0,0,0,54,0,0,0,117,0,154,0,253,0,142,0,5,0,0,0,60,0,207,0,167,0,138,0,177,0,0,0,0,0,116,0,131,0,0,0,36,0,218,0,0,0,124,0,0,0,0,0,0,0,0,0,61,0,51,0,190,0,0,0,240,0,62,0,21,0,0,0,203,0,81,0,71,0,0,0,56,0,0,0,37,0,190,0,0,0,84,0,93,0,0,0,0,0,0,0,127,0,0,0,38,0,250,0,5,0,0,0,0,0,204,0,176,0,215,0,79,0,104,0,128,0,1,0,108,0,235,0,238,0,228,0,104,0,42,0,142,0,165,0);
signal scenario_full  : scenario_type := (243,31,243,30,251,31,108,31,227,31,199,31,156,31,61,31,105,31,104,31,104,30,40,31,213,31,16,31,54,31,121,31,133,31,244,31,113,31,8,31,8,30,88,31,58,31,58,30,58,29,246,31,77,31,101,31,142,31,217,31,36,31,222,31,169,31,169,30,162,31,67,31,67,30,130,31,27,31,167,31,5,31,229,31,106,31,95,31,187,31,187,31,202,31,73,31,1,31,128,31,57,31,73,31,193,31,71,31,71,30,196,31,22,31,137,31,194,31,108,31,108,30,50,31,167,31,15,31,241,31,239,31,43,31,247,31,254,31,127,31,165,31,35,31,204,31,204,30,204,29,119,31,109,31,109,30,134,31,175,31,75,31,155,31,155,30,92,31,66,31,208,31,239,31,76,31,76,30,7,31,133,31,133,30,133,29,89,31,146,31,146,30,197,31,16,31,159,31,97,31,178,31,6,31,108,31,246,31,103,31,236,31,46,31,47,31,38,31,38,30,223,31,53,31,53,30,200,31,208,31,208,30,9,31,65,31,35,31,35,30,222,31,99,31,99,30,158,31,215,31,215,30,197,31,197,30,219,31,40,31,228,31,55,31,16,31,202,31,34,31,22,31,17,31,236,31,146,31,56,31,158,31,71,31,71,30,71,29,175,31,142,31,171,31,197,31,197,30,120,31,147,31,22,31,226,31,117,31,139,31,114,31,251,31,187,31,22,31,178,31,28,31,114,31,163,31,163,30,96,31,92,31,47,31,197,31,12,31,12,30,232,31,161,31,156,31,253,31,239,31,217,31,77,31,201,31,201,30,212,31,120,31,208,31,208,30,246,31,246,30,148,31,148,30,148,29,249,31,249,30,108,31,222,31,35,31,147,31,196,31,52,31,103,31,36,31,75,31,136,31,218,31,100,31,10,31,47,31,47,30,188,31,29,31,29,30,72,31,112,31,112,30,11,31,94,31,94,30,94,29,94,28,94,27,94,26,80,31,160,31,191,31,68,31,168,31,104,31,123,31,66,31,137,31,137,30,138,31,129,31,129,30,95,31,33,31,33,30,112,31,112,30,112,29,68,31,139,31,119,31,112,31,43,31,53,31,53,30,197,31,89,31,233,31,74,31,178,31,235,31,54,31,54,30,53,31,7,31,201,31,201,30,212,31,239,31,126,31,54,31,54,31,214,31,214,30,214,29,214,28,143,31,41,31,136,31,147,31,178,31,29,31,173,31,159,31,51,31,192,31,42,31,166,31,166,30,226,31,166,31,182,31,70,31,70,30,171,31,116,31,38,31,167,31,228,31,187,31,162,31,162,30,107,31,175,31,199,31,135,31,172,31,131,31,43,31,88,31,88,30,56,31,185,31,182,31,239,31,156,31,5,31,95,31,247,31,63,31,43,31,43,30,43,29,71,31,77,31,148,31,162,31,32,31,113,31,195,31,195,30,116,31,116,30,187,31,140,31,235,31,66,31,235,31,183,31,183,30,194,31,194,30,20,31,227,31,227,30,214,31,106,31,125,31,100,31,21,31,243,31,200,31,176,31,176,31,176,30,211,31,211,30,211,29,162,31,181,31,163,31,216,31,216,30,167,31,63,31,43,31,33,31,176,31,176,30,130,31,107,31,235,31,174,31,66,31,163,31,223,31,222,31,163,31,86,31,61,31,195,31,131,31,131,30,131,29,253,31,181,31,23,31,235,31,224,31,241,31,30,31,9,31,9,30,214,31,162,31,162,30,236,31,164,31,78,31,78,30,66,31,190,31,153,31,41,31,231,31,239,31,227,31,52,31,242,31,65,31,111,31,179,31,1,31,90,31,186,31,202,31,215,31,215,30,215,29,215,28,181,31,164,31,132,31,125,31,125,30,129,31,201,31,201,30,107,31,80,31,62,31,170,31,75,31,143,31,244,31,89,31,74,31,74,30,74,29,77,31,117,31,197,31,105,31,195,31,214,31,27,31,98,31,212,31,234,31,234,30,160,31,155,31,18,31,18,30,24,31,174,31,223,31,223,30,223,29,135,31,203,31,118,31,118,30,132,31,132,30,132,29,225,31,85,31,97,31,74,31,53,31,53,30,74,31,74,30,142,31,85,31,46,31,46,30,56,31,243,31,184,31,184,30,189,31,21,31,21,30,249,31,114,31,50,31,183,31,64,31,251,31,172,31,253,31,126,31,126,30,180,31,173,31,180,31,174,31,130,31,213,31,14,31,14,30,97,31,132,31,7,31,7,30,7,29,214,31,185,31,44,31,44,30,101,31,148,31,118,31,110,31,110,30,110,29,160,31,215,31,190,31,237,31,194,31,3,31,127,31,239,31,219,31,219,30,78,31,78,30,166,31,214,31,150,31,136,31,25,31,215,31,215,30,9,31,175,31,54,31,248,31,78,31,177,31,213,31,15,31,155,31,194,31,194,30,221,31,163,31,131,31,126,31,63,31,240,31,86,31,86,30,15,31,249,31,227,31,245,31,235,31,140,31,118,31,118,30,213,31,59,31,234,31,234,30,61,31,244,31,244,30,200,31,213,31,32,31,196,31,196,30,196,29,231,31,45,31,178,31,127,31,87,31,88,31,88,30,192,31,192,30,13,31,147,31,169,31,169,30,66,31,138,31,16,31,175,31,205,31,94,31,138,31,54,31,61,31,50,31,97,31,199,31,199,30,199,29,20,31,20,30,65,31,65,30,217,31,180,31,31,31,31,30,236,31,77,31,172,31,172,30,172,29,197,31,81,31,195,31,189,31,85,31,214,31,105,31,88,31,119,31,156,31,119,31,206,31,185,31,68,31,68,30,92,31,26,31,26,30,127,31,127,30,68,31,161,31,72,31,89,31,241,31,114,31,254,31,243,31,115,31,133,31,42,31,44,31,178,31,178,30,178,29,90,31,90,30,205,31,215,31,215,30,54,31,54,30,117,31,154,31,253,31,142,31,5,31,5,30,60,31,207,31,167,31,138,31,177,31,177,30,177,29,116,31,131,31,131,30,36,31,218,31,218,30,124,31,124,30,124,29,124,28,124,27,61,31,51,31,190,31,190,30,240,31,62,31,21,31,21,30,203,31,81,31,71,31,71,30,56,31,56,30,37,31,190,31,190,30,84,31,93,31,93,30,93,29,93,28,127,31,127,30,38,31,250,31,5,31,5,30,5,29,204,31,176,31,215,31,79,31,104,31,128,31,1,31,108,31,235,31,238,31,228,31,104,31,42,31,142,31,165,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
