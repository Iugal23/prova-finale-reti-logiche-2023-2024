-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 394;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (87,0,183,0,30,0,74,0,0,0,0,0,0,0,0,0,161,0,140,0,43,0,13,0,208,0,153,0,52,0,149,0,0,0,0,0,5,0,166,0,201,0,119,0,23,0,23,0,0,0,254,0,157,0,250,0,55,0,0,0,28,0,241,0,0,0,0,0,242,0,186,0,74,0,113,0,19,0,13,0,96,0,114,0,53,0,127,0,233,0,220,0,196,0,227,0,0,0,183,0,28,0,252,0,0,0,221,0,98,0,230,0,0,0,0,0,6,0,165,0,124,0,251,0,81,0,35,0,20,0,56,0,131,0,0,0,128,0,0,0,26,0,180,0,103,0,250,0,179,0,98,0,50,0,72,0,3,0,81,0,215,0,247,0,0,0,0,0,1,0,38,0,170,0,250,0,137,0,45,0,1,0,16,0,43,0,220,0,22,0,50,0,57,0,0,0,212,0,244,0,93,0,235,0,32,0,76,0,249,0,0,0,237,0,122,0,7,0,0,0,72,0,70,0,173,0,243,0,86,0,0,0,0,0,233,0,39,0,0,0,166,0,0,0,0,0,148,0,0,0,247,0,0,0,104,0,139,0,151,0,138,0,249,0,24,0,0,0,112,0,0,0,65,0,145,0,0,0,3,0,120,0,142,0,33,0,0,0,22,0,59,0,0,0,232,0,106,0,100,0,202,0,168,0,0,0,207,0,48,0,0,0,61,0,43,0,0,0,250,0,50,0,227,0,235,0,191,0,187,0,207,0,127,0,128,0,62,0,33,0,59,0,157,0,127,0,106,0,19,0,56,0,0,0,163,0,0,0,42,0,236,0,0,0,153,0,105,0,39,0,163,0,0,0,28,0,46,0,208,0,202,0,0,0,71,0,251,0,135,0,132,0,0,0,53,0,224,0,66,0,74,0,117,0,240,0,158,0,40,0,150,0,0,0,221,0,129,0,0,0,164,0,241,0,0,0,35,0,24,0,160,0,177,0,0,0,35,0,0,0,0,0,88,0,0,0,22,0,23,0,0,0,155,0,40,0,17,0,152,0,0,0,0,0,55,0,226,0,0,0,100,0,195,0,14,0,203,0,61,0,0,0,0,0,19,0,230,0,7,0,59,0,244,0,37,0,225,0,227,0,23,0,69,0,220,0,155,0,211,0,170,0,52,0,29,0,0,0,19,0,191,0,73,0,80,0,150,0,0,0,77,0,0,0,250,0,141,0,222,0,126,0,217,0,186,0,94,0,211,0,251,0,222,0,0,0,55,0,188,0,165,0,0,0,38,0,160,0,37,0,0,0,5,0,225,0,153,0,0,0,88,0,193,0,43,0,51,0,246,0,228,0,0,0,179,0,143,0,216,0,26,0,0,0,65,0,0,0,5,0,165,0,34,0,183,0,102,0,0,0,170,0,173,0,190,0,151,0,46,0,61,0,0,0,219,0,16,0,193,0,106,0,12,0,64,0,0,0,184,0,97,0,199,0,43,0,0,0,9,0,157,0,45,0,250,0,65,0,242,0,12,0,248,0,84,0,0,0,203,0,6,0,225,0,143,0,133,0,93,0,0,0,45,0,0,0,205,0,55,0,136,0,63,0,0,0,0,0,64,0,50,0,245,0,199,0,6,0,166,0,248,0,226,0,18,0,159,0,235,0,154,0,218,0,205,0,104,0,238,0,218,0,0,0,230,0,1,0,27,0,177,0,0,0,0,0,79,0,219,0,0,0,144,0,134,0,19,0,166,0,0,0,141,0,247,0,0,0,147,0,52,0,18,0,41,0,0,0);
signal scenario_full  : scenario_type := (87,31,183,31,30,31,74,31,74,30,74,29,74,28,74,27,161,31,140,31,43,31,13,31,208,31,153,31,52,31,149,31,149,30,149,29,5,31,166,31,201,31,119,31,23,31,23,31,23,30,254,31,157,31,250,31,55,31,55,30,28,31,241,31,241,30,241,29,242,31,186,31,74,31,113,31,19,31,13,31,96,31,114,31,53,31,127,31,233,31,220,31,196,31,227,31,227,30,183,31,28,31,252,31,252,30,221,31,98,31,230,31,230,30,230,29,6,31,165,31,124,31,251,31,81,31,35,31,20,31,56,31,131,31,131,30,128,31,128,30,26,31,180,31,103,31,250,31,179,31,98,31,50,31,72,31,3,31,81,31,215,31,247,31,247,30,247,29,1,31,38,31,170,31,250,31,137,31,45,31,1,31,16,31,43,31,220,31,22,31,50,31,57,31,57,30,212,31,244,31,93,31,235,31,32,31,76,31,249,31,249,30,237,31,122,31,7,31,7,30,72,31,70,31,173,31,243,31,86,31,86,30,86,29,233,31,39,31,39,30,166,31,166,30,166,29,148,31,148,30,247,31,247,30,104,31,139,31,151,31,138,31,249,31,24,31,24,30,112,31,112,30,65,31,145,31,145,30,3,31,120,31,142,31,33,31,33,30,22,31,59,31,59,30,232,31,106,31,100,31,202,31,168,31,168,30,207,31,48,31,48,30,61,31,43,31,43,30,250,31,50,31,227,31,235,31,191,31,187,31,207,31,127,31,128,31,62,31,33,31,59,31,157,31,127,31,106,31,19,31,56,31,56,30,163,31,163,30,42,31,236,31,236,30,153,31,105,31,39,31,163,31,163,30,28,31,46,31,208,31,202,31,202,30,71,31,251,31,135,31,132,31,132,30,53,31,224,31,66,31,74,31,117,31,240,31,158,31,40,31,150,31,150,30,221,31,129,31,129,30,164,31,241,31,241,30,35,31,24,31,160,31,177,31,177,30,35,31,35,30,35,29,88,31,88,30,22,31,23,31,23,30,155,31,40,31,17,31,152,31,152,30,152,29,55,31,226,31,226,30,100,31,195,31,14,31,203,31,61,31,61,30,61,29,19,31,230,31,7,31,59,31,244,31,37,31,225,31,227,31,23,31,69,31,220,31,155,31,211,31,170,31,52,31,29,31,29,30,19,31,191,31,73,31,80,31,150,31,150,30,77,31,77,30,250,31,141,31,222,31,126,31,217,31,186,31,94,31,211,31,251,31,222,31,222,30,55,31,188,31,165,31,165,30,38,31,160,31,37,31,37,30,5,31,225,31,153,31,153,30,88,31,193,31,43,31,51,31,246,31,228,31,228,30,179,31,143,31,216,31,26,31,26,30,65,31,65,30,5,31,165,31,34,31,183,31,102,31,102,30,170,31,173,31,190,31,151,31,46,31,61,31,61,30,219,31,16,31,193,31,106,31,12,31,64,31,64,30,184,31,97,31,199,31,43,31,43,30,9,31,157,31,45,31,250,31,65,31,242,31,12,31,248,31,84,31,84,30,203,31,6,31,225,31,143,31,133,31,93,31,93,30,45,31,45,30,205,31,55,31,136,31,63,31,63,30,63,29,64,31,50,31,245,31,199,31,6,31,166,31,248,31,226,31,18,31,159,31,235,31,154,31,218,31,205,31,104,31,238,31,218,31,218,30,230,31,1,31,27,31,177,31,177,30,177,29,79,31,219,31,219,30,144,31,134,31,19,31,166,31,166,30,141,31,247,31,247,30,147,31,52,31,18,31,41,31,41,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
