-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 438;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (168,0,91,0,132,0,191,0,0,0,0,0,91,0,86,0,150,0,187,0,107,0,75,0,3,0,17,0,168,0,184,0,50,0,155,0,53,0,159,0,81,0,149,0,55,0,0,0,131,0,119,0,0,0,32,0,0,0,239,0,204,0,147,0,3,0,208,0,160,0,254,0,184,0,13,0,0,0,116,0,90,0,247,0,0,0,203,0,0,0,0,0,167,0,97,0,228,0,212,0,95,0,0,0,0,0,197,0,63,0,0,0,129,0,0,0,103,0,88,0,126,0,134,0,61,0,191,0,249,0,65,0,57,0,255,0,190,0,57,0,216,0,18,0,94,0,0,0,252,0,32,0,149,0,17,0,168,0,65,0,217,0,239,0,0,0,177,0,102,0,202,0,87,0,0,0,0,0,166,0,233,0,176,0,38,0,58,0,0,0,114,0,68,0,189,0,36,0,104,0,244,0,86,0,210,0,111,0,84,0,188,0,29,0,73,0,217,0,155,0,116,0,209,0,228,0,0,0,119,0,146,0,183,0,50,0,0,0,166,0,0,0,95,0,0,0,8,0,208,0,173,0,231,0,138,0,71,0,221,0,173,0,243,0,0,0,209,0,11,0,205,0,244,0,120,0,162,0,24,0,94,0,249,0,53,0,0,0,0,0,99,0,103,0,205,0,114,0,213,0,45,0,137,0,36,0,171,0,185,0,0,0,0,0,80,0,238,0,15,0,208,0,14,0,190,0,81,0,26,0,92,0,173,0,75,0,16,0,92,0,237,0,0,0,193,0,0,0,4,0,201,0,65,0,201,0,58,0,39,0,0,0,233,0,126,0,0,0,10,0,109,0,205,0,118,0,0,0,0,0,79,0,178,0,154,0,17,0,0,0,143,0,196,0,48,0,168,0,70,0,0,0,21,0,0,0,137,0,146,0,48,0,111,0,14,0,108,0,186,0,234,0,128,0,88,0,158,0,0,0,0,0,119,0,155,0,89,0,6,0,91,0,128,0,109,0,0,0,190,0,54,0,203,0,253,0,179,0,162,0,0,0,220,0,119,0,159,0,0,0,103,0,60,0,73,0,183,0,252,0,59,0,45,0,37,0,19,0,117,0,95,0,77,0,98,0,0,0,43,0,10,0,135,0,150,0,126,0,112,0,9,0,214,0,157,0,247,0,80,0,132,0,143,0,2,0,205,0,168,0,0,0,0,0,23,0,170,0,236,0,26,0,0,0,134,0,206,0,210,0,193,0,36,0,107,0,133,0,231,0,0,0,139,0,229,0,12,0,167,0,0,0,125,0,16,0,243,0,148,0,101,0,52,0,221,0,252,0,0,0,56,0,116,0,224,0,27,0,185,0,48,0,33,0,0,0,0,0,235,0,73,0,246,0,153,0,1,0,219,0,154,0,0,0,151,0,3,0,8,0,15,0,195,0,34,0,126,0,214,0,117,0,219,0,0,0,71,0,136,0,228,0,70,0,244,0,221,0,27,0,171,0,203,0,129,0,145,0,121,0,23,0,242,0,251,0,142,0,70,0,116,0,67,0,0,0,231,0,78,0,128,0,0,0,159,0,174,0,165,0,164,0,124,0,194,0,56,0,167,0,27,0,0,0,248,0,72,0,49,0,0,0,0,0,112,0,71,0,76,0,129,0,0,0,227,0,100,0,93,0,197,0,243,0,139,0,94,0,0,0,125,0,75,0,44,0,8,0,13,0,113,0,137,0,78,0,0,0,161,0,180,0,25,0,0,0,0,0,65,0,0,0,213,0,0,0,136,0,179,0,0,0,1,0,128,0,42,0,0,0,238,0,162,0,177,0,0,0,7,0,87,0,80,0,171,0,150,0,0,0,238,0,190,0,71,0,17,0,83,0,58,0,0,0,0,0,90,0,87,0,154,0,133,0,7,0,0,0,161,0,0,0,210,0,0,0,0,0,0,0,15,0,147,0,51,0,0,0,62,0,0,0,220,0,13,0);
signal scenario_full  : scenario_type := (168,31,91,31,132,31,191,31,191,30,191,29,91,31,86,31,150,31,187,31,107,31,75,31,3,31,17,31,168,31,184,31,50,31,155,31,53,31,159,31,81,31,149,31,55,31,55,30,131,31,119,31,119,30,32,31,32,30,239,31,204,31,147,31,3,31,208,31,160,31,254,31,184,31,13,31,13,30,116,31,90,31,247,31,247,30,203,31,203,30,203,29,167,31,97,31,228,31,212,31,95,31,95,30,95,29,197,31,63,31,63,30,129,31,129,30,103,31,88,31,126,31,134,31,61,31,191,31,249,31,65,31,57,31,255,31,190,31,57,31,216,31,18,31,94,31,94,30,252,31,32,31,149,31,17,31,168,31,65,31,217,31,239,31,239,30,177,31,102,31,202,31,87,31,87,30,87,29,166,31,233,31,176,31,38,31,58,31,58,30,114,31,68,31,189,31,36,31,104,31,244,31,86,31,210,31,111,31,84,31,188,31,29,31,73,31,217,31,155,31,116,31,209,31,228,31,228,30,119,31,146,31,183,31,50,31,50,30,166,31,166,30,95,31,95,30,8,31,208,31,173,31,231,31,138,31,71,31,221,31,173,31,243,31,243,30,209,31,11,31,205,31,244,31,120,31,162,31,24,31,94,31,249,31,53,31,53,30,53,29,99,31,103,31,205,31,114,31,213,31,45,31,137,31,36,31,171,31,185,31,185,30,185,29,80,31,238,31,15,31,208,31,14,31,190,31,81,31,26,31,92,31,173,31,75,31,16,31,92,31,237,31,237,30,193,31,193,30,4,31,201,31,65,31,201,31,58,31,39,31,39,30,233,31,126,31,126,30,10,31,109,31,205,31,118,31,118,30,118,29,79,31,178,31,154,31,17,31,17,30,143,31,196,31,48,31,168,31,70,31,70,30,21,31,21,30,137,31,146,31,48,31,111,31,14,31,108,31,186,31,234,31,128,31,88,31,158,31,158,30,158,29,119,31,155,31,89,31,6,31,91,31,128,31,109,31,109,30,190,31,54,31,203,31,253,31,179,31,162,31,162,30,220,31,119,31,159,31,159,30,103,31,60,31,73,31,183,31,252,31,59,31,45,31,37,31,19,31,117,31,95,31,77,31,98,31,98,30,43,31,10,31,135,31,150,31,126,31,112,31,9,31,214,31,157,31,247,31,80,31,132,31,143,31,2,31,205,31,168,31,168,30,168,29,23,31,170,31,236,31,26,31,26,30,134,31,206,31,210,31,193,31,36,31,107,31,133,31,231,31,231,30,139,31,229,31,12,31,167,31,167,30,125,31,16,31,243,31,148,31,101,31,52,31,221,31,252,31,252,30,56,31,116,31,224,31,27,31,185,31,48,31,33,31,33,30,33,29,235,31,73,31,246,31,153,31,1,31,219,31,154,31,154,30,151,31,3,31,8,31,15,31,195,31,34,31,126,31,214,31,117,31,219,31,219,30,71,31,136,31,228,31,70,31,244,31,221,31,27,31,171,31,203,31,129,31,145,31,121,31,23,31,242,31,251,31,142,31,70,31,116,31,67,31,67,30,231,31,78,31,128,31,128,30,159,31,174,31,165,31,164,31,124,31,194,31,56,31,167,31,27,31,27,30,248,31,72,31,49,31,49,30,49,29,112,31,71,31,76,31,129,31,129,30,227,31,100,31,93,31,197,31,243,31,139,31,94,31,94,30,125,31,75,31,44,31,8,31,13,31,113,31,137,31,78,31,78,30,161,31,180,31,25,31,25,30,25,29,65,31,65,30,213,31,213,30,136,31,179,31,179,30,1,31,128,31,42,31,42,30,238,31,162,31,177,31,177,30,7,31,87,31,80,31,171,31,150,31,150,30,238,31,190,31,71,31,17,31,83,31,58,31,58,30,58,29,90,31,87,31,154,31,133,31,7,31,7,30,161,31,161,30,210,31,210,30,210,29,210,28,15,31,147,31,51,31,51,30,62,31,62,30,220,31,13,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
