-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 685;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (239,0,66,0,0,0,244,0,64,0,110,0,78,0,178,0,0,0,81,0,220,0,160,0,0,0,40,0,22,0,200,0,211,0,40,0,1,0,0,0,117,0,88,0,174,0,0,0,17,0,143,0,209,0,90,0,132,0,131,0,178,0,76,0,216,0,35,0,15,0,241,0,189,0,164,0,0,0,2,0,62,0,245,0,90,0,139,0,166,0,184,0,169,0,45,0,80,0,0,0,190,0,14,0,0,0,0,0,240,0,144,0,213,0,201,0,0,0,100,0,0,0,74,0,150,0,0,0,0,0,129,0,0,0,150,0,0,0,80,0,66,0,16,0,20,0,121,0,131,0,122,0,0,0,129,0,0,0,125,0,0,0,239,0,144,0,0,0,122,0,0,0,173,0,244,0,0,0,110,0,39,0,15,0,213,0,140,0,110,0,179,0,158,0,247,0,117,0,0,0,215,0,129,0,103,0,134,0,114,0,0,0,25,0,138,0,0,0,237,0,68,0,0,0,139,0,220,0,110,0,82,0,0,0,121,0,0,0,61,0,0,0,115,0,247,0,216,0,250,0,144,0,92,0,0,0,188,0,16,0,255,0,222,0,132,0,228,0,138,0,159,0,9,0,224,0,174,0,240,0,0,0,15,0,119,0,24,0,99,0,188,0,245,0,180,0,113,0,167,0,89,0,220,0,238,0,41,0,141,0,50,0,32,0,249,0,0,0,0,0,104,0,95,0,172,0,130,0,119,0,0,0,22,0,234,0,230,0,49,0,105,0,67,0,50,0,13,0,40,0,12,0,0,0,65,0,15,0,23,0,17,0,74,0,199,0,0,0,0,0,221,0,242,0,119,0,70,0,55,0,1,0,44,0,54,0,90,0,206,0,82,0,205,0,138,0,0,0,111,0,0,0,9,0,229,0,47,0,0,0,50,0,129,0,0,0,17,0,0,0,0,0,74,0,205,0,0,0,51,0,189,0,188,0,0,0,133,0,0,0,178,0,205,0,207,0,102,0,46,0,0,0,165,0,0,0,192,0,17,0,152,0,144,0,129,0,60,0,173,0,135,0,149,0,101,0,0,0,30,0,178,0,0,0,28,0,56,0,245,0,219,0,39,0,173,0,137,0,0,0,0,0,0,0,214,0,115,0,128,0,228,0,0,0,0,0,48,0,208,0,0,0,191,0,113,0,76,0,192,0,17,0,53,0,116,0,44,0,161,0,65,0,0,0,234,0,102,0,11,0,228,0,0,0,32,0,45,0,104,0,162,0,46,0,237,0,86,0,156,0,124,0,147,0,233,0,184,0,0,0,216,0,254,0,182,0,0,0,60,0,91,0,220,0,194,0,130,0,132,0,38,0,223,0,220,0,97,0,53,0,107,0,0,0,118,0,5,0,184,0,238,0,162,0,158,0,144,0,0,0,133,0,36,0,150,0,159,0,109,0,243,0,147,0,0,0,143,0,130,0,117,0,58,0,0,0,27,0,0,0,177,0,236,0,243,0,62,0,109,0,119,0,19,0,0,0,0,0,237,0,29,0,29,0,75,0,143,0,173,0,46,0,0,0,112,0,149,0,250,0,42,0,108,0,125,0,220,0,0,0,239,0,83,0,0,0,179,0,0,0,253,0,0,0,145,0,154,0,7,0,242,0,17,0,0,0,186,0,242,0,107,0,0,0,0,0,196,0,25,0,0,0,37,0,238,0,130,0,121,0,68,0,0,0,228,0,167,0,33,0,247,0,183,0,232,0,199,0,0,0,216,0,132,0,86,0,81,0,0,0,250,0,136,0,33,0,127,0,58,0,243,0,0,0,181,0,7,0,15,0,152,0,0,0,30,0,139,0,60,0,126,0,135,0,75,0,0,0,93,0,209,0,0,0,0,0,175,0,189,0,88,0,106,0,195,0,21,0,44,0,203,0,78,0,47,0,195,0,140,0,12,0,98,0,76,0,116,0,109,0,0,0,141,0,47,0,0,0,0,0,74,0,4,0,0,0,0,0,0,0,128,0,0,0,243,0,197,0,119,0,218,0,202,0,0,0,0,0,138,0,109,0,0,0,0,0,0,0,0,0,33,0,208,0,154,0,79,0,134,0,36,0,20,0,0,0,0,0,0,0,0,0,0,0,11,0,227,0,195,0,154,0,132,0,0,0,92,0,72,0,37,0,176,0,85,0,128,0,99,0,161,0,45,0,175,0,31,0,212,0,124,0,243,0,0,0,150,0,187,0,2,0,234,0,14,0,0,0,76,0,219,0,51,0,160,0,0,0,0,0,201,0,0,0,126,0,0,0,239,0,0,0,0,0,74,0,125,0,226,0,0,0,189,0,123,0,43,0,195,0,65,0,174,0,206,0,232,0,64,0,0,0,0,0,0,0,232,0,214,0,29,0,83,0,228,0,173,0,76,0,141,0,159,0,140,0,189,0,3,0,3,0,183,0,3,0,74,0,246,0,35,0,169,0,174,0,0,0,101,0,38,0,254,0,30,0,221,0,209,0,125,0,36,0,133,0,0,0,217,0,0,0,0,0,248,0,122,0,2,0,153,0,56,0,204,0,0,0,245,0,118,0,7,0,143,0,187,0,0,0,0,0,237,0,7,0,108,0,132,0,153,0,48,0,118,0,119,0,54,0,230,0,254,0,246,0,0,0,35,0,61,0,15,0,0,0,152,0,209,0,139,0,251,0,0,0,0,0,14,0,230,0,67,0,28,0,22,0,6,0,63,0,53,0,217,0,145,0,249,0,242,0,98,0,172,0,48,0,133,0,209,0,138,0,0,0,92,0,0,0,196,0,20,0,0,0,55,0,165,0,0,0,0,0,173,0,176,0,67,0,0,0,0,0,0,0,191,0,219,0,75,0,12,0,7,0,0,0,198,0,0,0,31,0,41,0,0,0,198,0,51,0,188,0,1,0,138,0,67,0,196,0,26,0,0,0,0,0,220,0,198,0,12,0,90,0,30,0,0,0,0,0,45,0,88,0,162,0,0,0,241,0,36,0,217,0,6,0,228,0,251,0,145,0,97,0,32,0,157,0,195,0,139,0,62,0,254,0,0,0,47,0,78,0,20,0,6,0,70,0);
signal scenario_full  : scenario_type := (239,31,66,31,66,30,244,31,64,31,110,31,78,31,178,31,178,30,81,31,220,31,160,31,160,30,40,31,22,31,200,31,211,31,40,31,1,31,1,30,117,31,88,31,174,31,174,30,17,31,143,31,209,31,90,31,132,31,131,31,178,31,76,31,216,31,35,31,15,31,241,31,189,31,164,31,164,30,2,31,62,31,245,31,90,31,139,31,166,31,184,31,169,31,45,31,80,31,80,30,190,31,14,31,14,30,14,29,240,31,144,31,213,31,201,31,201,30,100,31,100,30,74,31,150,31,150,30,150,29,129,31,129,30,150,31,150,30,80,31,66,31,16,31,20,31,121,31,131,31,122,31,122,30,129,31,129,30,125,31,125,30,239,31,144,31,144,30,122,31,122,30,173,31,244,31,244,30,110,31,39,31,15,31,213,31,140,31,110,31,179,31,158,31,247,31,117,31,117,30,215,31,129,31,103,31,134,31,114,31,114,30,25,31,138,31,138,30,237,31,68,31,68,30,139,31,220,31,110,31,82,31,82,30,121,31,121,30,61,31,61,30,115,31,247,31,216,31,250,31,144,31,92,31,92,30,188,31,16,31,255,31,222,31,132,31,228,31,138,31,159,31,9,31,224,31,174,31,240,31,240,30,15,31,119,31,24,31,99,31,188,31,245,31,180,31,113,31,167,31,89,31,220,31,238,31,41,31,141,31,50,31,32,31,249,31,249,30,249,29,104,31,95,31,172,31,130,31,119,31,119,30,22,31,234,31,230,31,49,31,105,31,67,31,50,31,13,31,40,31,12,31,12,30,65,31,15,31,23,31,17,31,74,31,199,31,199,30,199,29,221,31,242,31,119,31,70,31,55,31,1,31,44,31,54,31,90,31,206,31,82,31,205,31,138,31,138,30,111,31,111,30,9,31,229,31,47,31,47,30,50,31,129,31,129,30,17,31,17,30,17,29,74,31,205,31,205,30,51,31,189,31,188,31,188,30,133,31,133,30,178,31,205,31,207,31,102,31,46,31,46,30,165,31,165,30,192,31,17,31,152,31,144,31,129,31,60,31,173,31,135,31,149,31,101,31,101,30,30,31,178,31,178,30,28,31,56,31,245,31,219,31,39,31,173,31,137,31,137,30,137,29,137,28,214,31,115,31,128,31,228,31,228,30,228,29,48,31,208,31,208,30,191,31,113,31,76,31,192,31,17,31,53,31,116,31,44,31,161,31,65,31,65,30,234,31,102,31,11,31,228,31,228,30,32,31,45,31,104,31,162,31,46,31,237,31,86,31,156,31,124,31,147,31,233,31,184,31,184,30,216,31,254,31,182,31,182,30,60,31,91,31,220,31,194,31,130,31,132,31,38,31,223,31,220,31,97,31,53,31,107,31,107,30,118,31,5,31,184,31,238,31,162,31,158,31,144,31,144,30,133,31,36,31,150,31,159,31,109,31,243,31,147,31,147,30,143,31,130,31,117,31,58,31,58,30,27,31,27,30,177,31,236,31,243,31,62,31,109,31,119,31,19,31,19,30,19,29,237,31,29,31,29,31,75,31,143,31,173,31,46,31,46,30,112,31,149,31,250,31,42,31,108,31,125,31,220,31,220,30,239,31,83,31,83,30,179,31,179,30,253,31,253,30,145,31,154,31,7,31,242,31,17,31,17,30,186,31,242,31,107,31,107,30,107,29,196,31,25,31,25,30,37,31,238,31,130,31,121,31,68,31,68,30,228,31,167,31,33,31,247,31,183,31,232,31,199,31,199,30,216,31,132,31,86,31,81,31,81,30,250,31,136,31,33,31,127,31,58,31,243,31,243,30,181,31,7,31,15,31,152,31,152,30,30,31,139,31,60,31,126,31,135,31,75,31,75,30,93,31,209,31,209,30,209,29,175,31,189,31,88,31,106,31,195,31,21,31,44,31,203,31,78,31,47,31,195,31,140,31,12,31,98,31,76,31,116,31,109,31,109,30,141,31,47,31,47,30,47,29,74,31,4,31,4,30,4,29,4,28,128,31,128,30,243,31,197,31,119,31,218,31,202,31,202,30,202,29,138,31,109,31,109,30,109,29,109,28,109,27,33,31,208,31,154,31,79,31,134,31,36,31,20,31,20,30,20,29,20,28,20,27,20,26,11,31,227,31,195,31,154,31,132,31,132,30,92,31,72,31,37,31,176,31,85,31,128,31,99,31,161,31,45,31,175,31,31,31,212,31,124,31,243,31,243,30,150,31,187,31,2,31,234,31,14,31,14,30,76,31,219,31,51,31,160,31,160,30,160,29,201,31,201,30,126,31,126,30,239,31,239,30,239,29,74,31,125,31,226,31,226,30,189,31,123,31,43,31,195,31,65,31,174,31,206,31,232,31,64,31,64,30,64,29,64,28,232,31,214,31,29,31,83,31,228,31,173,31,76,31,141,31,159,31,140,31,189,31,3,31,3,31,183,31,3,31,74,31,246,31,35,31,169,31,174,31,174,30,101,31,38,31,254,31,30,31,221,31,209,31,125,31,36,31,133,31,133,30,217,31,217,30,217,29,248,31,122,31,2,31,153,31,56,31,204,31,204,30,245,31,118,31,7,31,143,31,187,31,187,30,187,29,237,31,7,31,108,31,132,31,153,31,48,31,118,31,119,31,54,31,230,31,254,31,246,31,246,30,35,31,61,31,15,31,15,30,152,31,209,31,139,31,251,31,251,30,251,29,14,31,230,31,67,31,28,31,22,31,6,31,63,31,53,31,217,31,145,31,249,31,242,31,98,31,172,31,48,31,133,31,209,31,138,31,138,30,92,31,92,30,196,31,20,31,20,30,55,31,165,31,165,30,165,29,173,31,176,31,67,31,67,30,67,29,67,28,191,31,219,31,75,31,12,31,7,31,7,30,198,31,198,30,31,31,41,31,41,30,198,31,51,31,188,31,1,31,138,31,67,31,196,31,26,31,26,30,26,29,220,31,198,31,12,31,90,31,30,31,30,30,30,29,45,31,88,31,162,31,162,30,241,31,36,31,217,31,6,31,228,31,251,31,145,31,97,31,32,31,157,31,195,31,139,31,62,31,254,31,254,30,47,31,78,31,20,31,6,31,70,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
