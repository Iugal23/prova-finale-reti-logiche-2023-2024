-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_531 is
end project_tb_531;

architecture project_tb_arch_531 of project_tb_531 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 803;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (22,0,184,0,120,0,233,0,0,0,2,0,0,0,219,0,40,0,99,0,204,0,64,0,140,0,212,0,210,0,0,0,22,0,104,0,50,0,0,0,228,0,0,0,72,0,209,0,194,0,109,0,243,0,0,0,72,0,169,0,1,0,0,0,246,0,11,0,29,0,244,0,143,0,139,0,0,0,95,0,162,0,178,0,154,0,30,0,140,0,88,0,0,0,199,0,5,0,169,0,162,0,233,0,92,0,19,0,193,0,0,0,89,0,234,0,244,0,68,0,13,0,0,0,251,0,0,0,165,0,196,0,231,0,63,0,72,0,19,0,243,0,215,0,189,0,56,0,133,0,255,0,240,0,64,0,95,0,85,0,155,0,0,0,16,0,0,0,160,0,238,0,109,0,124,0,80,0,24,0,253,0,185,0,42,0,246,0,0,0,251,0,36,0,219,0,0,0,137,0,52,0,0,0,229,0,165,0,21,0,0,0,98,0,134,0,227,0,235,0,134,0,63,0,39,0,96,0,91,0,0,0,109,0,0,0,0,0,102,0,97,0,252,0,114,0,48,0,0,0,231,0,50,0,43,0,0,0,181,0,39,0,101,0,18,0,182,0,108,0,190,0,21,0,0,0,55,0,249,0,182,0,68,0,150,0,178,0,0,0,41,0,0,0,210,0,0,0,36,0,217,0,0,0,197,0,224,0,207,0,66,0,108,0,0,0,0,0,0,0,61,0,80,0,0,0,39,0,0,0,0,0,0,0,0,0,165,0,113,0,117,0,119,0,203,0,38,0,0,0,186,0,236,0,190,0,35,0,0,0,2,0,129,0,245,0,117,0,193,0,229,0,133,0,217,0,26,0,151,0,22,0,155,0,25,0,172,0,103,0,229,0,71,0,116,0,197,0,47,0,114,0,151,0,58,0,92,0,0,0,53,0,115,0,240,0,191,0,249,0,130,0,0,0,199,0,7,0,34,0,29,0,0,0,209,0,248,0,6,0,255,0,0,0,78,0,0,0,218,0,0,0,229,0,209,0,6,0,247,0,73,0,81,0,10,0,196,0,189,0,221,0,0,0,154,0,46,0,0,0,1,0,45,0,36,0,194,0,238,0,141,0,137,0,21,0,254,0,98,0,133,0,234,0,2,0,215,0,12,0,136,0,254,0,208,0,101,0,178,0,44,0,183,0,195,0,24,0,198,0,133,0,188,0,246,0,93,0,90,0,0,0,149,0,76,0,100,0,135,0,122,0,0,0,2,0,35,0,107,0,0,0,54,0,113,0,0,0,161,0,106,0,33,0,93,0,238,0,15,0,26,0,193,0,61,0,41,0,186,0,0,0,78,0,8,0,211,0,130,0,208,0,0,0,0,0,184,0,114,0,23,0,0,0,15,0,182,0,135,0,68,0,182,0,194,0,255,0,9,0,0,0,158,0,0,0,0,0,0,0,27,0,0,0,198,0,141,0,171,0,0,0,131,0,238,0,234,0,37,0,251,0,207,0,0,0,165,0,0,0,9,0,254,0,121,0,0,0,239,0,10,0,173,0,176,0,160,0,218,0,254,0,138,0,98,0,0,0,157,0,206,0,0,0,0,0,95,0,102,0,98,0,139,0,90,0,27,0,249,0,171,0,133,0,22,0,0,0,69,0,0,0,95,0,58,0,13,0,58,0,58,0,39,0,63,0,2,0,20,0,128,0,47,0,193,0,26,0,105,0,117,0,105,0,168,0,49,0,151,0,70,0,181,0,31,0,219,0,129,0,248,0,121,0,74,0,0,0,186,0,4,0,0,0,225,0,205,0,184,0,229,0,0,0,60,0,171,0,220,0,247,0,39,0,199,0,184,0,173,0,0,0,6,0,0,0,0,0,203,0,134,0,60,0,141,0,0,0,0,0,86,0,4,0,103,0,254,0,135,0,197,0,1,0,0,0,222,0,1,0,0,0,5,0,147,0,253,0,128,0,128,0,5,0,244,0,0,0,100,0,0,0,135,0,0,0,0,0,77,0,0,0,0,0,37,0,25,0,155,0,97,0,57,0,88,0,0,0,74,0,55,0,156,0,161,0,174,0,0,0,54,0,216,0,118,0,247,0,212,0,164,0,205,0,240,0,133,0,50,0,22,0,14,0,0,0,0,0,224,0,99,0,220,0,65,0,189,0,74,0,163,0,83,0,207,0,142,0,161,0,6,0,32,0,122,0,60,0,195,0,85,0,95,0,119,0,205,0,222,0,0,0,212,0,0,0,242,0,0,0,214,0,240,0,0,0,165,0,135,0,171,0,152,0,166,0,9,0,155,0,0,0,0,0,248,0,185,0,34,0,51,0,45,0,0,0,169,0,0,0,0,0,173,0,72,0,165,0,95,0,54,0,0,0,166,0,152,0,107,0,187,0,0,0,0,0,55,0,79,0,0,0,0,0,103,0,169,0,62,0,112,0,0,0,205,0,188,0,159,0,172,0,36,0,0,0,0,0,0,0,73,0,132,0,62,0,20,0,66,0,82,0,0,0,107,0,195,0,0,0,237,0,18,0,230,0,16,0,92,0,87,0,82,0,217,0,213,0,78,0,0,0,206,0,213,0,23,0,111,0,160,0,0,0,143,0,135,0,243,0,105,0,0,0,239,0,57,0,33,0,175,0,64,0,0,0,36,0,243,0,2,0,137,0,0,0,117,0,108,0,9,0,171,0,149,0,125,0,90,0,0,0,97,0,0,0,3,0,75,0,202,0,161,0,105,0,0,0,107,0,6,0,0,0,50,0,0,0,0,0,196,0,0,0,226,0,176,0,161,0,26,0,0,0,0,0,0,0,0,0,38,0,20,0,238,0,0,0,67,0,155,0,162,0,83,0,117,0,0,0,5,0,56,0,113,0,154,0,76,0,36,0,113,0,225,0,118,0,9,0,225,0,185,0,0,0,0,0,0,0,104,0,52,0,90,0,0,0,0,0,17,0,229,0,0,0,145,0,227,0,72,0,0,0,0,0,11,0,0,0,255,0,172,0,155,0,240,0,255,0,196,0,118,0,226,0,201,0,133,0,0,0,0,0,35,0,232,0,206,0,166,0,59,0,106,0,117,0,231,0,224,0,0,0,124,0,241,0,212,0,226,0,33,0,103,0,241,0,158,0,64,0,19,0,158,0,193,0,159,0,161,0,147,0,11,0,118,0,59,0,240,0,109,0,0,0,72,0,155,0,214,0,0,0,0,0,248,0,162,0,16,0,92,0,27,0,141,0,164,0,0,0,192,0,0,0,134,0,0,0,111,0,71,0,212,0,109,0,188,0,17,0,56,0,202,0,0,0,0,0,180,0,190,0,32,0,118,0,35,0,145,0,0,0,17,0,45,0,175,0,111,0,137,0,241,0,207,0,134,0,0,0,74,0,86,0,50,0,45,0,161,0,0,0,106,0,220,0,83,0,92,0,190,0,184,0,48,0,71,0,227,0,57,0,25,0,86,0,59,0,99,0,0,0,47,0,59,0,116,0,108,0,66,0,64,0,0,0,147,0,0,0,27,0,97,0,0,0,230,0,0,0,70,0,223,0,207,0,250,0,146,0,170,0,0,0,62,0,0,0,223,0,0,0,0,0,18,0,0,0,78,0,0,0,0,0);
signal scenario_full  : scenario_type := (22,31,184,31,120,31,233,31,233,30,2,31,2,30,219,31,40,31,99,31,204,31,64,31,140,31,212,31,210,31,210,30,22,31,104,31,50,31,50,30,228,31,228,30,72,31,209,31,194,31,109,31,243,31,243,30,72,31,169,31,1,31,1,30,246,31,11,31,29,31,244,31,143,31,139,31,139,30,95,31,162,31,178,31,154,31,30,31,140,31,88,31,88,30,199,31,5,31,169,31,162,31,233,31,92,31,19,31,193,31,193,30,89,31,234,31,244,31,68,31,13,31,13,30,251,31,251,30,165,31,196,31,231,31,63,31,72,31,19,31,243,31,215,31,189,31,56,31,133,31,255,31,240,31,64,31,95,31,85,31,155,31,155,30,16,31,16,30,160,31,238,31,109,31,124,31,80,31,24,31,253,31,185,31,42,31,246,31,246,30,251,31,36,31,219,31,219,30,137,31,52,31,52,30,229,31,165,31,21,31,21,30,98,31,134,31,227,31,235,31,134,31,63,31,39,31,96,31,91,31,91,30,109,31,109,30,109,29,102,31,97,31,252,31,114,31,48,31,48,30,231,31,50,31,43,31,43,30,181,31,39,31,101,31,18,31,182,31,108,31,190,31,21,31,21,30,55,31,249,31,182,31,68,31,150,31,178,31,178,30,41,31,41,30,210,31,210,30,36,31,217,31,217,30,197,31,224,31,207,31,66,31,108,31,108,30,108,29,108,28,61,31,80,31,80,30,39,31,39,30,39,29,39,28,39,27,165,31,113,31,117,31,119,31,203,31,38,31,38,30,186,31,236,31,190,31,35,31,35,30,2,31,129,31,245,31,117,31,193,31,229,31,133,31,217,31,26,31,151,31,22,31,155,31,25,31,172,31,103,31,229,31,71,31,116,31,197,31,47,31,114,31,151,31,58,31,92,31,92,30,53,31,115,31,240,31,191,31,249,31,130,31,130,30,199,31,7,31,34,31,29,31,29,30,209,31,248,31,6,31,255,31,255,30,78,31,78,30,218,31,218,30,229,31,209,31,6,31,247,31,73,31,81,31,10,31,196,31,189,31,221,31,221,30,154,31,46,31,46,30,1,31,45,31,36,31,194,31,238,31,141,31,137,31,21,31,254,31,98,31,133,31,234,31,2,31,215,31,12,31,136,31,254,31,208,31,101,31,178,31,44,31,183,31,195,31,24,31,198,31,133,31,188,31,246,31,93,31,90,31,90,30,149,31,76,31,100,31,135,31,122,31,122,30,2,31,35,31,107,31,107,30,54,31,113,31,113,30,161,31,106,31,33,31,93,31,238,31,15,31,26,31,193,31,61,31,41,31,186,31,186,30,78,31,8,31,211,31,130,31,208,31,208,30,208,29,184,31,114,31,23,31,23,30,15,31,182,31,135,31,68,31,182,31,194,31,255,31,9,31,9,30,158,31,158,30,158,29,158,28,27,31,27,30,198,31,141,31,171,31,171,30,131,31,238,31,234,31,37,31,251,31,207,31,207,30,165,31,165,30,9,31,254,31,121,31,121,30,239,31,10,31,173,31,176,31,160,31,218,31,254,31,138,31,98,31,98,30,157,31,206,31,206,30,206,29,95,31,102,31,98,31,139,31,90,31,27,31,249,31,171,31,133,31,22,31,22,30,69,31,69,30,95,31,58,31,13,31,58,31,58,31,39,31,63,31,2,31,20,31,128,31,47,31,193,31,26,31,105,31,117,31,105,31,168,31,49,31,151,31,70,31,181,31,31,31,219,31,129,31,248,31,121,31,74,31,74,30,186,31,4,31,4,30,225,31,205,31,184,31,229,31,229,30,60,31,171,31,220,31,247,31,39,31,199,31,184,31,173,31,173,30,6,31,6,30,6,29,203,31,134,31,60,31,141,31,141,30,141,29,86,31,4,31,103,31,254,31,135,31,197,31,1,31,1,30,222,31,1,31,1,30,5,31,147,31,253,31,128,31,128,31,5,31,244,31,244,30,100,31,100,30,135,31,135,30,135,29,77,31,77,30,77,29,37,31,25,31,155,31,97,31,57,31,88,31,88,30,74,31,55,31,156,31,161,31,174,31,174,30,54,31,216,31,118,31,247,31,212,31,164,31,205,31,240,31,133,31,50,31,22,31,14,31,14,30,14,29,224,31,99,31,220,31,65,31,189,31,74,31,163,31,83,31,207,31,142,31,161,31,6,31,32,31,122,31,60,31,195,31,85,31,95,31,119,31,205,31,222,31,222,30,212,31,212,30,242,31,242,30,214,31,240,31,240,30,165,31,135,31,171,31,152,31,166,31,9,31,155,31,155,30,155,29,248,31,185,31,34,31,51,31,45,31,45,30,169,31,169,30,169,29,173,31,72,31,165,31,95,31,54,31,54,30,166,31,152,31,107,31,187,31,187,30,187,29,55,31,79,31,79,30,79,29,103,31,169,31,62,31,112,31,112,30,205,31,188,31,159,31,172,31,36,31,36,30,36,29,36,28,73,31,132,31,62,31,20,31,66,31,82,31,82,30,107,31,195,31,195,30,237,31,18,31,230,31,16,31,92,31,87,31,82,31,217,31,213,31,78,31,78,30,206,31,213,31,23,31,111,31,160,31,160,30,143,31,135,31,243,31,105,31,105,30,239,31,57,31,33,31,175,31,64,31,64,30,36,31,243,31,2,31,137,31,137,30,117,31,108,31,9,31,171,31,149,31,125,31,90,31,90,30,97,31,97,30,3,31,75,31,202,31,161,31,105,31,105,30,107,31,6,31,6,30,50,31,50,30,50,29,196,31,196,30,226,31,176,31,161,31,26,31,26,30,26,29,26,28,26,27,38,31,20,31,238,31,238,30,67,31,155,31,162,31,83,31,117,31,117,30,5,31,56,31,113,31,154,31,76,31,36,31,113,31,225,31,118,31,9,31,225,31,185,31,185,30,185,29,185,28,104,31,52,31,90,31,90,30,90,29,17,31,229,31,229,30,145,31,227,31,72,31,72,30,72,29,11,31,11,30,255,31,172,31,155,31,240,31,255,31,196,31,118,31,226,31,201,31,133,31,133,30,133,29,35,31,232,31,206,31,166,31,59,31,106,31,117,31,231,31,224,31,224,30,124,31,241,31,212,31,226,31,33,31,103,31,241,31,158,31,64,31,19,31,158,31,193,31,159,31,161,31,147,31,11,31,118,31,59,31,240,31,109,31,109,30,72,31,155,31,214,31,214,30,214,29,248,31,162,31,16,31,92,31,27,31,141,31,164,31,164,30,192,31,192,30,134,31,134,30,111,31,71,31,212,31,109,31,188,31,17,31,56,31,202,31,202,30,202,29,180,31,190,31,32,31,118,31,35,31,145,31,145,30,17,31,45,31,175,31,111,31,137,31,241,31,207,31,134,31,134,30,74,31,86,31,50,31,45,31,161,31,161,30,106,31,220,31,83,31,92,31,190,31,184,31,48,31,71,31,227,31,57,31,25,31,86,31,59,31,99,31,99,30,47,31,59,31,116,31,108,31,66,31,64,31,64,30,147,31,147,30,27,31,97,31,97,30,230,31,230,30,70,31,223,31,207,31,250,31,146,31,170,31,170,30,62,31,62,30,223,31,223,30,223,29,18,31,18,30,78,31,78,30,78,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
