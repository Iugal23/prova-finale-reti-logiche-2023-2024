-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 326;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (192,0,14,0,0,0,114,0,0,0,0,0,215,0,83,0,76,0,219,0,0,0,0,0,0,0,0,0,148,0,208,0,252,0,111,0,66,0,227,0,0,0,230,0,0,0,64,0,0,0,79,0,255,0,0,0,9,0,117,0,222,0,0,0,97,0,0,0,0,0,44,0,173,0,120,0,0,0,1,0,140,0,109,0,100,0,188,0,194,0,130,0,37,0,236,0,0,0,0,0,232,0,90,0,123,0,133,0,0,0,97,0,253,0,239,0,57,0,161,0,91,0,68,0,108,0,0,0,74,0,0,0,21,0,0,0,0,0,239,0,3,0,166,0,0,0,220,0,90,0,0,0,138,0,42,0,0,0,0,0,0,0,150,0,34,0,0,0,126,0,0,0,0,0,234,0,183,0,0,0,94,0,219,0,251,0,0,0,196,0,187,0,222,0,183,0,234,0,0,0,6,0,6,0,119,0,117,0,174,0,184,0,231,0,244,0,211,0,250,0,0,0,207,0,142,0,159,0,0,0,70,0,0,0,116,0,209,0,159,0,21,0,158,0,58,0,0,0,210,0,106,0,54,0,226,0,216,0,236,0,126,0,24,0,123,0,0,0,151,0,238,0,77,0,107,0,12,0,14,0,0,0,158,0,55,0,28,0,115,0,138,0,0,0,86,0,0,0,5,0,130,0,74,0,94,0,0,0,115,0,0,0,232,0,114,0,192,0,200,0,0,0,48,0,0,0,6,0,198,0,93,0,207,0,230,0,86,0,208,0,171,0,0,0,0,0,226,0,0,0,0,0,77,0,116,0,95,0,24,0,244,0,16,0,0,0,4,0,0,0,132,0,0,0,245,0,0,0,240,0,0,0,180,0,229,0,22,0,50,0,0,0,1,0,80,0,253,0,0,0,0,0,69,0,107,0,143,0,100,0,209,0,0,0,83,0,245,0,67,0,130,0,168,0,190,0,0,0,0,0,24,0,0,0,0,0,1,0,189,0,179,0,122,0,66,0,0,0,28,0,1,0,69,0,13,0,0,0,207,0,0,0,56,0,138,0,0,0,207,0,2,0,87,0,123,0,55,0,241,0,46,0,75,0,27,0,1,0,253,0,202,0,80,0,72,0,100,0,174,0,79,0,108,0,0,0,13,0,50,0,246,0,103,0,133,0,71,0,41,0,166,0,207,0,193,0,0,0,130,0,48,0,186,0,15,0,222,0,205,0,90,0,110,0,0,0,196,0,198,0,210,0,0,0,0,0,246,0,169,0,102,0,0,0,50,0,242,0,142,0,158,0,152,0,77,0,92,0,6,0,52,0,40,0,26,0,41,0,18,0,0,0,182,0,178,0,218,0,229,0,198,0,0,0,138,0,174,0,0,0,56,0,235,0,219,0,45,0,118,0,224,0,51,0,210,0,99,0,0,0,87,0,0,0,0,0,198,0,231,0,0,0,115,0,122,0,25,0,0,0,71,0);
signal scenario_full  : scenario_type := (192,31,14,31,14,30,114,31,114,30,114,29,215,31,83,31,76,31,219,31,219,30,219,29,219,28,219,27,148,31,208,31,252,31,111,31,66,31,227,31,227,30,230,31,230,30,64,31,64,30,79,31,255,31,255,30,9,31,117,31,222,31,222,30,97,31,97,30,97,29,44,31,173,31,120,31,120,30,1,31,140,31,109,31,100,31,188,31,194,31,130,31,37,31,236,31,236,30,236,29,232,31,90,31,123,31,133,31,133,30,97,31,253,31,239,31,57,31,161,31,91,31,68,31,108,31,108,30,74,31,74,30,21,31,21,30,21,29,239,31,3,31,166,31,166,30,220,31,90,31,90,30,138,31,42,31,42,30,42,29,42,28,150,31,34,31,34,30,126,31,126,30,126,29,234,31,183,31,183,30,94,31,219,31,251,31,251,30,196,31,187,31,222,31,183,31,234,31,234,30,6,31,6,31,119,31,117,31,174,31,184,31,231,31,244,31,211,31,250,31,250,30,207,31,142,31,159,31,159,30,70,31,70,30,116,31,209,31,159,31,21,31,158,31,58,31,58,30,210,31,106,31,54,31,226,31,216,31,236,31,126,31,24,31,123,31,123,30,151,31,238,31,77,31,107,31,12,31,14,31,14,30,158,31,55,31,28,31,115,31,138,31,138,30,86,31,86,30,5,31,130,31,74,31,94,31,94,30,115,31,115,30,232,31,114,31,192,31,200,31,200,30,48,31,48,30,6,31,198,31,93,31,207,31,230,31,86,31,208,31,171,31,171,30,171,29,226,31,226,30,226,29,77,31,116,31,95,31,24,31,244,31,16,31,16,30,4,31,4,30,132,31,132,30,245,31,245,30,240,31,240,30,180,31,229,31,22,31,50,31,50,30,1,31,80,31,253,31,253,30,253,29,69,31,107,31,143,31,100,31,209,31,209,30,83,31,245,31,67,31,130,31,168,31,190,31,190,30,190,29,24,31,24,30,24,29,1,31,189,31,179,31,122,31,66,31,66,30,28,31,1,31,69,31,13,31,13,30,207,31,207,30,56,31,138,31,138,30,207,31,2,31,87,31,123,31,55,31,241,31,46,31,75,31,27,31,1,31,253,31,202,31,80,31,72,31,100,31,174,31,79,31,108,31,108,30,13,31,50,31,246,31,103,31,133,31,71,31,41,31,166,31,207,31,193,31,193,30,130,31,48,31,186,31,15,31,222,31,205,31,90,31,110,31,110,30,196,31,198,31,210,31,210,30,210,29,246,31,169,31,102,31,102,30,50,31,242,31,142,31,158,31,152,31,77,31,92,31,6,31,52,31,40,31,26,31,41,31,18,31,18,30,182,31,178,31,218,31,229,31,198,31,198,30,138,31,174,31,174,30,56,31,235,31,219,31,45,31,118,31,224,31,51,31,210,31,99,31,99,30,87,31,87,30,87,29,198,31,231,31,231,30,115,31,122,31,25,31,25,30,71,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
