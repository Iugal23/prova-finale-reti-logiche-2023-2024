-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_968 is
end project_tb_968;

architecture project_tb_arch_968 of project_tb_968 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 652;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (91,0,227,0,0,0,255,0,0,0,95,0,208,0,0,0,0,0,155,0,232,0,19,0,70,0,66,0,18,0,97,0,0,0,57,0,78,0,99,0,201,0,133,0,217,0,95,0,104,0,0,0,194,0,183,0,208,0,221,0,0,0,63,0,80,0,13,0,10,0,192,0,115,0,136,0,44,0,9,0,243,0,160,0,230,0,53,0,0,0,87,0,115,0,102,0,134,0,0,0,53,0,0,0,246,0,203,0,216,0,194,0,76,0,41,0,194,0,0,0,55,0,133,0,94,0,130,0,227,0,240,0,0,0,68,0,106,0,133,0,96,0,169,0,107,0,145,0,122,0,0,0,201,0,114,0,76,0,218,0,123,0,26,0,188,0,106,0,144,0,185,0,59,0,242,0,40,0,122,0,115,0,238,0,184,0,167,0,38,0,88,0,244,0,71,0,20,0,0,0,96,0,0,0,72,0,186,0,162,0,0,0,152,0,64,0,229,0,53,0,117,0,31,0,183,0,208,0,138,0,0,0,100,0,128,0,121,0,29,0,30,0,71,0,0,0,152,0,154,0,15,0,58,0,60,0,108,0,72,0,0,0,0,0,0,0,179,0,81,0,180,0,106,0,86,0,139,0,46,0,40,0,96,0,0,0,0,0,124,0,0,0,134,0,197,0,160,0,75,0,0,0,0,0,0,0,220,0,83,0,159,0,238,0,0,0,47,0,10,0,48,0,39,0,0,0,211,0,203,0,111,0,44,0,211,0,9,0,151,0,29,0,11,0,229,0,114,0,109,0,96,0,130,0,0,0,210,0,131,0,182,0,219,0,197,0,252,0,0,0,75,0,35,0,5,0,102,0,238,0,192,0,203,0,29,0,0,0,149,0,152,0,104,0,0,0,0,0,45,0,0,0,103,0,12,0,0,0,152,0,253,0,196,0,161,0,0,0,223,0,176,0,87,0,106,0,221,0,97,0,192,0,158,0,61,0,89,0,27,0,0,0,226,0,183,0,0,0,151,0,0,0,0,0,206,0,55,0,166,0,55,0,206,0,132,0,82,0,0,0,78,0,156,0,196,0,0,0,151,0,132,0,34,0,0,0,31,0,120,0,0,0,0,0,41,0,143,0,244,0,0,0,68,0,0,0,254,0,13,0,137,0,0,0,206,0,179,0,61,0,249,0,203,0,192,0,0,0,252,0,0,0,125,0,155,0,191,0,117,0,252,0,232,0,151,0,165,0,190,0,0,0,0,0,0,0,0,0,55,0,122,0,2,0,0,0,214,0,138,0,95,0,0,0,234,0,251,0,239,0,247,0,47,0,0,0,62,0,153,0,170,0,180,0,29,0,0,0,137,0,251,0,251,0,119,0,0,0,75,0,152,0,0,0,0,0,108,0,0,0,143,0,0,0,90,0,14,0,207,0,96,0,11,0,153,0,215,0,87,0,248,0,199,0,203,0,202,0,113,0,228,0,98,0,19,0,190,0,137,0,2,0,0,0,160,0,75,0,142,0,0,0,107,0,249,0,86,0,169,0,4,0,142,0,188,0,34,0,147,0,158,0,65,0,237,0,0,0,196,0,0,0,36,0,222,0,175,0,236,0,0,0,232,0,37,0,215,0,79,0,226,0,10,0,0,0,148,0,226,0,0,0,218,0,36,0,202,0,116,0,34,0,107,0,160,0,0,0,0,0,103,0,89,0,207,0,242,0,63,0,243,0,96,0,12,0,31,0,36,0,24,0,0,0,203,0,36,0,0,0,0,0,0,0,133,0,86,0,24,0,0,0,164,0,226,0,16,0,13,0,57,0,12,0,158,0,0,0,4,0,0,0,0,0,5,0,136,0,82,0,0,0,68,0,135,0,22,0,254,0,117,0,35,0,107,0,146,0,171,0,0,0,219,0,152,0,0,0,215,0,15,0,168,0,93,0,21,0,134,0,0,0,0,0,219,0,0,0,106,0,65,0,150,0,0,0,0,0,0,0,207,0,0,0,207,0,122,0,0,0,213,0,0,0,0,0,81,0,3,0,0,0,165,0,56,0,172,0,96,0,0,0,0,0,136,0,149,0,0,0,181,0,220,0,136,0,83,0,229,0,142,0,0,0,0,0,132,0,78,0,209,0,36,0,68,0,131,0,159,0,0,0,150,0,176,0,49,0,148,0,28,0,133,0,70,0,218,0,0,0,164,0,0,0,251,0,79,0,10,0,33,0,192,0,81,0,252,0,164,0,253,0,223,0,203,0,97,0,111,0,208,0,15,0,64,0,66,0,59,0,152,0,40,0,119,0,0,0,172,0,54,0,51,0,68,0,85,0,243,0,34,0,179,0,188,0,15,0,107,0,164,0,20,0,130,0,1,0,161,0,133,0,0,0,48,0,21,0,0,0,90,0,200,0,138,0,168,0,13,0,39,0,78,0,0,0,238,0,132,0,33,0,193,0,9,0,90,0,216,0,0,0,212,0,54,0,183,0,198,0,0,0,232,0,0,0,0,0,27,0,0,0,0,0,177,0,129,0,146,0,103,0,203,0,70,0,0,0,140,0,45,0,0,0,163,0,46,0,110,0,0,0,251,0,34,0,0,0,92,0,254,0,20,0,164,0,69,0,83,0,105,0,0,0,109,0,0,0,77,0,24,0,0,0,73,0,37,0,227,0,210,0,39,0,0,0,73,0,106,0,54,0,0,0,91,0,0,0,3,0,139,0,234,0,178,0,0,0,0,0,126,0,82,0,117,0,0,0,154,0,162,0,35,0,255,0,73,0,199,0,22,0,46,0,110,0,74,0,225,0,87,0,16,0,20,0,192,0,25,0,224,0,236,0,95,0,172,0,117,0,240,0,255,0,123,0,208,0,229,0,123,0,197,0,120,0,168,0,245,0,0,0,8,0,159,0,241,0,210,0,0,0,148,0,174,0,0,0,211,0,1,0,97,0);
signal scenario_full  : scenario_type := (91,31,227,31,227,30,255,31,255,30,95,31,208,31,208,30,208,29,155,31,232,31,19,31,70,31,66,31,18,31,97,31,97,30,57,31,78,31,99,31,201,31,133,31,217,31,95,31,104,31,104,30,194,31,183,31,208,31,221,31,221,30,63,31,80,31,13,31,10,31,192,31,115,31,136,31,44,31,9,31,243,31,160,31,230,31,53,31,53,30,87,31,115,31,102,31,134,31,134,30,53,31,53,30,246,31,203,31,216,31,194,31,76,31,41,31,194,31,194,30,55,31,133,31,94,31,130,31,227,31,240,31,240,30,68,31,106,31,133,31,96,31,169,31,107,31,145,31,122,31,122,30,201,31,114,31,76,31,218,31,123,31,26,31,188,31,106,31,144,31,185,31,59,31,242,31,40,31,122,31,115,31,238,31,184,31,167,31,38,31,88,31,244,31,71,31,20,31,20,30,96,31,96,30,72,31,186,31,162,31,162,30,152,31,64,31,229,31,53,31,117,31,31,31,183,31,208,31,138,31,138,30,100,31,128,31,121,31,29,31,30,31,71,31,71,30,152,31,154,31,15,31,58,31,60,31,108,31,72,31,72,30,72,29,72,28,179,31,81,31,180,31,106,31,86,31,139,31,46,31,40,31,96,31,96,30,96,29,124,31,124,30,134,31,197,31,160,31,75,31,75,30,75,29,75,28,220,31,83,31,159,31,238,31,238,30,47,31,10,31,48,31,39,31,39,30,211,31,203,31,111,31,44,31,211,31,9,31,151,31,29,31,11,31,229,31,114,31,109,31,96,31,130,31,130,30,210,31,131,31,182,31,219,31,197,31,252,31,252,30,75,31,35,31,5,31,102,31,238,31,192,31,203,31,29,31,29,30,149,31,152,31,104,31,104,30,104,29,45,31,45,30,103,31,12,31,12,30,152,31,253,31,196,31,161,31,161,30,223,31,176,31,87,31,106,31,221,31,97,31,192,31,158,31,61,31,89,31,27,31,27,30,226,31,183,31,183,30,151,31,151,30,151,29,206,31,55,31,166,31,55,31,206,31,132,31,82,31,82,30,78,31,156,31,196,31,196,30,151,31,132,31,34,31,34,30,31,31,120,31,120,30,120,29,41,31,143,31,244,31,244,30,68,31,68,30,254,31,13,31,137,31,137,30,206,31,179,31,61,31,249,31,203,31,192,31,192,30,252,31,252,30,125,31,155,31,191,31,117,31,252,31,232,31,151,31,165,31,190,31,190,30,190,29,190,28,190,27,55,31,122,31,2,31,2,30,214,31,138,31,95,31,95,30,234,31,251,31,239,31,247,31,47,31,47,30,62,31,153,31,170,31,180,31,29,31,29,30,137,31,251,31,251,31,119,31,119,30,75,31,152,31,152,30,152,29,108,31,108,30,143,31,143,30,90,31,14,31,207,31,96,31,11,31,153,31,215,31,87,31,248,31,199,31,203,31,202,31,113,31,228,31,98,31,19,31,190,31,137,31,2,31,2,30,160,31,75,31,142,31,142,30,107,31,249,31,86,31,169,31,4,31,142,31,188,31,34,31,147,31,158,31,65,31,237,31,237,30,196,31,196,30,36,31,222,31,175,31,236,31,236,30,232,31,37,31,215,31,79,31,226,31,10,31,10,30,148,31,226,31,226,30,218,31,36,31,202,31,116,31,34,31,107,31,160,31,160,30,160,29,103,31,89,31,207,31,242,31,63,31,243,31,96,31,12,31,31,31,36,31,24,31,24,30,203,31,36,31,36,30,36,29,36,28,133,31,86,31,24,31,24,30,164,31,226,31,16,31,13,31,57,31,12,31,158,31,158,30,4,31,4,30,4,29,5,31,136,31,82,31,82,30,68,31,135,31,22,31,254,31,117,31,35,31,107,31,146,31,171,31,171,30,219,31,152,31,152,30,215,31,15,31,168,31,93,31,21,31,134,31,134,30,134,29,219,31,219,30,106,31,65,31,150,31,150,30,150,29,150,28,207,31,207,30,207,31,122,31,122,30,213,31,213,30,213,29,81,31,3,31,3,30,165,31,56,31,172,31,96,31,96,30,96,29,136,31,149,31,149,30,181,31,220,31,136,31,83,31,229,31,142,31,142,30,142,29,132,31,78,31,209,31,36,31,68,31,131,31,159,31,159,30,150,31,176,31,49,31,148,31,28,31,133,31,70,31,218,31,218,30,164,31,164,30,251,31,79,31,10,31,33,31,192,31,81,31,252,31,164,31,253,31,223,31,203,31,97,31,111,31,208,31,15,31,64,31,66,31,59,31,152,31,40,31,119,31,119,30,172,31,54,31,51,31,68,31,85,31,243,31,34,31,179,31,188,31,15,31,107,31,164,31,20,31,130,31,1,31,161,31,133,31,133,30,48,31,21,31,21,30,90,31,200,31,138,31,168,31,13,31,39,31,78,31,78,30,238,31,132,31,33,31,193,31,9,31,90,31,216,31,216,30,212,31,54,31,183,31,198,31,198,30,232,31,232,30,232,29,27,31,27,30,27,29,177,31,129,31,146,31,103,31,203,31,70,31,70,30,140,31,45,31,45,30,163,31,46,31,110,31,110,30,251,31,34,31,34,30,92,31,254,31,20,31,164,31,69,31,83,31,105,31,105,30,109,31,109,30,77,31,24,31,24,30,73,31,37,31,227,31,210,31,39,31,39,30,73,31,106,31,54,31,54,30,91,31,91,30,3,31,139,31,234,31,178,31,178,30,178,29,126,31,82,31,117,31,117,30,154,31,162,31,35,31,255,31,73,31,199,31,22,31,46,31,110,31,74,31,225,31,87,31,16,31,20,31,192,31,25,31,224,31,236,31,95,31,172,31,117,31,240,31,255,31,123,31,208,31,229,31,123,31,197,31,120,31,168,31,245,31,245,30,8,31,159,31,241,31,210,31,210,30,148,31,174,31,174,30,211,31,1,31,97,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
