-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 957;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,93,0,158,0,221,0,40,0,104,0,114,0,153,0,0,0,167,0,132,0,159,0,141,0,219,0,100,0,100,0,1,0,0,0,3,0,127,0,195,0,115,0,130,0,108,0,43,0,141,0,0,0,197,0,46,0,150,0,0,0,183,0,121,0,246,0,6,0,35,0,137,0,0,0,44,0,82,0,183,0,157,0,7,0,66,0,128,0,93,0,71,0,0,0,172,0,43,0,38,0,225,0,45,0,212,0,22,0,69,0,43,0,54,0,118,0,199,0,29,0,109,0,0,0,228,0,225,0,0,0,0,0,151,0,0,0,210,0,181,0,202,0,186,0,131,0,113,0,85,0,9,0,238,0,34,0,159,0,101,0,4,0,244,0,103,0,167,0,0,0,0,0,180,0,113,0,35,0,7,0,246,0,220,0,0,0,94,0,227,0,0,0,82,0,0,0,161,0,59,0,0,0,5,0,56,0,149,0,226,0,90,0,74,0,139,0,151,0,0,0,0,0,0,0,227,0,50,0,228,0,27,0,104,0,244,0,164,0,191,0,116,0,246,0,22,0,48,0,61,0,229,0,101,0,200,0,0,0,252,0,0,0,0,0,221,0,157,0,215,0,30,0,28,0,253,0,111,0,173,0,0,0,182,0,94,0,245,0,148,0,194,0,231,0,123,0,246,0,140,0,0,0,149,0,199,0,11,0,49,0,116,0,122,0,21,0,247,0,0,0,242,0,52,0,226,0,88,0,223,0,0,0,159,0,0,0,97,0,0,0,179,0,55,0,49,0,179,0,2,0,0,0,65,0,46,0,0,0,105,0,7,0,0,0,144,0,119,0,0,0,221,0,104,0,230,0,86,0,0,0,156,0,0,0,120,0,93,0,228,0,0,0,0,0,92,0,64,0,81,0,128,0,75,0,237,0,237,0,107,0,73,0,160,0,135,0,0,0,193,0,0,0,146,0,165,0,229,0,189,0,0,0,164,0,18,0,37,0,0,0,19,0,0,0,183,0,157,0,163,0,152,0,202,0,237,0,0,0,67,0,200,0,42,0,100,0,92,0,63,0,165,0,202,0,132,0,0,0,0,0,193,0,98,0,32,0,214,0,242,0,0,0,22,0,91,0,0,0,0,0,0,0,0,0,0,0,165,0,129,0,217,0,54,0,6,0,50,0,178,0,37,0,79,0,147,0,123,0,163,0,84,0,0,0,0,0,83,0,5,0,241,0,228,0,91,0,153,0,154,0,75,0,47,0,104,0,68,0,37,0,121,0,234,0,183,0,0,0,113,0,143,0,38,0,39,0,0,0,222,0,156,0,188,0,40,0,211,0,160,0,97,0,177,0,61,0,131,0,76,0,240,0,49,0,47,0,4,0,170,0,0,0,238,0,76,0,179,0,0,0,10,0,77,0,131,0,108,0,0,0,15,0,255,0,109,0,0,0,185,0,165,0,26,0,128,0,4,0,232,0,0,0,211,0,185,0,197,0,0,0,0,0,92,0,166,0,50,0,0,0,251,0,206,0,0,0,60,0,0,0,0,0,66,0,188,0,0,0,13,0,148,0,173,0,172,0,179,0,68,0,73,0,52,0,0,0,241,0,229,0,21,0,139,0,231,0,0,0,89,0,229,0,133,0,87,0,82,0,69,0,0,0,183,0,222,0,0,0,99,0,72,0,0,0,94,0,251,0,200,0,139,0,42,0,34,0,185,0,41,0,162,0,208,0,0,0,0,0,2,0,0,0,0,0,242,0,195,0,16,0,98,0,182,0,0,0,9,0,83,0,26,0,187,0,167,0,13,0,78,0,118,0,91,0,244,0,220,0,70,0,170,0,185,0,43,0,0,0,224,0,144,0,0,0,124,0,0,0,175,0,126,0,30,0,221,0,7,0,93,0,29,0,0,0,26,0,0,0,105,0,79,0,15,0,10,0,103,0,0,0,92,0,149,0,108,0,174,0,0,0,75,0,136,0,148,0,90,0,20,0,46,0,0,0,239,0,182,0,169,0,0,0,91,0,235,0,179,0,95,0,127,0,81,0,224,0,150,0,64,0,0,0,203,0,243,0,0,0,0,0,0,0,154,0,202,0,130,0,252,0,52,0,0,0,0,0,1,0,0,0,53,0,2,0,41,0,12,0,27,0,52,0,11,0,144,0,0,0,0,0,136,0,0,0,15,0,47,0,31,0,111,0,250,0,215,0,14,0,0,0,93,0,28,0,10,0,42,0,16,0,100,0,220,0,232,0,147,0,48,0,0,0,0,0,65,0,1,0,73,0,143,0,0,0,10,0,147,0,83,0,183,0,0,0,200,0,186,0,182,0,95,0,152,0,0,0,171,0,35,0,93,0,0,0,183,0,104,0,0,0,66,0,138,0,137,0,143,0,198,0,167,0,152,0,0,0,245,0,186,0,124,0,234,0,0,0,42,0,0,0,203,0,251,0,0,0,26,0,0,0,58,0,115,0,0,0,192,0,202,0,119,0,137,0,185,0,143,0,0,0,238,0,0,0,1,0,19,0,229,0,78,0,60,0,0,0,0,0,0,0,22,0,16,0,215,0,151,0,2,0,214,0,0,0,0,0,0,0,68,0,234,0,0,0,2,0,0,0,45,0,0,0,34,0,19,0,90,0,206,0,46,0,132,0,213,0,31,0,174,0,0,0,0,0,208,0,44,0,237,0,81,0,220,0,141,0,5,0,42,0,182,0,193,0,119,0,113,0,24,0,216,0,86,0,181,0,45,0,197,0,0,0,104,0,181,0,235,0,201,0,132,0,0,0,0,0,17,0,184,0,70,0,155,0,183,0,204,0,35,0,240,0,142,0,56,0,39,0,124,0,101,0,224,0,146,0,248,0,12,0,0,0,212,0,192,0,108,0,152,0,78,0,66,0,62,0,0,0,136,0,250,0,173,0,223,0,182,0,0,0,148,0,104,0,209,0,0,0,0,0,215,0,162,0,76,0,88,0,0,0,8,0,218,0,173,0,0,0,133,0,190,0,183,0,36,0,0,0,85,0,231,0,0,0,13,0,0,0,24,0,155,0,200,0,0,0,59,0,178,0,237,0,227,0,0,0,38,0,0,0,113,0,0,0,231,0,17,0,168,0,98,0,141,0,228,0,165,0,36,0,0,0,178,0,178,0,94,0,0,0,48,0,0,0,117,0,120,0,0,0,158,0,0,0,251,0,9,0,243,0,0,0,239,0,83,0,146,0,135,0,82,0,230,0,163,0,151,0,246,0,49,0,0,0,59,0,154,0,157,0,0,0,145,0,0,0,0,0,0,0,11,0,125,0,194,0,172,0,0,0,44,0,133,0,9,0,64,0,159,0,31,0,159,0,249,0,0,0,15,0,0,0,67,0,161,0,0,0,0,0,169,0,74,0,228,0,144,0,4,0,3,0,224,0,0,0,51,0,35,0,88,0,0,0,191,0,184,0,100,0,64,0,63,0,122,0,69,0,199,0,0,0,0,0,71,0,60,0,30,0,220,0,57,0,51,0,227,0,28,0,97,0,47,0,0,0,0,0,214,0,128,0,0,0,22,0,102,0,0,0,145,0,0,0,106,0,170,0,144,0,194,0,211,0,188,0,168,0,34,0,238,0,43,0,248,0,0,0,151,0,180,0,217,0,23,0,114,0,216,0,15,0,47,0,219,0,70,0,9,0,228,0,28,0,168,0,167,0,0,0,57,0,239,0,200,0,0,0,0,0,181,0,52,0,146,0,91,0,72,0,194,0,237,0,39,0,0,0,185,0,190,0,0,0,46,0,18,0,250,0,146,0,0,0,0,0,220,0,244,0,0,0,215,0,0,0,61,0,0,0,77,0,62,0,249,0,72,0,0,0,136,0,56,0,0,0,94,0,46,0,147,0,87,0,0,0,157,0,126,0,0,0,25,0,118,0,99,0,0,0,0,0,201,0,194,0,0,0,125,0,194,0,252,0,165,0,75,0,178,0,151,0,0,0,80,0,87,0,216,0,0,0,247,0,0,0,135,0,238,0,130,0,69,0,166,0,29,0,107,0,0,0,4,0,237,0,59,0,43,0,0,0,224,0,212,0,14,0,173,0,19,0,185,0,48,0,78,0,241,0,145,0,169,0,49,0,0,0,156,0,0,0,228,0,61,0,57,0,249,0,142,0,117,0,0,0,219,0,0,0,65,0,48,0,63,0,0,0,65,0,2,0,248,0,28,0,149,0,246,0,184,0,81,0,251,0,78,0,185,0,56,0,0,0,43,0,142,0,0,0,130,0,116,0,200,0,41,0,147,0,91,0,105,0,118,0,168,0,0,0,207,0);
signal scenario_full  : scenario_type := (0,0,93,31,158,31,221,31,40,31,104,31,114,31,153,31,153,30,167,31,132,31,159,31,141,31,219,31,100,31,100,31,1,31,1,30,3,31,127,31,195,31,115,31,130,31,108,31,43,31,141,31,141,30,197,31,46,31,150,31,150,30,183,31,121,31,246,31,6,31,35,31,137,31,137,30,44,31,82,31,183,31,157,31,7,31,66,31,128,31,93,31,71,31,71,30,172,31,43,31,38,31,225,31,45,31,212,31,22,31,69,31,43,31,54,31,118,31,199,31,29,31,109,31,109,30,228,31,225,31,225,30,225,29,151,31,151,30,210,31,181,31,202,31,186,31,131,31,113,31,85,31,9,31,238,31,34,31,159,31,101,31,4,31,244,31,103,31,167,31,167,30,167,29,180,31,113,31,35,31,7,31,246,31,220,31,220,30,94,31,227,31,227,30,82,31,82,30,161,31,59,31,59,30,5,31,56,31,149,31,226,31,90,31,74,31,139,31,151,31,151,30,151,29,151,28,227,31,50,31,228,31,27,31,104,31,244,31,164,31,191,31,116,31,246,31,22,31,48,31,61,31,229,31,101,31,200,31,200,30,252,31,252,30,252,29,221,31,157,31,215,31,30,31,28,31,253,31,111,31,173,31,173,30,182,31,94,31,245,31,148,31,194,31,231,31,123,31,246,31,140,31,140,30,149,31,199,31,11,31,49,31,116,31,122,31,21,31,247,31,247,30,242,31,52,31,226,31,88,31,223,31,223,30,159,31,159,30,97,31,97,30,179,31,55,31,49,31,179,31,2,31,2,30,65,31,46,31,46,30,105,31,7,31,7,30,144,31,119,31,119,30,221,31,104,31,230,31,86,31,86,30,156,31,156,30,120,31,93,31,228,31,228,30,228,29,92,31,64,31,81,31,128,31,75,31,237,31,237,31,107,31,73,31,160,31,135,31,135,30,193,31,193,30,146,31,165,31,229,31,189,31,189,30,164,31,18,31,37,31,37,30,19,31,19,30,183,31,157,31,163,31,152,31,202,31,237,31,237,30,67,31,200,31,42,31,100,31,92,31,63,31,165,31,202,31,132,31,132,30,132,29,193,31,98,31,32,31,214,31,242,31,242,30,22,31,91,31,91,30,91,29,91,28,91,27,91,26,165,31,129,31,217,31,54,31,6,31,50,31,178,31,37,31,79,31,147,31,123,31,163,31,84,31,84,30,84,29,83,31,5,31,241,31,228,31,91,31,153,31,154,31,75,31,47,31,104,31,68,31,37,31,121,31,234,31,183,31,183,30,113,31,143,31,38,31,39,31,39,30,222,31,156,31,188,31,40,31,211,31,160,31,97,31,177,31,61,31,131,31,76,31,240,31,49,31,47,31,4,31,170,31,170,30,238,31,76,31,179,31,179,30,10,31,77,31,131,31,108,31,108,30,15,31,255,31,109,31,109,30,185,31,165,31,26,31,128,31,4,31,232,31,232,30,211,31,185,31,197,31,197,30,197,29,92,31,166,31,50,31,50,30,251,31,206,31,206,30,60,31,60,30,60,29,66,31,188,31,188,30,13,31,148,31,173,31,172,31,179,31,68,31,73,31,52,31,52,30,241,31,229,31,21,31,139,31,231,31,231,30,89,31,229,31,133,31,87,31,82,31,69,31,69,30,183,31,222,31,222,30,99,31,72,31,72,30,94,31,251,31,200,31,139,31,42,31,34,31,185,31,41,31,162,31,208,31,208,30,208,29,2,31,2,30,2,29,242,31,195,31,16,31,98,31,182,31,182,30,9,31,83,31,26,31,187,31,167,31,13,31,78,31,118,31,91,31,244,31,220,31,70,31,170,31,185,31,43,31,43,30,224,31,144,31,144,30,124,31,124,30,175,31,126,31,30,31,221,31,7,31,93,31,29,31,29,30,26,31,26,30,105,31,79,31,15,31,10,31,103,31,103,30,92,31,149,31,108,31,174,31,174,30,75,31,136,31,148,31,90,31,20,31,46,31,46,30,239,31,182,31,169,31,169,30,91,31,235,31,179,31,95,31,127,31,81,31,224,31,150,31,64,31,64,30,203,31,243,31,243,30,243,29,243,28,154,31,202,31,130,31,252,31,52,31,52,30,52,29,1,31,1,30,53,31,2,31,41,31,12,31,27,31,52,31,11,31,144,31,144,30,144,29,136,31,136,30,15,31,47,31,31,31,111,31,250,31,215,31,14,31,14,30,93,31,28,31,10,31,42,31,16,31,100,31,220,31,232,31,147,31,48,31,48,30,48,29,65,31,1,31,73,31,143,31,143,30,10,31,147,31,83,31,183,31,183,30,200,31,186,31,182,31,95,31,152,31,152,30,171,31,35,31,93,31,93,30,183,31,104,31,104,30,66,31,138,31,137,31,143,31,198,31,167,31,152,31,152,30,245,31,186,31,124,31,234,31,234,30,42,31,42,30,203,31,251,31,251,30,26,31,26,30,58,31,115,31,115,30,192,31,202,31,119,31,137,31,185,31,143,31,143,30,238,31,238,30,1,31,19,31,229,31,78,31,60,31,60,30,60,29,60,28,22,31,16,31,215,31,151,31,2,31,214,31,214,30,214,29,214,28,68,31,234,31,234,30,2,31,2,30,45,31,45,30,34,31,19,31,90,31,206,31,46,31,132,31,213,31,31,31,174,31,174,30,174,29,208,31,44,31,237,31,81,31,220,31,141,31,5,31,42,31,182,31,193,31,119,31,113,31,24,31,216,31,86,31,181,31,45,31,197,31,197,30,104,31,181,31,235,31,201,31,132,31,132,30,132,29,17,31,184,31,70,31,155,31,183,31,204,31,35,31,240,31,142,31,56,31,39,31,124,31,101,31,224,31,146,31,248,31,12,31,12,30,212,31,192,31,108,31,152,31,78,31,66,31,62,31,62,30,136,31,250,31,173,31,223,31,182,31,182,30,148,31,104,31,209,31,209,30,209,29,215,31,162,31,76,31,88,31,88,30,8,31,218,31,173,31,173,30,133,31,190,31,183,31,36,31,36,30,85,31,231,31,231,30,13,31,13,30,24,31,155,31,200,31,200,30,59,31,178,31,237,31,227,31,227,30,38,31,38,30,113,31,113,30,231,31,17,31,168,31,98,31,141,31,228,31,165,31,36,31,36,30,178,31,178,31,94,31,94,30,48,31,48,30,117,31,120,31,120,30,158,31,158,30,251,31,9,31,243,31,243,30,239,31,83,31,146,31,135,31,82,31,230,31,163,31,151,31,246,31,49,31,49,30,59,31,154,31,157,31,157,30,145,31,145,30,145,29,145,28,11,31,125,31,194,31,172,31,172,30,44,31,133,31,9,31,64,31,159,31,31,31,159,31,249,31,249,30,15,31,15,30,67,31,161,31,161,30,161,29,169,31,74,31,228,31,144,31,4,31,3,31,224,31,224,30,51,31,35,31,88,31,88,30,191,31,184,31,100,31,64,31,63,31,122,31,69,31,199,31,199,30,199,29,71,31,60,31,30,31,220,31,57,31,51,31,227,31,28,31,97,31,47,31,47,30,47,29,214,31,128,31,128,30,22,31,102,31,102,30,145,31,145,30,106,31,170,31,144,31,194,31,211,31,188,31,168,31,34,31,238,31,43,31,248,31,248,30,151,31,180,31,217,31,23,31,114,31,216,31,15,31,47,31,219,31,70,31,9,31,228,31,28,31,168,31,167,31,167,30,57,31,239,31,200,31,200,30,200,29,181,31,52,31,146,31,91,31,72,31,194,31,237,31,39,31,39,30,185,31,190,31,190,30,46,31,18,31,250,31,146,31,146,30,146,29,220,31,244,31,244,30,215,31,215,30,61,31,61,30,77,31,62,31,249,31,72,31,72,30,136,31,56,31,56,30,94,31,46,31,147,31,87,31,87,30,157,31,126,31,126,30,25,31,118,31,99,31,99,30,99,29,201,31,194,31,194,30,125,31,194,31,252,31,165,31,75,31,178,31,151,31,151,30,80,31,87,31,216,31,216,30,247,31,247,30,135,31,238,31,130,31,69,31,166,31,29,31,107,31,107,30,4,31,237,31,59,31,43,31,43,30,224,31,212,31,14,31,173,31,19,31,185,31,48,31,78,31,241,31,145,31,169,31,49,31,49,30,156,31,156,30,228,31,61,31,57,31,249,31,142,31,117,31,117,30,219,31,219,30,65,31,48,31,63,31,63,30,65,31,2,31,248,31,28,31,149,31,246,31,184,31,81,31,251,31,78,31,185,31,56,31,56,30,43,31,142,31,142,30,130,31,116,31,200,31,41,31,147,31,91,31,105,31,118,31,168,31,168,30,207,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
