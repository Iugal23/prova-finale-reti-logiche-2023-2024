-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_200 is
end project_tb_200;

architecture project_tb_arch_200 of project_tb_200 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 531;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (247,0,142,0,106,0,0,0,0,0,62,0,66,0,230,0,165,0,184,0,182,0,59,0,94,0,180,0,0,0,0,0,201,0,7,0,73,0,43,0,55,0,183,0,106,0,0,0,0,0,150,0,44,0,187,0,223,0,0,0,19,0,234,0,214,0,194,0,55,0,32,0,160,0,242,0,213,0,0,0,0,0,180,0,0,0,14,0,246,0,129,0,0,0,147,0,0,0,0,0,113,0,78,0,25,0,143,0,0,0,34,0,159,0,31,0,60,0,245,0,96,0,190,0,40,0,14,0,38,0,136,0,0,0,146,0,227,0,187,0,85,0,0,0,197,0,152,0,56,0,229,0,0,0,0,0,220,0,169,0,127,0,152,0,46,0,7,0,216,0,19,0,26,0,0,0,48,0,49,0,0,0,251,0,2,0,98,0,240,0,6,0,155,0,208,0,129,0,102,0,65,0,142,0,187,0,10,0,203,0,137,0,221,0,77,0,152,0,55,0,99,0,144,0,5,0,147,0,147,0,0,0,67,0,117,0,122,0,0,0,211,0,224,0,139,0,0,0,55,0,133,0,0,0,85,0,0,0,129,0,99,0,178,0,35,0,206,0,0,0,254,0,225,0,199,0,120,0,0,0,80,0,241,0,3,0,16,0,0,0,75,0,207,0,138,0,3,0,72,0,195,0,154,0,212,0,92,0,245,0,0,0,24,0,235,0,144,0,207,0,249,0,12,0,69,0,56,0,146,0,73,0,218,0,0,0,22,0,0,0,163,0,8,0,0,0,146,0,100,0,0,0,90,0,222,0,0,0,0,0,0,0,0,0,178,0,0,0,142,0,65,0,0,0,0,0,0,0,245,0,255,0,0,0,0,0,0,0,69,0,195,0,160,0,138,0,0,0,54,0,0,0,10,0,19,0,94,0,0,0,102,0,38,0,0,0,77,0,64,0,182,0,32,0,0,0,236,0,223,0,22,0,56,0,0,0,37,0,0,0,24,0,94,0,115,0,97,0,104,0,151,0,0,0,138,0,152,0,17,0,138,0,212,0,133,0,125,0,47,0,58,0,155,0,231,0,25,0,166,0,215,0,247,0,20,0,205,0,0,0,186,0,26,0,0,0,0,0,183,0,220,0,44,0,96,0,0,0,0,0,0,0,99,0,223,0,113,0,178,0,98,0,40,0,253,0,237,0,104,0,0,0,78,0,57,0,79,0,81,0,126,0,45,0,248,0,7,0,169,0,210,0,148,0,47,0,130,0,245,0,136,0,44,0,234,0,0,0,163,0,197,0,39,0,102,0,0,0,0,0,150,0,95,0,171,0,37,0,66,0,164,0,189,0,213,0,101,0,141,0,133,0,167,0,67,0,155,0,0,0,188,0,195,0,42,0,221,0,0,0,61,0,0,0,0,0,124,0,32,0,149,0,0,0,4,0,0,0,0,0,160,0,0,0,15,0,3,0,116,0,0,0,0,0,58,0,0,0,123,0,202,0,140,0,233,0,37,0,44,0,9,0,135,0,0,0,227,0,0,0,92,0,0,0,0,0,195,0,0,0,125,0,16,0,87,0,103,0,149,0,0,0,0,0,0,0,0,0,127,0,91,0,162,0,0,0,6,0,246,0,95,0,181,0,0,0,129,0,121,0,121,0,221,0,88,0,244,0,0,0,0,0,201,0,0,0,249,0,101,0,0,0,0,0,211,0,71,0,225,0,136,0,0,0,91,0,148,0,109,0,0,0,106,0,183,0,0,0,0,0,116,0,183,0,0,0,220,0,155,0,129,0,125,0,156,0,242,0,198,0,0,0,253,0,27,0,0,0,190,0,69,0,176,0,4,0,196,0,57,0,0,0,42,0,201,0,201,0,0,0,188,0,80,0,139,0,0,0,159,0,0,0,148,0,94,0,175,0,0,0,190,0,0,0,0,0,48,0,103,0,186,0,141,0,64,0,1,0,20,0,194,0,103,0,148,0,0,0,0,0,133,0,112,0,75,0,5,0,9,0,0,0,185,0,31,0,229,0,0,0,164,0,0,0,0,0,0,0,169,0,0,0,139,0,74,0,76,0,33,0,115,0,101,0,51,0,0,0,93,0,222,0,165,0,188,0,81,0,0,0,68,0,35,0,0,0,177,0,0,0,151,0,78,0,192,0,0,0,196,0,174,0,226,0,247,0,133,0,157,0,108,0,79,0,14,0,171,0,0,0,0,0,35,0,147,0,71,0,59,0,185,0,214,0,98,0,41,0,0,0,0,0,0,0,182,0,60,0,171,0,134,0,94,0,144,0,68,0,15,0,0,0,207,0,98,0,170,0,0,0,64,0,194,0,207,0,117,0,192,0,88,0,83,0,159,0,225,0,0,0,0,0,169,0,176,0,111,0,71,0,215,0);
signal scenario_full  : scenario_type := (247,31,142,31,106,31,106,30,106,29,62,31,66,31,230,31,165,31,184,31,182,31,59,31,94,31,180,31,180,30,180,29,201,31,7,31,73,31,43,31,55,31,183,31,106,31,106,30,106,29,150,31,44,31,187,31,223,31,223,30,19,31,234,31,214,31,194,31,55,31,32,31,160,31,242,31,213,31,213,30,213,29,180,31,180,30,14,31,246,31,129,31,129,30,147,31,147,30,147,29,113,31,78,31,25,31,143,31,143,30,34,31,159,31,31,31,60,31,245,31,96,31,190,31,40,31,14,31,38,31,136,31,136,30,146,31,227,31,187,31,85,31,85,30,197,31,152,31,56,31,229,31,229,30,229,29,220,31,169,31,127,31,152,31,46,31,7,31,216,31,19,31,26,31,26,30,48,31,49,31,49,30,251,31,2,31,98,31,240,31,6,31,155,31,208,31,129,31,102,31,65,31,142,31,187,31,10,31,203,31,137,31,221,31,77,31,152,31,55,31,99,31,144,31,5,31,147,31,147,31,147,30,67,31,117,31,122,31,122,30,211,31,224,31,139,31,139,30,55,31,133,31,133,30,85,31,85,30,129,31,99,31,178,31,35,31,206,31,206,30,254,31,225,31,199,31,120,31,120,30,80,31,241,31,3,31,16,31,16,30,75,31,207,31,138,31,3,31,72,31,195,31,154,31,212,31,92,31,245,31,245,30,24,31,235,31,144,31,207,31,249,31,12,31,69,31,56,31,146,31,73,31,218,31,218,30,22,31,22,30,163,31,8,31,8,30,146,31,100,31,100,30,90,31,222,31,222,30,222,29,222,28,222,27,178,31,178,30,142,31,65,31,65,30,65,29,65,28,245,31,255,31,255,30,255,29,255,28,69,31,195,31,160,31,138,31,138,30,54,31,54,30,10,31,19,31,94,31,94,30,102,31,38,31,38,30,77,31,64,31,182,31,32,31,32,30,236,31,223,31,22,31,56,31,56,30,37,31,37,30,24,31,94,31,115,31,97,31,104,31,151,31,151,30,138,31,152,31,17,31,138,31,212,31,133,31,125,31,47,31,58,31,155,31,231,31,25,31,166,31,215,31,247,31,20,31,205,31,205,30,186,31,26,31,26,30,26,29,183,31,220,31,44,31,96,31,96,30,96,29,96,28,99,31,223,31,113,31,178,31,98,31,40,31,253,31,237,31,104,31,104,30,78,31,57,31,79,31,81,31,126,31,45,31,248,31,7,31,169,31,210,31,148,31,47,31,130,31,245,31,136,31,44,31,234,31,234,30,163,31,197,31,39,31,102,31,102,30,102,29,150,31,95,31,171,31,37,31,66,31,164,31,189,31,213,31,101,31,141,31,133,31,167,31,67,31,155,31,155,30,188,31,195,31,42,31,221,31,221,30,61,31,61,30,61,29,124,31,32,31,149,31,149,30,4,31,4,30,4,29,160,31,160,30,15,31,3,31,116,31,116,30,116,29,58,31,58,30,123,31,202,31,140,31,233,31,37,31,44,31,9,31,135,31,135,30,227,31,227,30,92,31,92,30,92,29,195,31,195,30,125,31,16,31,87,31,103,31,149,31,149,30,149,29,149,28,149,27,127,31,91,31,162,31,162,30,6,31,246,31,95,31,181,31,181,30,129,31,121,31,121,31,221,31,88,31,244,31,244,30,244,29,201,31,201,30,249,31,101,31,101,30,101,29,211,31,71,31,225,31,136,31,136,30,91,31,148,31,109,31,109,30,106,31,183,31,183,30,183,29,116,31,183,31,183,30,220,31,155,31,129,31,125,31,156,31,242,31,198,31,198,30,253,31,27,31,27,30,190,31,69,31,176,31,4,31,196,31,57,31,57,30,42,31,201,31,201,31,201,30,188,31,80,31,139,31,139,30,159,31,159,30,148,31,94,31,175,31,175,30,190,31,190,30,190,29,48,31,103,31,186,31,141,31,64,31,1,31,20,31,194,31,103,31,148,31,148,30,148,29,133,31,112,31,75,31,5,31,9,31,9,30,185,31,31,31,229,31,229,30,164,31,164,30,164,29,164,28,169,31,169,30,139,31,74,31,76,31,33,31,115,31,101,31,51,31,51,30,93,31,222,31,165,31,188,31,81,31,81,30,68,31,35,31,35,30,177,31,177,30,151,31,78,31,192,31,192,30,196,31,174,31,226,31,247,31,133,31,157,31,108,31,79,31,14,31,171,31,171,30,171,29,35,31,147,31,71,31,59,31,185,31,214,31,98,31,41,31,41,30,41,29,41,28,182,31,60,31,171,31,134,31,94,31,144,31,68,31,15,31,15,30,207,31,98,31,170,31,170,30,64,31,194,31,207,31,117,31,192,31,88,31,83,31,159,31,225,31,225,30,225,29,169,31,176,31,111,31,71,31,215,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
