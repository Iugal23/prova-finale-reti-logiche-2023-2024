-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_860 is
end project_tb_860;

architecture project_tb_arch_860 of project_tb_860 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 550;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (201,0,171,0,98,0,230,0,0,0,37,0,203,0,192,0,136,0,107,0,0,0,16,0,0,0,0,0,156,0,117,0,0,0,77,0,200,0,45,0,0,0,106,0,202,0,72,0,60,0,36,0,3,0,0,0,55,0,0,0,0,0,86,0,0,0,0,0,115,0,0,0,33,0,163,0,48,0,251,0,70,0,77,0,219,0,167,0,0,0,113,0,229,0,214,0,110,0,239,0,132,0,111,0,0,0,115,0,0,0,166,0,107,0,0,0,0,0,0,0,229,0,246,0,0,0,0,0,0,0,104,0,52,0,216,0,239,0,158,0,197,0,212,0,48,0,195,0,31,0,0,0,0,0,136,0,7,0,0,0,149,0,0,0,104,0,183,0,8,0,0,0,201,0,213,0,243,0,204,0,180,0,2,0,252,0,92,0,64,0,81,0,41,0,0,0,71,0,63,0,0,0,140,0,0,0,0,0,203,0,0,0,213,0,114,0,0,0,77,0,109,0,18,0,16,0,85,0,0,0,235,0,211,0,98,0,156,0,166,0,246,0,13,0,240,0,202,0,16,0,53,0,146,0,154,0,34,0,213,0,114,0,0,0,252,0,54,0,0,0,0,0,60,0,205,0,129,0,240,0,11,0,0,0,0,0,6,0,140,0,0,0,57,0,46,0,0,0,63,0,107,0,183,0,0,0,185,0,210,0,155,0,144,0,94,0,36,0,255,0,234,0,201,0,66,0,198,0,161,0,115,0,12,0,190,0,242,0,140,0,71,0,25,0,162,0,0,0,174,0,89,0,84,0,43,0,78,0,0,0,22,0,0,0,104,0,172,0,77,0,7,0,54,0,113,0,0,0,0,0,157,0,195,0,121,0,142,0,230,0,31,0,77,0,45,0,247,0,35,0,142,0,173,0,4,0,183,0,225,0,251,0,0,0,175,0,94,0,184,0,240,0,95,0,208,0,4,0,176,0,0,0,33,0,242,0,78,0,0,0,0,0,134,0,0,0,252,0,246,0,211,0,150,0,0,0,0,0,56,0,0,0,87,0,58,0,232,0,2,0,5,0,0,0,0,0,135,0,77,0,136,0,0,0,220,0,220,0,195,0,223,0,62,0,105,0,88,0,75,0,73,0,90,0,176,0,0,0,0,0,179,0,155,0,88,0,117,0,52,0,0,0,148,0,0,0,79,0,42,0,0,0,222,0,179,0,0,0,230,0,77,0,62,0,79,0,25,0,162,0,215,0,133,0,25,0,173,0,121,0,124,0,137,0,155,0,0,0,92,0,142,0,211,0,134,0,78,0,245,0,69,0,36,0,185,0,111,0,96,0,225,0,1,0,171,0,124,0,208,0,65,0,112,0,115,0,131,0,224,0,6,0,39,0,32,0,0,0,76,0,36,0,113,0,136,0,157,0,200,0,126,0,0,0,86,0,0,0,62,0,149,0,59,0,219,0,168,0,150,0,148,0,101,0,171,0,242,0,0,0,81,0,106,0,93,0,86,0,25,0,0,0,166,0,0,0,36,0,231,0,207,0,51,0,0,0,111,0,0,0,209,0,231,0,109,0,0,0,238,0,180,0,171,0,228,0,148,0,38,0,242,0,220,0,0,0,221,0,144,0,187,0,80,0,142,0,0,0,63,0,0,0,48,0,146,0,0,0,173,0,0,0,22,0,0,0,58,0,74,0,186,0,0,0,0,0,0,0,123,0,145,0,251,0,252,0,0,0,0,0,237,0,114,0,69,0,103,0,198,0,15,0,0,0,88,0,31,0,137,0,237,0,223,0,50,0,19,0,160,0,182,0,0,0,0,0,229,0,143,0,129,0,0,0,71,0,208,0,0,0,0,0,208,0,220,0,68,0,25,0,0,0,212,0,0,0,45,0,98,0,221,0,200,0,232,0,46,0,244,0,0,0,65,0,246,0,56,0,152,0,0,0,0,0,22,0,196,0,27,0,69,0,189,0,58,0,182,0,242,0,108,0,138,0,120,0,17,0,0,0,94,0,228,0,93,0,0,0,100,0,12,0,196,0,144,0,118,0,135,0,201,0,157,0,128,0,0,0,162,0,0,0,116,0,197,0,20,0,2,0,33,0,92,0,0,0,171,0,169,0,38,0,0,0,151,0,251,0,145,0,0,0,0,0,78,0,163,0,213,0,0,0,13,0,205,0,186,0,238,0,164,0,243,0,137,0,227,0,242,0,49,0,186,0,60,0,193,0,236,0,217,0,96,0,245,0,155,0,0,0,205,0,62,0,143,0,117,0,167,0,0,0,111,0,204,0,0,0,44,0,229,0,170,0,212,0,158,0,0,0,239,0,0,0,29,0,0,0,109,0,50,0,9,0,35,0,203,0,233,0,226,0,148,0,97,0,245,0,9,0,234,0,131,0,29,0,8,0,32,0,0,0,160,0,24,0,112,0,0,0,3,0,0,0,119,0,189,0,141,0,19,0,0,0,0,0,248,0,244,0);
signal scenario_full  : scenario_type := (201,31,171,31,98,31,230,31,230,30,37,31,203,31,192,31,136,31,107,31,107,30,16,31,16,30,16,29,156,31,117,31,117,30,77,31,200,31,45,31,45,30,106,31,202,31,72,31,60,31,36,31,3,31,3,30,55,31,55,30,55,29,86,31,86,30,86,29,115,31,115,30,33,31,163,31,48,31,251,31,70,31,77,31,219,31,167,31,167,30,113,31,229,31,214,31,110,31,239,31,132,31,111,31,111,30,115,31,115,30,166,31,107,31,107,30,107,29,107,28,229,31,246,31,246,30,246,29,246,28,104,31,52,31,216,31,239,31,158,31,197,31,212,31,48,31,195,31,31,31,31,30,31,29,136,31,7,31,7,30,149,31,149,30,104,31,183,31,8,31,8,30,201,31,213,31,243,31,204,31,180,31,2,31,252,31,92,31,64,31,81,31,41,31,41,30,71,31,63,31,63,30,140,31,140,30,140,29,203,31,203,30,213,31,114,31,114,30,77,31,109,31,18,31,16,31,85,31,85,30,235,31,211,31,98,31,156,31,166,31,246,31,13,31,240,31,202,31,16,31,53,31,146,31,154,31,34,31,213,31,114,31,114,30,252,31,54,31,54,30,54,29,60,31,205,31,129,31,240,31,11,31,11,30,11,29,6,31,140,31,140,30,57,31,46,31,46,30,63,31,107,31,183,31,183,30,185,31,210,31,155,31,144,31,94,31,36,31,255,31,234,31,201,31,66,31,198,31,161,31,115,31,12,31,190,31,242,31,140,31,71,31,25,31,162,31,162,30,174,31,89,31,84,31,43,31,78,31,78,30,22,31,22,30,104,31,172,31,77,31,7,31,54,31,113,31,113,30,113,29,157,31,195,31,121,31,142,31,230,31,31,31,77,31,45,31,247,31,35,31,142,31,173,31,4,31,183,31,225,31,251,31,251,30,175,31,94,31,184,31,240,31,95,31,208,31,4,31,176,31,176,30,33,31,242,31,78,31,78,30,78,29,134,31,134,30,252,31,246,31,211,31,150,31,150,30,150,29,56,31,56,30,87,31,58,31,232,31,2,31,5,31,5,30,5,29,135,31,77,31,136,31,136,30,220,31,220,31,195,31,223,31,62,31,105,31,88,31,75,31,73,31,90,31,176,31,176,30,176,29,179,31,155,31,88,31,117,31,52,31,52,30,148,31,148,30,79,31,42,31,42,30,222,31,179,31,179,30,230,31,77,31,62,31,79,31,25,31,162,31,215,31,133,31,25,31,173,31,121,31,124,31,137,31,155,31,155,30,92,31,142,31,211,31,134,31,78,31,245,31,69,31,36,31,185,31,111,31,96,31,225,31,1,31,171,31,124,31,208,31,65,31,112,31,115,31,131,31,224,31,6,31,39,31,32,31,32,30,76,31,36,31,113,31,136,31,157,31,200,31,126,31,126,30,86,31,86,30,62,31,149,31,59,31,219,31,168,31,150,31,148,31,101,31,171,31,242,31,242,30,81,31,106,31,93,31,86,31,25,31,25,30,166,31,166,30,36,31,231,31,207,31,51,31,51,30,111,31,111,30,209,31,231,31,109,31,109,30,238,31,180,31,171,31,228,31,148,31,38,31,242,31,220,31,220,30,221,31,144,31,187,31,80,31,142,31,142,30,63,31,63,30,48,31,146,31,146,30,173,31,173,30,22,31,22,30,58,31,74,31,186,31,186,30,186,29,186,28,123,31,145,31,251,31,252,31,252,30,252,29,237,31,114,31,69,31,103,31,198,31,15,31,15,30,88,31,31,31,137,31,237,31,223,31,50,31,19,31,160,31,182,31,182,30,182,29,229,31,143,31,129,31,129,30,71,31,208,31,208,30,208,29,208,31,220,31,68,31,25,31,25,30,212,31,212,30,45,31,98,31,221,31,200,31,232,31,46,31,244,31,244,30,65,31,246,31,56,31,152,31,152,30,152,29,22,31,196,31,27,31,69,31,189,31,58,31,182,31,242,31,108,31,138,31,120,31,17,31,17,30,94,31,228,31,93,31,93,30,100,31,12,31,196,31,144,31,118,31,135,31,201,31,157,31,128,31,128,30,162,31,162,30,116,31,197,31,20,31,2,31,33,31,92,31,92,30,171,31,169,31,38,31,38,30,151,31,251,31,145,31,145,30,145,29,78,31,163,31,213,31,213,30,13,31,205,31,186,31,238,31,164,31,243,31,137,31,227,31,242,31,49,31,186,31,60,31,193,31,236,31,217,31,96,31,245,31,155,31,155,30,205,31,62,31,143,31,117,31,167,31,167,30,111,31,204,31,204,30,44,31,229,31,170,31,212,31,158,31,158,30,239,31,239,30,29,31,29,30,109,31,50,31,9,31,35,31,203,31,233,31,226,31,148,31,97,31,245,31,9,31,234,31,131,31,29,31,8,31,32,31,32,30,160,31,24,31,112,31,112,30,3,31,3,30,119,31,189,31,141,31,19,31,19,30,19,29,248,31,244,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
