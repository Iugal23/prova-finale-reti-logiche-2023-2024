-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_524 is
end project_tb_524;

architecture project_tb_arch_524 of project_tb_524 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 679;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (254,0,0,0,0,0,210,0,0,0,99,0,102,0,107,0,38,0,104,0,223,0,185,0,0,0,243,0,252,0,139,0,177,0,174,0,95,0,215,0,161,0,214,0,164,0,0,0,241,0,0,0,53,0,184,0,102,0,158,0,0,0,143,0,186,0,185,0,136,0,165,0,0,0,70,0,130,0,169,0,47,0,59,0,77,0,120,0,0,0,176,0,9,0,140,0,14,0,102,0,146,0,65,0,63,0,0,0,98,0,0,0,0,0,0,0,122,0,112,0,177,0,0,0,64,0,42,0,87,0,180,0,80,0,105,0,153,0,51,0,219,0,45,0,0,0,158,0,15,0,252,0,176,0,70,0,4,0,254,0,0,0,7,0,251,0,197,0,241,0,31,0,0,0,217,0,126,0,39,0,28,0,12,0,162,0,5,0,15,0,76,0,3,0,91,0,0,0,0,0,219,0,40,0,0,0,0,0,239,0,49,0,0,0,146,0,224,0,155,0,126,0,0,0,133,0,107,0,111,0,26,0,1,0,169,0,46,0,8,0,141,0,55,0,201,0,0,0,87,0,60,0,117,0,157,0,0,0,184,0,160,0,79,0,155,0,87,0,27,0,216,0,13,0,151,0,239,0,94,0,160,0,154,0,212,0,0,0,149,0,221,0,15,0,137,0,185,0,0,0,242,0,21,0,0,0,23,0,224,0,250,0,162,0,146,0,100,0,123,0,116,0,66,0,12,0,215,0,245,0,4,0,229,0,194,0,189,0,70,0,202,0,94,0,113,0,172,0,0,0,244,0,16,0,71,0,222,0,169,0,0,0,38,0,55,0,84,0,136,0,68,0,36,0,79,0,0,0,161,0,6,0,30,0,85,0,0,0,201,0,215,0,116,0,0,0,232,0,33,0,149,0,102,0,23,0,0,0,218,0,128,0,51,0,148,0,196,0,58,0,65,0,32,0,183,0,206,0,201,0,1,0,0,0,192,0,34,0,0,0,168,0,253,0,162,0,0,0,90,0,198,0,0,0,244,0,129,0,11,0,118,0,0,0,76,0,0,0,0,0,142,0,14,0,0,0,211,0,0,0,179,0,11,0,139,0,208,0,39,0,157,0,142,0,176,0,212,0,130,0,0,0,49,0,119,0,0,0,58,0,234,0,0,0,0,0,0,0,163,0,162,0,44,0,173,0,54,0,156,0,0,0,204,0,172,0,52,0,15,0,93,0,77,0,13,0,253,0,176,0,0,0,131,0,26,0,120,0,220,0,212,0,0,0,0,0,225,0,85,0,9,0,120,0,77,0,113,0,181,0,234,0,0,0,124,0,0,0,237,0,132,0,165,0,4,0,250,0,0,0,243,0,8,0,180,0,0,0,230,0,221,0,65,0,0,0,239,0,240,0,183,0,152,0,208,0,168,0,166,0,8,0,17,0,75,0,89,0,86,0,173,0,0,0,0,0,0,0,95,0,168,0,64,0,158,0,255,0,38,0,28,0,26,0,6,0,42,0,139,0,188,0,202,0,233,0,69,0,0,0,100,0,0,0,77,0,5,0,10,0,0,0,0,0,182,0,0,0,0,0,179,0,124,0,252,0,41,0,79,0,0,0,201,0,98,0,141,0,175,0,140,0,187,0,151,0,0,0,121,0,232,0,133,0,106,0,203,0,146,0,40,0,168,0,138,0,12,0,133,0,108,0,119,0,0,0,195,0,0,0,137,0,98,0,0,0,100,0,0,0,241,0,202,0,218,0,135,0,3,0,0,0,224,0,210,0,43,0,78,0,0,0,137,0,0,0,0,0,1,0,224,0,70,0,139,0,97,0,155,0,246,0,0,0,0,0,79,0,151,0,0,0,0,0,124,0,0,0,235,0,161,0,96,0,76,0,132,0,74,0,0,0,0,0,78,0,129,0,0,0,55,0,201,0,88,0,0,0,188,0,44,0,194,0,97,0,157,0,162,0,97,0,0,0,0,0,106,0,140,0,54,0,0,0,133,0,159,0,245,0,115,0,241,0,200,0,172,0,5,0,0,0,152,0,165,0,87,0,161,0,157,0,62,0,235,0,69,0,0,0,116,0,88,0,50,0,0,0,85,0,0,0,83,0,0,0,7,0,244,0,26,0,0,0,172,0,170,0,83,0,0,0,0,0,191,0,32,0,154,0,125,0,126,0,0,0,16,0,0,0,183,0,0,0,12,0,182,0,194,0,174,0,222,0,52,0,20,0,171,0,71,0,154,0,227,0,88,0,107,0,106,0,0,0,248,0,156,0,195,0,164,0,0,0,37,0,0,0,240,0,72,0,130,0,250,0,0,0,236,0,134,0,240,0,10,0,129,0,131,0,0,0,19,0,202,0,50,0,249,0,97,0,1,0,205,0,42,0,0,0,213,0,0,0,27,0,0,0,82,0,189,0,166,0,118,0,242,0,239,0,127,0,46,0,194,0,175,0,27,0,9,0,56,0,24,0,30,0,0,0,104,0,176,0,99,0,0,0,23,0,0,0,31,0,88,0,181,0,57,0,185,0,0,0,97,0,220,0,209,0,222,0,161,0,77,0,138,0,119,0,32,0,239,0,197,0,131,0,0,0,30,0,0,0,196,0,0,0,90,0,164,0,17,0,107,0,254,0,117,0,94,0,226,0,248,0,12,0,213,0,92,0,38,0,0,0,142,0,0,0,0,0,230,0,215,0,161,0,42,0,139,0,221,0,232,0,0,0,0,0,106,0,0,0,109,0,128,0,188,0,4,0,236,0,0,0,213,0,253,0,159,0,224,0,0,0,53,0,135,0,151,0,238,0,126,0,0,0,93,0,176,0,112,0,171,0,8,0,97,0,141,0,190,0,210,0,196,0,99,0,0,0,83,0,86,0,63,0,0,0,247,0,213,0,221,0,4,0,196,0,206,0,252,0,129,0,87,0,207,0,198,0,0,0,198,0,164,0,238,0,50,0,71,0,0,0,139,0,28,0,195,0,193,0,0,0,0,0,133,0,52,0,84,0,16,0,0,0,237,0,71,0,37,0,248,0,226,0,2,0,160,0,83,0,0,0,69,0);
signal scenario_full  : scenario_type := (254,31,254,30,254,29,210,31,210,30,99,31,102,31,107,31,38,31,104,31,223,31,185,31,185,30,243,31,252,31,139,31,177,31,174,31,95,31,215,31,161,31,214,31,164,31,164,30,241,31,241,30,53,31,184,31,102,31,158,31,158,30,143,31,186,31,185,31,136,31,165,31,165,30,70,31,130,31,169,31,47,31,59,31,77,31,120,31,120,30,176,31,9,31,140,31,14,31,102,31,146,31,65,31,63,31,63,30,98,31,98,30,98,29,98,28,122,31,112,31,177,31,177,30,64,31,42,31,87,31,180,31,80,31,105,31,153,31,51,31,219,31,45,31,45,30,158,31,15,31,252,31,176,31,70,31,4,31,254,31,254,30,7,31,251,31,197,31,241,31,31,31,31,30,217,31,126,31,39,31,28,31,12,31,162,31,5,31,15,31,76,31,3,31,91,31,91,30,91,29,219,31,40,31,40,30,40,29,239,31,49,31,49,30,146,31,224,31,155,31,126,31,126,30,133,31,107,31,111,31,26,31,1,31,169,31,46,31,8,31,141,31,55,31,201,31,201,30,87,31,60,31,117,31,157,31,157,30,184,31,160,31,79,31,155,31,87,31,27,31,216,31,13,31,151,31,239,31,94,31,160,31,154,31,212,31,212,30,149,31,221,31,15,31,137,31,185,31,185,30,242,31,21,31,21,30,23,31,224,31,250,31,162,31,146,31,100,31,123,31,116,31,66,31,12,31,215,31,245,31,4,31,229,31,194,31,189,31,70,31,202,31,94,31,113,31,172,31,172,30,244,31,16,31,71,31,222,31,169,31,169,30,38,31,55,31,84,31,136,31,68,31,36,31,79,31,79,30,161,31,6,31,30,31,85,31,85,30,201,31,215,31,116,31,116,30,232,31,33,31,149,31,102,31,23,31,23,30,218,31,128,31,51,31,148,31,196,31,58,31,65,31,32,31,183,31,206,31,201,31,1,31,1,30,192,31,34,31,34,30,168,31,253,31,162,31,162,30,90,31,198,31,198,30,244,31,129,31,11,31,118,31,118,30,76,31,76,30,76,29,142,31,14,31,14,30,211,31,211,30,179,31,11,31,139,31,208,31,39,31,157,31,142,31,176,31,212,31,130,31,130,30,49,31,119,31,119,30,58,31,234,31,234,30,234,29,234,28,163,31,162,31,44,31,173,31,54,31,156,31,156,30,204,31,172,31,52,31,15,31,93,31,77,31,13,31,253,31,176,31,176,30,131,31,26,31,120,31,220,31,212,31,212,30,212,29,225,31,85,31,9,31,120,31,77,31,113,31,181,31,234,31,234,30,124,31,124,30,237,31,132,31,165,31,4,31,250,31,250,30,243,31,8,31,180,31,180,30,230,31,221,31,65,31,65,30,239,31,240,31,183,31,152,31,208,31,168,31,166,31,8,31,17,31,75,31,89,31,86,31,173,31,173,30,173,29,173,28,95,31,168,31,64,31,158,31,255,31,38,31,28,31,26,31,6,31,42,31,139,31,188,31,202,31,233,31,69,31,69,30,100,31,100,30,77,31,5,31,10,31,10,30,10,29,182,31,182,30,182,29,179,31,124,31,252,31,41,31,79,31,79,30,201,31,98,31,141,31,175,31,140,31,187,31,151,31,151,30,121,31,232,31,133,31,106,31,203,31,146,31,40,31,168,31,138,31,12,31,133,31,108,31,119,31,119,30,195,31,195,30,137,31,98,31,98,30,100,31,100,30,241,31,202,31,218,31,135,31,3,31,3,30,224,31,210,31,43,31,78,31,78,30,137,31,137,30,137,29,1,31,224,31,70,31,139,31,97,31,155,31,246,31,246,30,246,29,79,31,151,31,151,30,151,29,124,31,124,30,235,31,161,31,96,31,76,31,132,31,74,31,74,30,74,29,78,31,129,31,129,30,55,31,201,31,88,31,88,30,188,31,44,31,194,31,97,31,157,31,162,31,97,31,97,30,97,29,106,31,140,31,54,31,54,30,133,31,159,31,245,31,115,31,241,31,200,31,172,31,5,31,5,30,152,31,165,31,87,31,161,31,157,31,62,31,235,31,69,31,69,30,116,31,88,31,50,31,50,30,85,31,85,30,83,31,83,30,7,31,244,31,26,31,26,30,172,31,170,31,83,31,83,30,83,29,191,31,32,31,154,31,125,31,126,31,126,30,16,31,16,30,183,31,183,30,12,31,182,31,194,31,174,31,222,31,52,31,20,31,171,31,71,31,154,31,227,31,88,31,107,31,106,31,106,30,248,31,156,31,195,31,164,31,164,30,37,31,37,30,240,31,72,31,130,31,250,31,250,30,236,31,134,31,240,31,10,31,129,31,131,31,131,30,19,31,202,31,50,31,249,31,97,31,1,31,205,31,42,31,42,30,213,31,213,30,27,31,27,30,82,31,189,31,166,31,118,31,242,31,239,31,127,31,46,31,194,31,175,31,27,31,9,31,56,31,24,31,30,31,30,30,104,31,176,31,99,31,99,30,23,31,23,30,31,31,88,31,181,31,57,31,185,31,185,30,97,31,220,31,209,31,222,31,161,31,77,31,138,31,119,31,32,31,239,31,197,31,131,31,131,30,30,31,30,30,196,31,196,30,90,31,164,31,17,31,107,31,254,31,117,31,94,31,226,31,248,31,12,31,213,31,92,31,38,31,38,30,142,31,142,30,142,29,230,31,215,31,161,31,42,31,139,31,221,31,232,31,232,30,232,29,106,31,106,30,109,31,128,31,188,31,4,31,236,31,236,30,213,31,253,31,159,31,224,31,224,30,53,31,135,31,151,31,238,31,126,31,126,30,93,31,176,31,112,31,171,31,8,31,97,31,141,31,190,31,210,31,196,31,99,31,99,30,83,31,86,31,63,31,63,30,247,31,213,31,221,31,4,31,196,31,206,31,252,31,129,31,87,31,207,31,198,31,198,30,198,31,164,31,238,31,50,31,71,31,71,30,139,31,28,31,195,31,193,31,193,30,193,29,133,31,52,31,84,31,16,31,16,30,237,31,71,31,37,31,248,31,226,31,2,31,160,31,83,31,83,30,69,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
