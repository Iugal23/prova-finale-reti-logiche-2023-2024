-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_492 is
end project_tb_492;

architecture project_tb_arch_492 of project_tb_492 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 914;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (220,0,205,0,0,0,0,0,0,0,36,0,213,0,0,0,183,0,0,0,27,0,173,0,0,0,47,0,183,0,122,0,0,0,0,0,157,0,124,0,24,0,87,0,176,0,43,0,204,0,68,0,16,0,107,0,195,0,242,0,0,0,0,0,136,0,0,0,100,0,147,0,0,0,167,0,240,0,118,0,29,0,0,0,47,0,0,0,0,0,23,0,136,0,0,0,203,0,0,0,184,0,167,0,103,0,0,0,115,0,78,0,222,0,0,0,55,0,142,0,105,0,0,0,63,0,45,0,157,0,214,0,1,0,169,0,0,0,123,0,12,0,110,0,22,0,127,0,0,0,199,0,185,0,119,0,53,0,143,0,93,0,111,0,28,0,194,0,106,0,252,0,103,0,33,0,97,0,252,0,191,0,19,0,74,0,212,0,146,0,66,0,194,0,226,0,55,0,246,0,203,0,123,0,202,0,248,0,211,0,0,0,0,0,149,0,25,0,172,0,91,0,228,0,53,0,142,0,0,0,233,0,0,0,79,0,227,0,0,0,148,0,241,0,0,0,229,0,0,0,134,0,0,0,71,0,81,0,78,0,0,0,30,0,151,0,217,0,22,0,65,0,115,0,72,0,0,0,0,0,110,0,4,0,0,0,0,0,0,0,94,0,157,0,254,0,95,0,135,0,65,0,21,0,109,0,248,0,0,0,155,0,223,0,103,0,250,0,254,0,0,0,0,0,123,0,223,0,0,0,62,0,0,0,151,0,63,0,0,0,0,0,181,0,125,0,79,0,32,0,19,0,131,0,84,0,0,0,104,0,143,0,65,0,129,0,0,0,200,0,0,0,0,0,170,0,0,0,80,0,83,0,204,0,14,0,56,0,76,0,178,0,0,0,106,0,141,0,86,0,121,0,217,0,91,0,147,0,51,0,0,0,49,0,234,0,255,0,171,0,129,0,26,0,53,0,0,0,97,0,0,0,249,0,123,0,194,0,51,0,0,0,0,0,228,0,120,0,58,0,44,0,171,0,0,0,49,0,60,0,90,0,139,0,139,0,254,0,0,0,23,0,2,0,0,0,131,0,0,0,32,0,193,0,114,0,0,0,0,0,0,0,130,0,225,0,138,0,10,0,92,0,0,0,191,0,90,0,0,0,200,0,0,0,89,0,0,0,0,0,185,0,211,0,109,0,166,0,141,0,37,0,73,0,213,0,103,0,0,0,67,0,101,0,143,0,248,0,36,0,147,0,164,0,220,0,252,0,214,0,187,0,164,0,231,0,0,0,143,0,73,0,202,0,168,0,245,0,175,0,145,0,91,0,5,0,69,0,0,0,67,0,0,0,0,0,0,0,37,0,62,0,193,0,178,0,131,0,119,0,132,0,16,0,125,0,0,0,6,0,218,0,163,0,226,0,0,0,70,0,146,0,45,0,37,0,0,0,0,0,212,0,82,0,115,0,65,0,0,0,61,0,186,0,0,0,189,0,233,0,0,0,132,0,234,0,147,0,20,0,44,0,0,0,115,0,0,0,11,0,45,0,193,0,174,0,135,0,215,0,190,0,124,0,89,0,50,0,154,0,98,0,0,0,25,0,63,0,43,0,157,0,81,0,184,0,0,0,0,0,0,0,169,0,251,0,118,0,0,0,0,0,0,0,234,0,163,0,219,0,174,0,17,0,119,0,210,0,0,0,0,0,192,0,169,0,106,0,86,0,176,0,0,0,150,0,0,0,193,0,5,0,216,0,66,0,6,0,125,0,74,0,66,0,0,0,103,0,0,0,50,0,65,0,174,0,84,0,174,0,178,0,147,0,88,0,3,0,69,0,34,0,0,0,185,0,200,0,157,0,227,0,226,0,50,0,204,0,98,0,52,0,0,0,211,0,43,0,0,0,171,0,60,0,67,0,14,0,57,0,0,0,0,0,145,0,59,0,0,0,252,0,84,0,14,0,91,0,0,0,156,0,0,0,45,0,230,0,143,0,0,0,244,0,161,0,166,0,232,0,212,0,0,0,186,0,196,0,0,0,228,0,0,0,0,0,63,0,15,0,116,0,70,0,46,0,0,0,0,0,9,0,51,0,217,0,1,0,0,0,186,0,0,0,46,0,35,0,127,0,0,0,8,0,78,0,0,0,0,0,0,0,175,0,124,0,44,0,32,0,87,0,179,0,137,0,246,0,235,0,204,0,107,0,72,0,188,0,184,0,10,0,0,0,105,0,99,0,248,0,45,0,193,0,55,0,162,0,219,0,0,0,146,0,166,0,166,0,4,0,43,0,0,0,15,0,0,0,202,0,219,0,72,0,52,0,203,0,79,0,190,0,144,0,0,0,232,0,38,0,5,0,199,0,54,0,98,0,0,0,83,0,167,0,134,0,0,0,241,0,28,0,121,0,184,0,95,0,208,0,0,0,145,0,246,0,41,0,0,0,80,0,97,0,7,0,13,0,187,0,62,0,219,0,187,0,100,0,221,0,233,0,151,0,0,0,147,0,39,0,159,0,171,0,248,0,43,0,0,0,116,0,37,0,0,0,0,0,34,0,144,0,5,0,88,0,144,0,115,0,185,0,225,0,126,0,147,0,97,0,117,0,210,0,14,0,43,0,249,0,0,0,236,0,233,0,141,0,5,0,18,0,54,0,102,0,129,0,115,0,86,0,136,0,252,0,88,0,0,0,56,0,254,0,0,0,4,0,226,0,0,0,71,0,165,0,59,0,32,0,124,0,9,0,0,0,103,0,0,0,64,0,128,0,55,0,64,0,0,0,123,0,0,0,85,0,0,0,139,0,27,0,65,0,200,0,0,0,0,0,69,0,115,0,119,0,113,0,122,0,216,0,249,0,0,0,0,0,0,0,23,0,43,0,203,0,212,0,0,0,245,0,150,0,245,0,193,0,0,0,251,0,127,0,11,0,227,0,254,0,237,0,153,0,0,0,165,0,67,0,254,0,186,0,68,0,90,0,33,0,155,0,101,0,13,0,0,0,0,0,11,0,152,0,143,0,71,0,35,0,14,0,158,0,204,0,248,0,187,0,249,0,89,0,41,0,207,0,194,0,248,0,2,0,0,0,206,0,0,0,130,0,130,0,191,0,0,0,153,0,226,0,73,0,166,0,236,0,157,0,115,0,0,0,111,0,81,0,80,0,238,0,167,0,254,0,243,0,0,0,179,0,143,0,235,0,73,0,142,0,107,0,0,0,205,0,3,0,5,0,0,0,133,0,154,0,130,0,180,0,72,0,199,0,4,0,146,0,0,0,0,0,120,0,92,0,0,0,105,0,251,0,77,0,198,0,60,0,170,0,236,0,0,0,85,0,0,0,163,0,100,0,32,0,179,0,80,0,122,0,197,0,25,0,191,0,49,0,79,0,105,0,1,0,62,0,0,0,134,0,78,0,135,0,0,0,252,0,0,0,94,0,54,0,131,0,0,0,0,0,15,0,0,0,248,0,0,0,0,0,170,0,233,0,253,0,0,0,28,0,236,0,210,0,66,0,54,0,180,0,241,0,0,0,61,0,153,0,161,0,207,0,97,0,89,0,0,0,0,0,157,0,215,0,10,0,46,0,74,0,32,0,189,0,0,0,62,0,0,0,0,0,34,0,0,0,107,0,30,0,153,0,133,0,0,0,179,0,84,0,0,0,68,0,0,0,0,0,25,0,63,0,176,0,254,0,220,0,0,0,0,0,247,0,173,0,2,0,82,0,247,0,225,0,25,0,146,0,3,0,191,0,188,0,56,0,0,0,200,0,167,0,0,0,186,0,253,0,0,0,86,0,66,0,175,0,47,0,121,0,122,0,186,0,37,0,149,0,62,0,28,0,126,0,3,0,30,0,200,0,29,0,92,0,54,0,213,0,0,0,135,0,0,0,248,0,21,0,96,0,121,0,40,0,109,0,121,0,213,0,0,0,0,0,0,0,153,0,249,0,0,0,118,0,179,0,93,0,136,0,25,0,237,0,150,0,172,0,0,0,3,0,0,0,0,0,0,0,213,0,165,0,0,0,155,0,145,0,0,0,233,0,0,0,177,0,0,0,142,0,253,0,86,0,26,0,0,0,78,0,191,0,220,0,18,0,6,0,21,0,159,0,40,0,62,0,233,0);
signal scenario_full  : scenario_type := (220,31,205,31,205,30,205,29,205,28,36,31,213,31,213,30,183,31,183,30,27,31,173,31,173,30,47,31,183,31,122,31,122,30,122,29,157,31,124,31,24,31,87,31,176,31,43,31,204,31,68,31,16,31,107,31,195,31,242,31,242,30,242,29,136,31,136,30,100,31,147,31,147,30,167,31,240,31,118,31,29,31,29,30,47,31,47,30,47,29,23,31,136,31,136,30,203,31,203,30,184,31,167,31,103,31,103,30,115,31,78,31,222,31,222,30,55,31,142,31,105,31,105,30,63,31,45,31,157,31,214,31,1,31,169,31,169,30,123,31,12,31,110,31,22,31,127,31,127,30,199,31,185,31,119,31,53,31,143,31,93,31,111,31,28,31,194,31,106,31,252,31,103,31,33,31,97,31,252,31,191,31,19,31,74,31,212,31,146,31,66,31,194,31,226,31,55,31,246,31,203,31,123,31,202,31,248,31,211,31,211,30,211,29,149,31,25,31,172,31,91,31,228,31,53,31,142,31,142,30,233,31,233,30,79,31,227,31,227,30,148,31,241,31,241,30,229,31,229,30,134,31,134,30,71,31,81,31,78,31,78,30,30,31,151,31,217,31,22,31,65,31,115,31,72,31,72,30,72,29,110,31,4,31,4,30,4,29,4,28,94,31,157,31,254,31,95,31,135,31,65,31,21,31,109,31,248,31,248,30,155,31,223,31,103,31,250,31,254,31,254,30,254,29,123,31,223,31,223,30,62,31,62,30,151,31,63,31,63,30,63,29,181,31,125,31,79,31,32,31,19,31,131,31,84,31,84,30,104,31,143,31,65,31,129,31,129,30,200,31,200,30,200,29,170,31,170,30,80,31,83,31,204,31,14,31,56,31,76,31,178,31,178,30,106,31,141,31,86,31,121,31,217,31,91,31,147,31,51,31,51,30,49,31,234,31,255,31,171,31,129,31,26,31,53,31,53,30,97,31,97,30,249,31,123,31,194,31,51,31,51,30,51,29,228,31,120,31,58,31,44,31,171,31,171,30,49,31,60,31,90,31,139,31,139,31,254,31,254,30,23,31,2,31,2,30,131,31,131,30,32,31,193,31,114,31,114,30,114,29,114,28,130,31,225,31,138,31,10,31,92,31,92,30,191,31,90,31,90,30,200,31,200,30,89,31,89,30,89,29,185,31,211,31,109,31,166,31,141,31,37,31,73,31,213,31,103,31,103,30,67,31,101,31,143,31,248,31,36,31,147,31,164,31,220,31,252,31,214,31,187,31,164,31,231,31,231,30,143,31,73,31,202,31,168,31,245,31,175,31,145,31,91,31,5,31,69,31,69,30,67,31,67,30,67,29,67,28,37,31,62,31,193,31,178,31,131,31,119,31,132,31,16,31,125,31,125,30,6,31,218,31,163,31,226,31,226,30,70,31,146,31,45,31,37,31,37,30,37,29,212,31,82,31,115,31,65,31,65,30,61,31,186,31,186,30,189,31,233,31,233,30,132,31,234,31,147,31,20,31,44,31,44,30,115,31,115,30,11,31,45,31,193,31,174,31,135,31,215,31,190,31,124,31,89,31,50,31,154,31,98,31,98,30,25,31,63,31,43,31,157,31,81,31,184,31,184,30,184,29,184,28,169,31,251,31,118,31,118,30,118,29,118,28,234,31,163,31,219,31,174,31,17,31,119,31,210,31,210,30,210,29,192,31,169,31,106,31,86,31,176,31,176,30,150,31,150,30,193,31,5,31,216,31,66,31,6,31,125,31,74,31,66,31,66,30,103,31,103,30,50,31,65,31,174,31,84,31,174,31,178,31,147,31,88,31,3,31,69,31,34,31,34,30,185,31,200,31,157,31,227,31,226,31,50,31,204,31,98,31,52,31,52,30,211,31,43,31,43,30,171,31,60,31,67,31,14,31,57,31,57,30,57,29,145,31,59,31,59,30,252,31,84,31,14,31,91,31,91,30,156,31,156,30,45,31,230,31,143,31,143,30,244,31,161,31,166,31,232,31,212,31,212,30,186,31,196,31,196,30,228,31,228,30,228,29,63,31,15,31,116,31,70,31,46,31,46,30,46,29,9,31,51,31,217,31,1,31,1,30,186,31,186,30,46,31,35,31,127,31,127,30,8,31,78,31,78,30,78,29,78,28,175,31,124,31,44,31,32,31,87,31,179,31,137,31,246,31,235,31,204,31,107,31,72,31,188,31,184,31,10,31,10,30,105,31,99,31,248,31,45,31,193,31,55,31,162,31,219,31,219,30,146,31,166,31,166,31,4,31,43,31,43,30,15,31,15,30,202,31,219,31,72,31,52,31,203,31,79,31,190,31,144,31,144,30,232,31,38,31,5,31,199,31,54,31,98,31,98,30,83,31,167,31,134,31,134,30,241,31,28,31,121,31,184,31,95,31,208,31,208,30,145,31,246,31,41,31,41,30,80,31,97,31,7,31,13,31,187,31,62,31,219,31,187,31,100,31,221,31,233,31,151,31,151,30,147,31,39,31,159,31,171,31,248,31,43,31,43,30,116,31,37,31,37,30,37,29,34,31,144,31,5,31,88,31,144,31,115,31,185,31,225,31,126,31,147,31,97,31,117,31,210,31,14,31,43,31,249,31,249,30,236,31,233,31,141,31,5,31,18,31,54,31,102,31,129,31,115,31,86,31,136,31,252,31,88,31,88,30,56,31,254,31,254,30,4,31,226,31,226,30,71,31,165,31,59,31,32,31,124,31,9,31,9,30,103,31,103,30,64,31,128,31,55,31,64,31,64,30,123,31,123,30,85,31,85,30,139,31,27,31,65,31,200,31,200,30,200,29,69,31,115,31,119,31,113,31,122,31,216,31,249,31,249,30,249,29,249,28,23,31,43,31,203,31,212,31,212,30,245,31,150,31,245,31,193,31,193,30,251,31,127,31,11,31,227,31,254,31,237,31,153,31,153,30,165,31,67,31,254,31,186,31,68,31,90,31,33,31,155,31,101,31,13,31,13,30,13,29,11,31,152,31,143,31,71,31,35,31,14,31,158,31,204,31,248,31,187,31,249,31,89,31,41,31,207,31,194,31,248,31,2,31,2,30,206,31,206,30,130,31,130,31,191,31,191,30,153,31,226,31,73,31,166,31,236,31,157,31,115,31,115,30,111,31,81,31,80,31,238,31,167,31,254,31,243,31,243,30,179,31,143,31,235,31,73,31,142,31,107,31,107,30,205,31,3,31,5,31,5,30,133,31,154,31,130,31,180,31,72,31,199,31,4,31,146,31,146,30,146,29,120,31,92,31,92,30,105,31,251,31,77,31,198,31,60,31,170,31,236,31,236,30,85,31,85,30,163,31,100,31,32,31,179,31,80,31,122,31,197,31,25,31,191,31,49,31,79,31,105,31,1,31,62,31,62,30,134,31,78,31,135,31,135,30,252,31,252,30,94,31,54,31,131,31,131,30,131,29,15,31,15,30,248,31,248,30,248,29,170,31,233,31,253,31,253,30,28,31,236,31,210,31,66,31,54,31,180,31,241,31,241,30,61,31,153,31,161,31,207,31,97,31,89,31,89,30,89,29,157,31,215,31,10,31,46,31,74,31,32,31,189,31,189,30,62,31,62,30,62,29,34,31,34,30,107,31,30,31,153,31,133,31,133,30,179,31,84,31,84,30,68,31,68,30,68,29,25,31,63,31,176,31,254,31,220,31,220,30,220,29,247,31,173,31,2,31,82,31,247,31,225,31,25,31,146,31,3,31,191,31,188,31,56,31,56,30,200,31,167,31,167,30,186,31,253,31,253,30,86,31,66,31,175,31,47,31,121,31,122,31,186,31,37,31,149,31,62,31,28,31,126,31,3,31,30,31,200,31,29,31,92,31,54,31,213,31,213,30,135,31,135,30,248,31,21,31,96,31,121,31,40,31,109,31,121,31,213,31,213,30,213,29,213,28,153,31,249,31,249,30,118,31,179,31,93,31,136,31,25,31,237,31,150,31,172,31,172,30,3,31,3,30,3,29,3,28,213,31,165,31,165,30,155,31,145,31,145,30,233,31,233,30,177,31,177,30,142,31,253,31,86,31,26,31,26,30,78,31,191,31,220,31,18,31,6,31,21,31,159,31,40,31,62,31,233,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
