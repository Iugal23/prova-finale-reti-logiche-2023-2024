-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 775;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (203,0,101,0,73,0,223,0,195,0,116,0,23,0,125,0,189,0,24,0,240,0,73,0,125,0,69,0,14,0,68,0,67,0,168,0,193,0,138,0,65,0,234,0,216,0,107,0,184,0,226,0,21,0,172,0,129,0,23,0,234,0,251,0,224,0,135,0,35,0,203,0,188,0,87,0,225,0,174,0,192,0,41,0,55,0,0,0,12,0,243,0,27,0,205,0,231,0,17,0,50,0,131,0,158,0,71,0,18,0,91,0,31,0,135,0,68,0,90,0,169,0,0,0,156,0,0,0,250,0,180,0,210,0,35,0,73,0,0,0,0,0,0,0,143,0,223,0,142,0,0,0,0,0,0,0,0,0,0,0,28,0,160,0,0,0,239,0,228,0,95,0,60,0,0,0,134,0,216,0,42,0,223,0,147,0,222,0,178,0,0,0,164,0,0,0,189,0,161,0,228,0,114,0,69,0,128,0,43,0,0,0,75,0,218,0,79,0,2,0,4,0,173,0,160,0,210,0,41,0,6,0,0,0,88,0,162,0,146,0,250,0,1,0,215,0,46,0,34,0,223,0,110,0,87,0,121,0,232,0,0,0,78,0,128,0,126,0,0,0,187,0,76,0,139,0,46,0,216,0,0,0,34,0,21,0,36,0,138,0,148,0,46,0,42,0,77,0,94,0,0,0,19,0,40,0,87,0,62,0,246,0,231,0,150,0,244,0,173,0,252,0,32,0,248,0,175,0,0,0,209,0,100,0,80,0,189,0,251,0,244,0,0,0,48,0,149,0,80,0,16,0,0,0,219,0,230,0,146,0,125,0,66,0,179,0,166,0,1,0,16,0,29,0,134,0,82,0,10,0,204,0,94,0,0,0,190,0,178,0,239,0,71,0,204,0,228,0,12,0,126,0,125,0,0,0,2,0,19,0,93,0,155,0,178,0,0,0,184,0,23,0,6,0,8,0,180,0,48,0,174,0,50,0,135,0,171,0,204,0,0,0,108,0,171,0,0,0,172,0,49,0,0,0,193,0,238,0,0,0,225,0,222,0,219,0,123,0,171,0,84,0,56,0,0,0,0,0,0,0,0,0,66,0,43,0,182,0,159,0,235,0,51,0,222,0,168,0,0,0,34,0,150,0,162,0,220,0,0,0,4,0,61,0,0,0,20,0,142,0,224,0,204,0,130,0,0,0,192,0,40,0,49,0,238,0,236,0,78,0,136,0,248,0,0,0,22,0,231,0,86,0,101,0,0,0,8,0,230,0,0,0,95,0,239,0,15,0,121,0,154,0,137,0,250,0,0,0,70,0,168,0,178,0,74,0,0,0,0,0,30,0,0,0,122,0,111,0,36,0,228,0,11,0,61,0,212,0,35,0,0,0,0,0,137,0,153,0,93,0,5,0,0,0,0,0,0,0,99,0,0,0,237,0,43,0,141,0,72,0,4,0,123,0,125,0,19,0,0,0,32,0,160,0,238,0,0,0,241,0,0,0,208,0,243,0,0,0,228,0,243,0,95,0,4,0,66,0,156,0,95,0,136,0,0,0,187,0,0,0,53,0,231,0,1,0,0,0,102,0,102,0,50,0,0,0,138,0,102,0,0,0,0,0,26,0,0,0,110,0,0,0,104,0,66,0,228,0,0,0,41,0,0,0,143,0,60,0,9,0,19,0,249,0,133,0,227,0,235,0,205,0,186,0,51,0,90,0,14,0,50,0,212,0,124,0,89,0,199,0,210,0,123,0,243,0,21,0,0,0,0,0,123,0,171,0,39,0,2,0,121,0,232,0,224,0,0,0,0,0,39,0,0,0,50,0,39,0,38,0,0,0,26,0,158,0,0,0,217,0,65,0,43,0,59,0,13,0,129,0,71,0,0,0,221,0,194,0,0,0,98,0,226,0,32,0,0,0,107,0,49,0,0,0,124,0,36,0,56,0,119,0,0,0,7,0,78,0,103,0,13,0,228,0,195,0,205,0,163,0,111,0,113,0,124,0,80,0,0,0,0,0,192,0,211,0,0,0,28,0,221,0,0,0,120,0,85,0,198,0,0,0,183,0,151,0,147,0,0,0,0,0,25,0,102,0,0,0,69,0,219,0,113,0,124,0,215,0,0,0,100,0,0,0,100,0,134,0,190,0,134,0,151,0,0,0,0,0,0,0,141,0,221,0,64,0,59,0,48,0,0,0,69,0,123,0,254,0,239,0,208,0,83,0,64,0,75,0,175,0,216,0,191,0,146,0,31,0,106,0,0,0,0,0,66,0,33,0,144,0,199,0,255,0,0,0,42,0,134,0,249,0,87,0,33,0,8,0,157,0,201,0,150,0,234,0,225,0,92,0,217,0,11,0,65,0,0,0,242,0,109,0,237,0,0,0,88,0,217,0,187,0,0,0,96,0,56,0,0,0,242,0,73,0,177,0,162,0,47,0,123,0,140,0,101,0,73,0,253,0,170,0,0,0,199,0,45,0,0,0,91,0,116,0,16,0,205,0,217,0,98,0,162,0,154,0,252,0,23,0,145,0,55,0,53,0,64,0,34,0,0,0,115,0,0,0,0,0,60,0,98,0,77,0,96,0,236,0,237,0,0,0,63,0,227,0,178,0,0,0,63,0,66,0,219,0,67,0,33,0,89,0,209,0,13,0,248,0,183,0,74,0,51,0,0,0,0,0,137,0,0,0,126,0,0,0,231,0,85,0,0,0,177,0,143,0,191,0,187,0,46,0,161,0,27,0,0,0,75,0,91,0,76,0,237,0,0,0,59,0,174,0,244,0,74,0,0,0,230,0,122,0,156,0,1,0,5,0,207,0,94,0,236,0,134,0,35,0,23,0,44,0,32,0,0,0,164,0,126,0,25,0,148,0,195,0,166,0,218,0,0,0,199,0,54,0,106,0,92,0,7,0,161,0,171,0,83,0,229,0,2,0,0,0,134,0,243,0,219,0,190,0,105,0,170,0,52,0,0,0,122,0,176,0,0,0,0,0,0,0,104,0,112,0,117,0,26,0,105,0,206,0,47,0,151,0,162,0,182,0,26,0,74,0,205,0,84,0,0,0,118,0,80,0,0,0,200,0,124,0,102,0,0,0,31,0,192,0,214,0,227,0,0,0,224,0,165,0,228,0,0,0,109,0,125,0,100,0,0,0,107,0,89,0,255,0,0,0,0,0,243,0,242,0,17,0,18,0,43,0,211,0,0,0,0,0,46,0,235,0,0,0,68,0,23,0,214,0,70,0,206,0,220,0,0,0,223,0,21,0,251,0,221,0,117,0,137,0,175,0,0,0,121,0,0,0,0,0,18,0,46,0,0,0,182,0,242,0,0,0,0,0,175,0,123,0,65,0,184,0,0,0,130,0,0,0,204,0,128,0,178,0,8,0,67,0,0,0,240,0,0,0,0,0,226,0,163,0,143,0,211,0,63,0,123,0,84,0,123,0,248,0,94,0,150,0,252,0,33,0,17,0,175,0,0,0,0,0,0,0);
signal scenario_full  : scenario_type := (203,31,101,31,73,31,223,31,195,31,116,31,23,31,125,31,189,31,24,31,240,31,73,31,125,31,69,31,14,31,68,31,67,31,168,31,193,31,138,31,65,31,234,31,216,31,107,31,184,31,226,31,21,31,172,31,129,31,23,31,234,31,251,31,224,31,135,31,35,31,203,31,188,31,87,31,225,31,174,31,192,31,41,31,55,31,55,30,12,31,243,31,27,31,205,31,231,31,17,31,50,31,131,31,158,31,71,31,18,31,91,31,31,31,135,31,68,31,90,31,169,31,169,30,156,31,156,30,250,31,180,31,210,31,35,31,73,31,73,30,73,29,73,28,143,31,223,31,142,31,142,30,142,29,142,28,142,27,142,26,28,31,160,31,160,30,239,31,228,31,95,31,60,31,60,30,134,31,216,31,42,31,223,31,147,31,222,31,178,31,178,30,164,31,164,30,189,31,161,31,228,31,114,31,69,31,128,31,43,31,43,30,75,31,218,31,79,31,2,31,4,31,173,31,160,31,210,31,41,31,6,31,6,30,88,31,162,31,146,31,250,31,1,31,215,31,46,31,34,31,223,31,110,31,87,31,121,31,232,31,232,30,78,31,128,31,126,31,126,30,187,31,76,31,139,31,46,31,216,31,216,30,34,31,21,31,36,31,138,31,148,31,46,31,42,31,77,31,94,31,94,30,19,31,40,31,87,31,62,31,246,31,231,31,150,31,244,31,173,31,252,31,32,31,248,31,175,31,175,30,209,31,100,31,80,31,189,31,251,31,244,31,244,30,48,31,149,31,80,31,16,31,16,30,219,31,230,31,146,31,125,31,66,31,179,31,166,31,1,31,16,31,29,31,134,31,82,31,10,31,204,31,94,31,94,30,190,31,178,31,239,31,71,31,204,31,228,31,12,31,126,31,125,31,125,30,2,31,19,31,93,31,155,31,178,31,178,30,184,31,23,31,6,31,8,31,180,31,48,31,174,31,50,31,135,31,171,31,204,31,204,30,108,31,171,31,171,30,172,31,49,31,49,30,193,31,238,31,238,30,225,31,222,31,219,31,123,31,171,31,84,31,56,31,56,30,56,29,56,28,56,27,66,31,43,31,182,31,159,31,235,31,51,31,222,31,168,31,168,30,34,31,150,31,162,31,220,31,220,30,4,31,61,31,61,30,20,31,142,31,224,31,204,31,130,31,130,30,192,31,40,31,49,31,238,31,236,31,78,31,136,31,248,31,248,30,22,31,231,31,86,31,101,31,101,30,8,31,230,31,230,30,95,31,239,31,15,31,121,31,154,31,137,31,250,31,250,30,70,31,168,31,178,31,74,31,74,30,74,29,30,31,30,30,122,31,111,31,36,31,228,31,11,31,61,31,212,31,35,31,35,30,35,29,137,31,153,31,93,31,5,31,5,30,5,29,5,28,99,31,99,30,237,31,43,31,141,31,72,31,4,31,123,31,125,31,19,31,19,30,32,31,160,31,238,31,238,30,241,31,241,30,208,31,243,31,243,30,228,31,243,31,95,31,4,31,66,31,156,31,95,31,136,31,136,30,187,31,187,30,53,31,231,31,1,31,1,30,102,31,102,31,50,31,50,30,138,31,102,31,102,30,102,29,26,31,26,30,110,31,110,30,104,31,66,31,228,31,228,30,41,31,41,30,143,31,60,31,9,31,19,31,249,31,133,31,227,31,235,31,205,31,186,31,51,31,90,31,14,31,50,31,212,31,124,31,89,31,199,31,210,31,123,31,243,31,21,31,21,30,21,29,123,31,171,31,39,31,2,31,121,31,232,31,224,31,224,30,224,29,39,31,39,30,50,31,39,31,38,31,38,30,26,31,158,31,158,30,217,31,65,31,43,31,59,31,13,31,129,31,71,31,71,30,221,31,194,31,194,30,98,31,226,31,32,31,32,30,107,31,49,31,49,30,124,31,36,31,56,31,119,31,119,30,7,31,78,31,103,31,13,31,228,31,195,31,205,31,163,31,111,31,113,31,124,31,80,31,80,30,80,29,192,31,211,31,211,30,28,31,221,31,221,30,120,31,85,31,198,31,198,30,183,31,151,31,147,31,147,30,147,29,25,31,102,31,102,30,69,31,219,31,113,31,124,31,215,31,215,30,100,31,100,30,100,31,134,31,190,31,134,31,151,31,151,30,151,29,151,28,141,31,221,31,64,31,59,31,48,31,48,30,69,31,123,31,254,31,239,31,208,31,83,31,64,31,75,31,175,31,216,31,191,31,146,31,31,31,106,31,106,30,106,29,66,31,33,31,144,31,199,31,255,31,255,30,42,31,134,31,249,31,87,31,33,31,8,31,157,31,201,31,150,31,234,31,225,31,92,31,217,31,11,31,65,31,65,30,242,31,109,31,237,31,237,30,88,31,217,31,187,31,187,30,96,31,56,31,56,30,242,31,73,31,177,31,162,31,47,31,123,31,140,31,101,31,73,31,253,31,170,31,170,30,199,31,45,31,45,30,91,31,116,31,16,31,205,31,217,31,98,31,162,31,154,31,252,31,23,31,145,31,55,31,53,31,64,31,34,31,34,30,115,31,115,30,115,29,60,31,98,31,77,31,96,31,236,31,237,31,237,30,63,31,227,31,178,31,178,30,63,31,66,31,219,31,67,31,33,31,89,31,209,31,13,31,248,31,183,31,74,31,51,31,51,30,51,29,137,31,137,30,126,31,126,30,231,31,85,31,85,30,177,31,143,31,191,31,187,31,46,31,161,31,27,31,27,30,75,31,91,31,76,31,237,31,237,30,59,31,174,31,244,31,74,31,74,30,230,31,122,31,156,31,1,31,5,31,207,31,94,31,236,31,134,31,35,31,23,31,44,31,32,31,32,30,164,31,126,31,25,31,148,31,195,31,166,31,218,31,218,30,199,31,54,31,106,31,92,31,7,31,161,31,171,31,83,31,229,31,2,31,2,30,134,31,243,31,219,31,190,31,105,31,170,31,52,31,52,30,122,31,176,31,176,30,176,29,176,28,104,31,112,31,117,31,26,31,105,31,206,31,47,31,151,31,162,31,182,31,26,31,74,31,205,31,84,31,84,30,118,31,80,31,80,30,200,31,124,31,102,31,102,30,31,31,192,31,214,31,227,31,227,30,224,31,165,31,228,31,228,30,109,31,125,31,100,31,100,30,107,31,89,31,255,31,255,30,255,29,243,31,242,31,17,31,18,31,43,31,211,31,211,30,211,29,46,31,235,31,235,30,68,31,23,31,214,31,70,31,206,31,220,31,220,30,223,31,21,31,251,31,221,31,117,31,137,31,175,31,175,30,121,31,121,30,121,29,18,31,46,31,46,30,182,31,242,31,242,30,242,29,175,31,123,31,65,31,184,31,184,30,130,31,130,30,204,31,128,31,178,31,8,31,67,31,67,30,240,31,240,30,240,29,226,31,163,31,143,31,211,31,63,31,123,31,84,31,123,31,248,31,94,31,150,31,252,31,33,31,17,31,175,31,175,30,175,29,175,28);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
