-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_455 is
end project_tb_455;

architecture project_tb_arch_455 of project_tb_455 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 895;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,136,0,52,0,51,0,19,0,72,0,140,0,213,0,213,0,174,0,0,0,0,0,92,0,79,0,54,0,0,0,187,0,170,0,228,0,0,0,0,0,0,0,78,0,11,0,130,0,106,0,0,0,1,0,67,0,189,0,0,0,0,0,172,0,216,0,0,0,0,0,249,0,52,0,149,0,137,0,42,0,190,0,115,0,170,0,172,0,70,0,140,0,89,0,8,0,167,0,206,0,0,0,181,0,0,0,12,0,43,0,0,0,11,0,13,0,139,0,169,0,197,0,108,0,96,0,0,0,31,0,218,0,39,0,224,0,0,0,26,0,221,0,100,0,0,0,0,0,111,0,140,0,72,0,21,0,180,0,0,0,38,0,133,0,28,0,225,0,121,0,228,0,83,0,35,0,37,0,250,0,0,0,220,0,0,0,0,0,3,0,131,0,147,0,177,0,187,0,21,0,0,0,48,0,213,0,0,0,0,0,219,0,0,0,201,0,253,0,2,0,194,0,81,0,99,0,0,0,0,0,5,0,99,0,48,0,38,0,45,0,129,0,136,0,43,0,229,0,169,0,149,0,177,0,96,0,223,0,231,0,9,0,56,0,215,0,109,0,75,0,118,0,0,0,26,0,124,0,0,0,221,0,206,0,0,0,114,0,1,0,187,0,30,0,11,0,192,0,172,0,0,0,66,0,0,0,39,0,0,0,194,0,55,0,224,0,0,0,249,0,103,0,70,0,68,0,46,0,185,0,79,0,144,0,67,0,190,0,0,0,84,0,0,0,70,0,103,0,246,0,66,0,0,0,0,0,30,0,177,0,0,0,68,0,67,0,240,0,83,0,23,0,225,0,146,0,68,0,126,0,68,0,97,0,61,0,33,0,0,0,0,0,0,0,78,0,121,0,150,0,244,0,11,0,104,0,198,0,195,0,0,0,0,0,237,0,200,0,130,0,0,0,77,0,220,0,0,0,10,0,0,0,232,0,51,0,0,0,221,0,208,0,226,0,0,0,143,0,0,0,0,0,243,0,194,0,0,0,0,0,172,0,207,0,245,0,91,0,16,0,0,0,172,0,126,0,201,0,255,0,0,0,5,0,121,0,120,0,139,0,72,0,218,0,164,0,24,0,134,0,199,0,0,0,188,0,219,0,210,0,0,0,81,0,181,0,66,0,173,0,201,0,3,0,186,0,10,0,0,0,91,0,170,0,91,0,228,0,0,0,23,0,141,0,210,0,53,0,201,0,42,0,204,0,29,0,114,0,0,0,63,0,59,0,79,0,186,0,235,0,0,0,0,0,233,0,135,0,0,0,106,0,0,0,52,0,247,0,0,0,250,0,115,0,226,0,151,0,0,0,5,0,140,0,138,0,88,0,171,0,217,0,59,0,174,0,79,0,252,0,29,0,18,0,126,0,248,0,240,0,70,0,120,0,89,0,8,0,0,0,0,0,142,0,68,0,86,0,77,0,0,0,0,0,250,0,213,0,155,0,104,0,219,0,209,0,0,0,18,0,30,0,101,0,203,0,0,0,198,0,78,0,124,0,18,0,110,0,246,0,0,0,36,0,14,0,41,0,255,0,3,0,42,0,198,0,105,0,175,0,0,0,126,0,174,0,7,0,14,0,218,0,177,0,94,0,70,0,85,0,194,0,201,0,0,0,139,0,237,0,108,0,89,0,230,0,60,0,160,0,189,0,0,0,113,0,100,0,186,0,0,0,201,0,27,0,199,0,0,0,0,0,159,0,0,0,242,0,182,0,18,0,128,0,237,0,0,0,94,0,92,0,157,0,16,0,121,0,136,0,131,0,40,0,91,0,63,0,12,0,0,0,9,0,0,0,254,0,0,0,175,0,97,0,147,0,0,0,171,0,61,0,151,0,186,0,0,0,136,0,29,0,53,0,40,0,9,0,103,0,0,0,238,0,155,0,0,0,221,0,70,0,29,0,215,0,133,0,125,0,230,0,65,0,86,0,0,0,144,0,0,0,139,0,148,0,248,0,0,0,71,0,235,0,118,0,0,0,205,0,75,0,86,0,33,0,138,0,14,0,0,0,11,0,49,0,0,0,211,0,0,0,189,0,116,0,0,0,173,0,19,0,159,0,2,0,149,0,47,0,104,0,102,0,109,0,0,0,0,0,122,0,3,0,0,0,106,0,150,0,213,0,196,0,190,0,75,0,249,0,97,0,2,0,206,0,0,0,149,0,217,0,101,0,16,0,105,0,0,0,69,0,114,0,195,0,28,0,76,0,9,0,202,0,157,0,5,0,24,0,111,0,0,0,137,0,45,0,99,0,0,0,0,0,55,0,0,0,74,0,4,0,0,0,254,0,159,0,243,0,71,0,44,0,27,0,76,0,0,0,94,0,217,0,84,0,152,0,160,0,15,0,54,0,47,0,93,0,207,0,0,0,0,0,239,0,108,0,193,0,86,0,147,0,0,0,0,0,138,0,46,0,0,0,56,0,2,0,108,0,0,0,1,0,93,0,115,0,188,0,42,0,112,0,0,0,181,0,0,0,61,0,140,0,12,0,113,0,0,0,252,0,135,0,0,0,232,0,0,0,196,0,99,0,210,0,99,0,0,0,176,0,182,0,76,0,81,0,108,0,242,0,172,0,104,0,0,0,189,0,253,0,242,0,177,0,48,0,120,0,49,0,0,0,40,0,0,0,54,0,78,0,0,0,0,0,175,0,0,0,220,0,254,0,0,0,159,0,65,0,204,0,79,0,131,0,102,0,76,0,0,0,0,0,115,0,91,0,23,0,44,0,138,0,0,0,90,0,0,0,13,0,160,0,155,0,200,0,0,0,187,0,151,0,252,0,88,0,251,0,0,0,41,0,70,0,178,0,162,0,36,0,119,0,0,0,63,0,0,0,0,0,6,0,16,0,133,0,0,0,185,0,121,0,245,0,0,0,123,0,0,0,242,0,106,0,0,0,252,0,96,0,202,0,0,0,237,0,65,0,249,0,77,0,242,0,200,0,142,0,49,0,0,0,169,0,64,0,235,0,105,0,85,0,225,0,232,0,174,0,184,0,0,0,9,0,183,0,178,0,124,0,170,0,0,0,27,0,17,0,85,0,197,0,41,0,180,0,126,0,212,0,221,0,186,0,253,0,224,0,0,0,195,0,4,0,178,0,45,0,164,0,232,0,122,0,172,0,237,0,121,0,191,0,98,0,189,0,20,0,0,0,130,0,12,0,179,0,104,0,56,0,81,0,253,0,79,0,136,0,63,0,146,0,16,0,14,0,83,0,0,0,122,0,0,0,129,0,0,0,30,0,248,0,58,0,0,0,179,0,181,0,116,0,65,0,0,0,0,0,236,0,124,0,209,0,25,0,26,0,0,0,189,0,218,0,185,0,154,0,19,0,13,0,218,0,33,0,0,0,0,0,196,0,78,0,148,0,175,0,0,0,152,0,212,0,0,0,114,0,247,0,167,0,175,0,59,0,154,0,84,0,151,0,141,0,241,0,63,0,224,0,169,0,146,0,40,0,69,0,0,0,47,0,94,0,217,0,196,0,0,0,0,0,146,0,226,0,93,0,121,0,51,0,208,0,117,0,233,0,231,0,0,0,200,0,69,0,70,0,17,0,248,0,113,0,44,0,245,0,221,0,247,0,30,0,48,0,72,0,55,0,0,0,79,0,68,0,227,0,188,0,107,0,116,0,212,0,0,0,88,0,0,0,190,0,79,0,253,0,95,0,107,0,0,0,15,0,0,0,0,0,61,0,74,0,6,0,125,0,171,0,229,0,123,0,100,0,246,0,50,0,50,0,18,0,237,0,77,0,6,0,36,0,0,0,239,0,251,0,199,0,127,0,132,0,53,0,0,0,68,0,0,0,198,0,147,0,167,0,144,0,15,0,221,0,108,0,234,0,0,0,110,0,30,0,121,0,211,0,232,0,22,0,188,0,9,0,60,0,187,0,82,0,139,0,119,0,123,0,0,0,75,0,255,0,110,0,3,0,184,0,82,0,0,0,98,0,45,0,0,0,4,0,2,0,247,0);
signal scenario_full  : scenario_type := (0,0,136,31,52,31,51,31,19,31,72,31,140,31,213,31,213,31,174,31,174,30,174,29,92,31,79,31,54,31,54,30,187,31,170,31,228,31,228,30,228,29,228,28,78,31,11,31,130,31,106,31,106,30,1,31,67,31,189,31,189,30,189,29,172,31,216,31,216,30,216,29,249,31,52,31,149,31,137,31,42,31,190,31,115,31,170,31,172,31,70,31,140,31,89,31,8,31,167,31,206,31,206,30,181,31,181,30,12,31,43,31,43,30,11,31,13,31,139,31,169,31,197,31,108,31,96,31,96,30,31,31,218,31,39,31,224,31,224,30,26,31,221,31,100,31,100,30,100,29,111,31,140,31,72,31,21,31,180,31,180,30,38,31,133,31,28,31,225,31,121,31,228,31,83,31,35,31,37,31,250,31,250,30,220,31,220,30,220,29,3,31,131,31,147,31,177,31,187,31,21,31,21,30,48,31,213,31,213,30,213,29,219,31,219,30,201,31,253,31,2,31,194,31,81,31,99,31,99,30,99,29,5,31,99,31,48,31,38,31,45,31,129,31,136,31,43,31,229,31,169,31,149,31,177,31,96,31,223,31,231,31,9,31,56,31,215,31,109,31,75,31,118,31,118,30,26,31,124,31,124,30,221,31,206,31,206,30,114,31,1,31,187,31,30,31,11,31,192,31,172,31,172,30,66,31,66,30,39,31,39,30,194,31,55,31,224,31,224,30,249,31,103,31,70,31,68,31,46,31,185,31,79,31,144,31,67,31,190,31,190,30,84,31,84,30,70,31,103,31,246,31,66,31,66,30,66,29,30,31,177,31,177,30,68,31,67,31,240,31,83,31,23,31,225,31,146,31,68,31,126,31,68,31,97,31,61,31,33,31,33,30,33,29,33,28,78,31,121,31,150,31,244,31,11,31,104,31,198,31,195,31,195,30,195,29,237,31,200,31,130,31,130,30,77,31,220,31,220,30,10,31,10,30,232,31,51,31,51,30,221,31,208,31,226,31,226,30,143,31,143,30,143,29,243,31,194,31,194,30,194,29,172,31,207,31,245,31,91,31,16,31,16,30,172,31,126,31,201,31,255,31,255,30,5,31,121,31,120,31,139,31,72,31,218,31,164,31,24,31,134,31,199,31,199,30,188,31,219,31,210,31,210,30,81,31,181,31,66,31,173,31,201,31,3,31,186,31,10,31,10,30,91,31,170,31,91,31,228,31,228,30,23,31,141,31,210,31,53,31,201,31,42,31,204,31,29,31,114,31,114,30,63,31,59,31,79,31,186,31,235,31,235,30,235,29,233,31,135,31,135,30,106,31,106,30,52,31,247,31,247,30,250,31,115,31,226,31,151,31,151,30,5,31,140,31,138,31,88,31,171,31,217,31,59,31,174,31,79,31,252,31,29,31,18,31,126,31,248,31,240,31,70,31,120,31,89,31,8,31,8,30,8,29,142,31,68,31,86,31,77,31,77,30,77,29,250,31,213,31,155,31,104,31,219,31,209,31,209,30,18,31,30,31,101,31,203,31,203,30,198,31,78,31,124,31,18,31,110,31,246,31,246,30,36,31,14,31,41,31,255,31,3,31,42,31,198,31,105,31,175,31,175,30,126,31,174,31,7,31,14,31,218,31,177,31,94,31,70,31,85,31,194,31,201,31,201,30,139,31,237,31,108,31,89,31,230,31,60,31,160,31,189,31,189,30,113,31,100,31,186,31,186,30,201,31,27,31,199,31,199,30,199,29,159,31,159,30,242,31,182,31,18,31,128,31,237,31,237,30,94,31,92,31,157,31,16,31,121,31,136,31,131,31,40,31,91,31,63,31,12,31,12,30,9,31,9,30,254,31,254,30,175,31,97,31,147,31,147,30,171,31,61,31,151,31,186,31,186,30,136,31,29,31,53,31,40,31,9,31,103,31,103,30,238,31,155,31,155,30,221,31,70,31,29,31,215,31,133,31,125,31,230,31,65,31,86,31,86,30,144,31,144,30,139,31,148,31,248,31,248,30,71,31,235,31,118,31,118,30,205,31,75,31,86,31,33,31,138,31,14,31,14,30,11,31,49,31,49,30,211,31,211,30,189,31,116,31,116,30,173,31,19,31,159,31,2,31,149,31,47,31,104,31,102,31,109,31,109,30,109,29,122,31,3,31,3,30,106,31,150,31,213,31,196,31,190,31,75,31,249,31,97,31,2,31,206,31,206,30,149,31,217,31,101,31,16,31,105,31,105,30,69,31,114,31,195,31,28,31,76,31,9,31,202,31,157,31,5,31,24,31,111,31,111,30,137,31,45,31,99,31,99,30,99,29,55,31,55,30,74,31,4,31,4,30,254,31,159,31,243,31,71,31,44,31,27,31,76,31,76,30,94,31,217,31,84,31,152,31,160,31,15,31,54,31,47,31,93,31,207,31,207,30,207,29,239,31,108,31,193,31,86,31,147,31,147,30,147,29,138,31,46,31,46,30,56,31,2,31,108,31,108,30,1,31,93,31,115,31,188,31,42,31,112,31,112,30,181,31,181,30,61,31,140,31,12,31,113,31,113,30,252,31,135,31,135,30,232,31,232,30,196,31,99,31,210,31,99,31,99,30,176,31,182,31,76,31,81,31,108,31,242,31,172,31,104,31,104,30,189,31,253,31,242,31,177,31,48,31,120,31,49,31,49,30,40,31,40,30,54,31,78,31,78,30,78,29,175,31,175,30,220,31,254,31,254,30,159,31,65,31,204,31,79,31,131,31,102,31,76,31,76,30,76,29,115,31,91,31,23,31,44,31,138,31,138,30,90,31,90,30,13,31,160,31,155,31,200,31,200,30,187,31,151,31,252,31,88,31,251,31,251,30,41,31,70,31,178,31,162,31,36,31,119,31,119,30,63,31,63,30,63,29,6,31,16,31,133,31,133,30,185,31,121,31,245,31,245,30,123,31,123,30,242,31,106,31,106,30,252,31,96,31,202,31,202,30,237,31,65,31,249,31,77,31,242,31,200,31,142,31,49,31,49,30,169,31,64,31,235,31,105,31,85,31,225,31,232,31,174,31,184,31,184,30,9,31,183,31,178,31,124,31,170,31,170,30,27,31,17,31,85,31,197,31,41,31,180,31,126,31,212,31,221,31,186,31,253,31,224,31,224,30,195,31,4,31,178,31,45,31,164,31,232,31,122,31,172,31,237,31,121,31,191,31,98,31,189,31,20,31,20,30,130,31,12,31,179,31,104,31,56,31,81,31,253,31,79,31,136,31,63,31,146,31,16,31,14,31,83,31,83,30,122,31,122,30,129,31,129,30,30,31,248,31,58,31,58,30,179,31,181,31,116,31,65,31,65,30,65,29,236,31,124,31,209,31,25,31,26,31,26,30,189,31,218,31,185,31,154,31,19,31,13,31,218,31,33,31,33,30,33,29,196,31,78,31,148,31,175,31,175,30,152,31,212,31,212,30,114,31,247,31,167,31,175,31,59,31,154,31,84,31,151,31,141,31,241,31,63,31,224,31,169,31,146,31,40,31,69,31,69,30,47,31,94,31,217,31,196,31,196,30,196,29,146,31,226,31,93,31,121,31,51,31,208,31,117,31,233,31,231,31,231,30,200,31,69,31,70,31,17,31,248,31,113,31,44,31,245,31,221,31,247,31,30,31,48,31,72,31,55,31,55,30,79,31,68,31,227,31,188,31,107,31,116,31,212,31,212,30,88,31,88,30,190,31,79,31,253,31,95,31,107,31,107,30,15,31,15,30,15,29,61,31,74,31,6,31,125,31,171,31,229,31,123,31,100,31,246,31,50,31,50,31,18,31,237,31,77,31,6,31,36,31,36,30,239,31,251,31,199,31,127,31,132,31,53,31,53,30,68,31,68,30,198,31,147,31,167,31,144,31,15,31,221,31,108,31,234,31,234,30,110,31,30,31,121,31,211,31,232,31,22,31,188,31,9,31,60,31,187,31,82,31,139,31,119,31,123,31,123,30,75,31,255,31,110,31,3,31,184,31,82,31,82,30,98,31,45,31,45,30,4,31,2,31,247,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
