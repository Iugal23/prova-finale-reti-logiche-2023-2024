-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 659;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (245,0,251,0,24,0,23,0,88,0,21,0,249,0,184,0,134,0,161,0,111,0,153,0,246,0,169,0,154,0,12,0,126,0,255,0,48,0,144,0,0,0,0,0,162,0,243,0,106,0,152,0,207,0,147,0,0,0,145,0,97,0,0,0,0,0,124,0,28,0,0,0,116,0,253,0,233,0,221,0,144,0,0,0,140,0,242,0,0,0,151,0,204,0,25,0,130,0,105,0,235,0,0,0,0,0,194,0,113,0,169,0,0,0,0,0,69,0,46,0,102,0,0,0,129,0,0,0,0,0,0,0,233,0,178,0,112,0,37,0,146,0,88,0,0,0,0,0,216,0,84,0,0,0,121,0,0,0,68,0,91,0,63,0,0,0,137,0,56,0,254,0,0,0,55,0,119,0,51,0,76,0,208,0,168,0,182,0,159,0,100,0,92,0,84,0,233,0,13,0,80,0,102,0,195,0,6,0,204,0,0,0,14,0,41,0,95,0,0,0,69,0,196,0,144,0,0,0,193,0,84,0,0,0,0,0,187,0,215,0,154,0,116,0,100,0,0,0,0,0,164,0,73,0,84,0,0,0,169,0,174,0,85,0,128,0,0,0,185,0,126,0,0,0,85,0,209,0,0,0,162,0,66,0,0,0,211,0,0,0,65,0,55,0,254,0,250,0,20,0,0,0,225,0,144,0,0,0,187,0,0,0,232,0,11,0,151,0,158,0,0,0,125,0,167,0,193,0,160,0,0,0,170,0,0,0,215,0,242,0,118,0,59,0,14,0,165,0,174,0,190,0,248,0,186,0,85,0,161,0,0,0,154,0,0,0,160,0,35,0,44,0,0,0,187,0,70,0,194,0,190,0,150,0,21,0,241,0,208,0,63,0,247,0,0,0,255,0,0,0,79,0,139,0,199,0,0,0,151,0,244,0,249,0,75,0,0,0,165,0,221,0,147,0,14,0,28,0,252,0,112,0,0,0,248,0,202,0,128,0,169,0,0,0,195,0,89,0,92,0,186,0,211,0,215,0,95,0,130,0,66,0,224,0,66,0,234,0,162,0,0,0,238,0,140,0,250,0,184,0,159,0,227,0,0,0,137,0,79,0,75,0,69,0,244,0,47,0,157,0,0,0,168,0,73,0,173,0,0,0,0,0,0,0,120,0,99,0,0,0,110,0,0,0,0,0,55,0,189,0,154,0,158,0,143,0,0,0,0,0,0,0,135,0,182,0,123,0,172,0,88,0,0,0,89,0,156,0,153,0,243,0,65,0,226,0,38,0,0,0,123,0,231,0,252,0,8,0,0,0,104,0,216,0,78,0,0,0,96,0,141,0,0,0,242,0,213,0,159,0,174,0,147,0,146,0,142,0,142,0,0,0,64,0,216,0,78,0,33,0,0,0,79,0,64,0,56,0,43,0,15,0,17,0,0,0,0,0,223,0,191,0,42,0,193,0,173,0,110,0,231,0,46,0,47,0,80,0,53,0,7,0,239,0,64,0,6,0,31,0,49,0,15,0,0,0,0,0,158,0,97,0,98,0,22,0,107,0,252,0,21,0,255,0,175,0,171,0,125,0,91,0,121,0,68,0,4,0,0,0,239,0,198,0,207,0,0,0,35,0,174,0,0,0,157,0,93,0,0,0,203,0,28,0,238,0,243,0,32,0,3,0,0,0,82,0,194,0,254,0,117,0,76,0,0,0,119,0,45,0,127,0,143,0,146,0,77,0,107,0,111,0,39,0,164,0,229,0,0,0,237,0,96,0,42,0,240,0,167,0,28,0,138,0,0,0,107,0,248,0,12,0,23,0,170,0,124,0,0,0,249,0,70,0,79,0,35,0,0,0,142,0,0,0,0,0,0,0,0,0,73,0,74,0,252,0,47,0,0,0,175,0,0,0,227,0,0,0,0,0,221,0,144,0,56,0,245,0,87,0,0,0,159,0,0,0,138,0,191,0,131,0,13,0,205,0,65,0,0,0,195,0,174,0,38,0,0,0,210,0,227,0,221,0,78,0,131,0,46,0,85,0,33,0,46,0,74,0,146,0,216,0,189,0,96,0,205,0,101,0,0,0,71,0,0,0,58,0,0,0,34,0,0,0,121,0,150,0,84,0,0,0,43,0,14,0,134,0,55,0,218,0,165,0,0,0,74,0,222,0,0,0,155,0,202,0,127,0,217,0,0,0,196,0,246,0,88,0,0,0,121,0,107,0,213,0,0,0,229,0,236,0,173,0,245,0,13,0,0,0,4,0,218,0,134,0,234,0,89,0,131,0,0,0,103,0,41,0,243,0,157,0,29,0,254,0,41,0,210,0,179,0,14,0,213,0,148,0,105,0,0,0,214,0,111,0,206,0,108,0,113,0,0,0,149,0,108,0,0,0,86,0,0,0,0,0,0,0,191,0,0,0,68,0,247,0,99,0,126,0,241,0,19,0,233,0,0,0,0,0,55,0,180,0,48,0,147,0,10,0,0,0,181,0,0,0,18,0,148,0,254,0,74,0,7,0,7,0,112,0,0,0,25,0,0,0,3,0,69,0,91,0,255,0,0,0,108,0,34,0,62,0,0,0,0,0,0,0,191,0,20,0,154,0,35,0,217,0,0,0,202,0,110,0,0,0,65,0,236,0,0,0,213,0,238,0,82,0,103,0,135,0,71,0,55,0,0,0,174,0,231,0,74,0,127,0,105,0,0,0,69,0,227,0,115,0,215,0,243,0,139,0,160,0,0,0,23,0,61,0,137,0,40,0,118,0,193,0,0,0,195,0,0,0,247,0,255,0,0,0,168,0,255,0,0,0,113,0,99,0,82,0,16,0,196,0,238,0,0,0,171,0,241,0,18,0,0,0,23,0,145,0,74,0,89,0,38,0,249,0,0,0,1,0,14,0,0,0,111,0,67,0,0,0,247,0,243,0,167,0,179,0,48,0,156,0,121,0,24,0,205,0,0,0,94,0,0,0);
signal scenario_full  : scenario_type := (245,31,251,31,24,31,23,31,88,31,21,31,249,31,184,31,134,31,161,31,111,31,153,31,246,31,169,31,154,31,12,31,126,31,255,31,48,31,144,31,144,30,144,29,162,31,243,31,106,31,152,31,207,31,147,31,147,30,145,31,97,31,97,30,97,29,124,31,28,31,28,30,116,31,253,31,233,31,221,31,144,31,144,30,140,31,242,31,242,30,151,31,204,31,25,31,130,31,105,31,235,31,235,30,235,29,194,31,113,31,169,31,169,30,169,29,69,31,46,31,102,31,102,30,129,31,129,30,129,29,129,28,233,31,178,31,112,31,37,31,146,31,88,31,88,30,88,29,216,31,84,31,84,30,121,31,121,30,68,31,91,31,63,31,63,30,137,31,56,31,254,31,254,30,55,31,119,31,51,31,76,31,208,31,168,31,182,31,159,31,100,31,92,31,84,31,233,31,13,31,80,31,102,31,195,31,6,31,204,31,204,30,14,31,41,31,95,31,95,30,69,31,196,31,144,31,144,30,193,31,84,31,84,30,84,29,187,31,215,31,154,31,116,31,100,31,100,30,100,29,164,31,73,31,84,31,84,30,169,31,174,31,85,31,128,31,128,30,185,31,126,31,126,30,85,31,209,31,209,30,162,31,66,31,66,30,211,31,211,30,65,31,55,31,254,31,250,31,20,31,20,30,225,31,144,31,144,30,187,31,187,30,232,31,11,31,151,31,158,31,158,30,125,31,167,31,193,31,160,31,160,30,170,31,170,30,215,31,242,31,118,31,59,31,14,31,165,31,174,31,190,31,248,31,186,31,85,31,161,31,161,30,154,31,154,30,160,31,35,31,44,31,44,30,187,31,70,31,194,31,190,31,150,31,21,31,241,31,208,31,63,31,247,31,247,30,255,31,255,30,79,31,139,31,199,31,199,30,151,31,244,31,249,31,75,31,75,30,165,31,221,31,147,31,14,31,28,31,252,31,112,31,112,30,248,31,202,31,128,31,169,31,169,30,195,31,89,31,92,31,186,31,211,31,215,31,95,31,130,31,66,31,224,31,66,31,234,31,162,31,162,30,238,31,140,31,250,31,184,31,159,31,227,31,227,30,137,31,79,31,75,31,69,31,244,31,47,31,157,31,157,30,168,31,73,31,173,31,173,30,173,29,173,28,120,31,99,31,99,30,110,31,110,30,110,29,55,31,189,31,154,31,158,31,143,31,143,30,143,29,143,28,135,31,182,31,123,31,172,31,88,31,88,30,89,31,156,31,153,31,243,31,65,31,226,31,38,31,38,30,123,31,231,31,252,31,8,31,8,30,104,31,216,31,78,31,78,30,96,31,141,31,141,30,242,31,213,31,159,31,174,31,147,31,146,31,142,31,142,31,142,30,64,31,216,31,78,31,33,31,33,30,79,31,64,31,56,31,43,31,15,31,17,31,17,30,17,29,223,31,191,31,42,31,193,31,173,31,110,31,231,31,46,31,47,31,80,31,53,31,7,31,239,31,64,31,6,31,31,31,49,31,15,31,15,30,15,29,158,31,97,31,98,31,22,31,107,31,252,31,21,31,255,31,175,31,171,31,125,31,91,31,121,31,68,31,4,31,4,30,239,31,198,31,207,31,207,30,35,31,174,31,174,30,157,31,93,31,93,30,203,31,28,31,238,31,243,31,32,31,3,31,3,30,82,31,194,31,254,31,117,31,76,31,76,30,119,31,45,31,127,31,143,31,146,31,77,31,107,31,111,31,39,31,164,31,229,31,229,30,237,31,96,31,42,31,240,31,167,31,28,31,138,31,138,30,107,31,248,31,12,31,23,31,170,31,124,31,124,30,249,31,70,31,79,31,35,31,35,30,142,31,142,30,142,29,142,28,142,27,73,31,74,31,252,31,47,31,47,30,175,31,175,30,227,31,227,30,227,29,221,31,144,31,56,31,245,31,87,31,87,30,159,31,159,30,138,31,191,31,131,31,13,31,205,31,65,31,65,30,195,31,174,31,38,31,38,30,210,31,227,31,221,31,78,31,131,31,46,31,85,31,33,31,46,31,74,31,146,31,216,31,189,31,96,31,205,31,101,31,101,30,71,31,71,30,58,31,58,30,34,31,34,30,121,31,150,31,84,31,84,30,43,31,14,31,134,31,55,31,218,31,165,31,165,30,74,31,222,31,222,30,155,31,202,31,127,31,217,31,217,30,196,31,246,31,88,31,88,30,121,31,107,31,213,31,213,30,229,31,236,31,173,31,245,31,13,31,13,30,4,31,218,31,134,31,234,31,89,31,131,31,131,30,103,31,41,31,243,31,157,31,29,31,254,31,41,31,210,31,179,31,14,31,213,31,148,31,105,31,105,30,214,31,111,31,206,31,108,31,113,31,113,30,149,31,108,31,108,30,86,31,86,30,86,29,86,28,191,31,191,30,68,31,247,31,99,31,126,31,241,31,19,31,233,31,233,30,233,29,55,31,180,31,48,31,147,31,10,31,10,30,181,31,181,30,18,31,148,31,254,31,74,31,7,31,7,31,112,31,112,30,25,31,25,30,3,31,69,31,91,31,255,31,255,30,108,31,34,31,62,31,62,30,62,29,62,28,191,31,20,31,154,31,35,31,217,31,217,30,202,31,110,31,110,30,65,31,236,31,236,30,213,31,238,31,82,31,103,31,135,31,71,31,55,31,55,30,174,31,231,31,74,31,127,31,105,31,105,30,69,31,227,31,115,31,215,31,243,31,139,31,160,31,160,30,23,31,61,31,137,31,40,31,118,31,193,31,193,30,195,31,195,30,247,31,255,31,255,30,168,31,255,31,255,30,113,31,99,31,82,31,16,31,196,31,238,31,238,30,171,31,241,31,18,31,18,30,23,31,145,31,74,31,89,31,38,31,249,31,249,30,1,31,14,31,14,30,111,31,67,31,67,30,247,31,243,31,167,31,179,31,48,31,156,31,121,31,24,31,205,31,205,30,94,31,94,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
