-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_28 is
end project_tb_28;

architecture project_tb_arch_28 of project_tb_28 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 180;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,94,0,29,0,169,0,186,0,46,0,174,0,150,0,141,0,144,0,50,0,1,0,0,0,228,0,20,0,0,0,165,0,56,0,158,0,180,0,171,0,76,0,222,0,77,0,70,0,131,0,0,0,134,0,218,0,195,0,188,0,9,0,146,0,45,0,178,0,240,0,49,0,84,0,56,0,205,0,249,0,146,0,0,0,101,0,85,0,42,0,32,0,159,0,55,0,24,0,0,0,0,0,155,0,80,0,0,0,28,0,3,0,0,0,36,0,189,0,87,0,37,0,216,0,9,0,243,0,84,0,49,0,18,0,106,0,16,0,191,0,53,0,185,0,120,0,89,0,226,0,25,0,63,0,226,0,184,0,106,0,49,0,192,0,0,0,205,0,0,0,169,0,19,0,80,0,209,0,102,0,0,0,159,0,71,0,107,0,134,0,2,0,161,0,242,0,179,0,0,0,221,0,136,0,211,0,160,0,235,0,7,0,195,0,50,0,49,0,81,0,0,0,21,0,196,0,0,0,72,0,122,0,15,0,0,0,20,0,16,0,28,0,0,0,183,0,217,0,34,0,196,0,0,0,22,0,0,0,0,0,22,0,255,0,104,0,140,0,0,0,47,0,0,0,54,0,0,0,234,0,0,0,39,0,190,0,193,0,249,0,206,0,101,0,0,0,3,0,117,0,131,0,28,0,233,0,0,0,0,0,230,0,0,0,191,0,65,0,0,0,39,0,88,0,20,0,87,0,244,0,238,0,102,0,135,0,237,0,76,0,0,0,225,0,227,0,3,0,239,0,0,0,9,0,0,0);
signal scenario_full  : scenario_type := (0,0,0,0,94,31,29,31,169,31,186,31,46,31,174,31,150,31,141,31,144,31,50,31,1,31,1,30,228,31,20,31,20,30,165,31,56,31,158,31,180,31,171,31,76,31,222,31,77,31,70,31,131,31,131,30,134,31,218,31,195,31,188,31,9,31,146,31,45,31,178,31,240,31,49,31,84,31,56,31,205,31,249,31,146,31,146,30,101,31,85,31,42,31,32,31,159,31,55,31,24,31,24,30,24,29,155,31,80,31,80,30,28,31,3,31,3,30,36,31,189,31,87,31,37,31,216,31,9,31,243,31,84,31,49,31,18,31,106,31,16,31,191,31,53,31,185,31,120,31,89,31,226,31,25,31,63,31,226,31,184,31,106,31,49,31,192,31,192,30,205,31,205,30,169,31,19,31,80,31,209,31,102,31,102,30,159,31,71,31,107,31,134,31,2,31,161,31,242,31,179,31,179,30,221,31,136,31,211,31,160,31,235,31,7,31,195,31,50,31,49,31,81,31,81,30,21,31,196,31,196,30,72,31,122,31,15,31,15,30,20,31,16,31,28,31,28,30,183,31,217,31,34,31,196,31,196,30,22,31,22,30,22,29,22,31,255,31,104,31,140,31,140,30,47,31,47,30,54,31,54,30,234,31,234,30,39,31,190,31,193,31,249,31,206,31,101,31,101,30,3,31,117,31,131,31,28,31,233,31,233,30,233,29,230,31,230,30,191,31,65,31,65,30,39,31,88,31,20,31,87,31,244,31,238,31,102,31,135,31,237,31,76,31,76,30,225,31,227,31,3,31,239,31,239,30,9,31,9,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
