-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 915;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (186,0,223,0,0,0,240,0,0,0,252,0,220,0,171,0,111,0,36,0,169,0,108,0,175,0,98,0,0,0,15,0,81,0,0,0,120,0,38,0,234,0,176,0,252,0,7,0,0,0,241,0,172,0,112,0,0,0,0,0,83,0,50,0,157,0,197,0,27,0,219,0,229,0,0,0,223,0,125,0,183,0,95,0,71,0,182,0,0,0,45,0,4,0,0,0,173,0,0,0,13,0,16,0,235,0,118,0,0,0,0,0,71,0,76,0,7,0,29,0,11,0,100,0,68,0,43,0,95,0,132,0,83,0,24,0,0,0,233,0,119,0,91,0,199,0,0,0,23,0,0,0,87,0,107,0,192,0,205,0,154,0,59,0,127,0,81,0,0,0,209,0,171,0,251,0,78,0,0,0,0,0,148,0,250,0,153,0,180,0,55,0,123,0,78,0,0,0,180,0,218,0,205,0,48,0,212,0,0,0,17,0,162,0,233,0,213,0,0,0,168,0,129,0,101,0,78,0,148,0,194,0,126,0,249,0,179,0,4,0,0,0,26,0,187,0,89,0,47,0,0,0,132,0,214,0,0,0,83,0,69,0,219,0,60,0,134,0,0,0,63,0,0,0,108,0,0,0,23,0,31,0,52,0,245,0,46,0,37,0,214,0,169,0,199,0,31,0,199,0,42,0,28,0,141,0,131,0,168,0,206,0,32,0,50,0,0,0,0,0,14,0,0,0,43,0,229,0,82,0,206,0,0,0,0,0,0,0,0,0,250,0,51,0,0,0,134,0,0,0,192,0,125,0,174,0,32,0,101,0,0,0,239,0,177,0,118,0,117,0,185,0,0,0,13,0,0,0,0,0,241,0,80,0,92,0,75,0,0,0,32,0,86,0,167,0,166,0,141,0,144,0,131,0,46,0,0,0,0,0,60,0,0,0,13,0,54,0,31,0,47,0,4,0,225,0,0,0,44,0,112,0,80,0,126,0,0,0,95,0,0,0,196,0,63,0,83,0,105,0,145,0,0,0,0,0,0,0,21,0,58,0,31,0,79,0,206,0,151,0,131,0,227,0,0,0,244,0,0,0,0,0,208,0,28,0,151,0,216,0,249,0,120,0,212,0,0,0,169,0,67,0,221,0,241,0,100,0,146,0,18,0,108,0,0,0,0,0,59,0,97,0,11,0,144,0,105,0,23,0,0,0,0,0,207,0,55,0,0,0,0,0,87,0,151,0,63,0,85,0,163,0,252,0,242,0,143,0,13,0,61,0,38,0,106,0,231,0,104,0,34,0,160,0,157,0,5,0,0,0,0,0,149,0,82,0,0,0,29,0,0,0,186,0,70,0,243,0,231,0,0,0,77,0,0,0,232,0,161,0,212,0,249,0,216,0,0,0,1,0,54,0,247,0,99,0,87,0,58,0,214,0,0,0,4,0,213,0,2,0,7,0,162,0,176,0,9,0,244,0,0,0,200,0,0,0,168,0,124,0,0,0,157,0,0,0,90,0,228,0,192,0,200,0,0,0,13,0,18,0,0,0,222,0,247,0,200,0,121,0,239,0,21,0,135,0,125,0,76,0,27,0,0,0,0,0,0,0,104,0,0,0,237,0,193,0,51,0,0,0,17,0,0,0,196,0,0,0,167,0,146,0,174,0,64,0,158,0,95,0,27,0,113,0,150,0,0,0,104,0,157,0,0,0,0,0,48,0,13,0,84,0,180,0,45,0,181,0,80,0,168,0,162,0,214,0,168,0,54,0,81,0,174,0,0,0,105,0,51,0,245,0,0,0,0,0,235,0,75,0,41,0,63,0,177,0,0,0,0,0,213,0,110,0,239,0,177,0,71,0,168,0,206,0,80,0,156,0,14,0,0,0,104,0,0,0,0,0,156,0,0,0,145,0,226,0,163,0,0,0,34,0,5,0,41,0,18,0,127,0,253,0,253,0,147,0,0,0,24,0,213,0,177,0,165,0,129,0,0,0,171,0,35,0,23,0,0,0,56,0,201,0,211,0,14,0,58,0,110,0,104,0,8,0,161,0,0,0,195,0,227,0,110,0,241,0,0,0,85,0,207,0,196,0,108,0,227,0,58,0,125,0,115,0,44,0,44,0,0,0,139,0,248,0,124,0,67,0,79,0,97,0,205,0,178,0,152,0,245,0,27,0,77,0,0,0,129,0,232,0,187,0,134,0,34,0,0,0,45,0,23,0,0,0,203,0,221,0,197,0,93,0,24,0,76,0,173,0,106,0,202,0,247,0,0,0,203,0,120,0,225,0,0,0,64,0,161,0,0,0,153,0,227,0,224,0,165,0,0,0,66,0,221,0,106,0,209,0,40,0,0,0,24,0,27,0,227,0,80,0,247,0,101,0,179,0,116,0,46,0,0,0,63,0,0,0,0,0,92,0,161,0,215,0,157,0,192,0,37,0,8,0,104,0,204,0,137,0,21,0,91,0,228,0,94,0,8,0,170,0,0,0,157,0,188,0,152,0,149,0,139,0,0,0,105,0,0,0,169,0,121,0,47,0,14,0,0,0,184,0,0,0,228,0,89,0,198,0,24,0,203,0,249,0,192,0,206,0,0,0,157,0,244,0,202,0,60,0,28,0,55,0,103,0,83,0,228,0,83,0,44,0,125,0,108,0,0,0,0,0,158,0,0,0,228,0,36,0,83,0,123,0,126,0,47,0,181,0,58,0,8,0,93,0,0,0,187,0,111,0,0,0,221,0,124,0,190,0,149,0,142,0,0,0,214,0,15,0,0,0,152,0,146,0,155,0,0,0,0,0,106,0,49,0,0,0,0,0,0,0,150,0,248,0,82,0,113,0,135,0,0,0,0,0,25,0,214,0,180,0,148,0,49,0,69,0,199,0,218,0,0,0,0,0,191,0,202,0,42,0,120,0,0,0,0,0,175,0,203,0,8,0,0,0,144,0,239,0,0,0,24,0,154,0,0,0,241,0,0,0,5,0,0,0,0,0,110,0,162,0,220,0,51,0,76,0,0,0,103,0,168,0,0,0,243,0,67,0,142,0,242,0,104,0,113,0,0,0,142,0,44,0,166,0,0,0,148,0,124,0,230,0,9,0,175,0,19,0,219,0,29,0,197,0,79,0,0,0,53,0,0,0,25,0,180,0,16,0,97,0,0,0,37,0,101,0,67,0,0,0,0,0,61,0,130,0,106,0,28,0,188,0,193,0,140,0,0,0,129,0,214,0,248,0,0,0,1,0,0,0,158,0,0,0,242,0,124,0,106,0,17,0,151,0,0,0,0,0,168,0,45,0,202,0,125,0,0,0,90,0,0,0,0,0,13,0,119,0,153,0,201,0,117,0,173,0,185,0,196,0,222,0,156,0,95,0,139,0,193,0,68,0,217,0,63,0,71,0,126,0,192,0,157,0,42,0,75,0,209,0,0,0,109,0,0,0,147,0,206,0,112,0,154,0,211,0,57,0,179,0,165,0,0,0,72,0,210,0,100,0,192,0,26,0,51,0,174,0,219,0,165,0,0,0,127,0,232,0,190,0,252,0,131,0,110,0,0,0,159,0,110,0,0,0,105,0,173,0,0,0,0,0,100,0,138,0,0,0,142,0,141,0,78,0,50,0,0,0,171,0,105,0,0,0,8,0,71,0,231,0,0,0,85,0,21,0,0,0,159,0,135,0,119,0,0,0,55,0,171,0,78,0,185,0,240,0,211,0,132,0,101,0,14,0,115,0,0,0,241,0,125,0,73,0,187,0,210,0,97,0,200,0,20,0,0,0,13,0,74,0,0,0,0,0,198,0,165,0,38,0,248,0,133,0,118,0,2,0,229,0,0,0,132,0,251,0,0,0,129,0,152,0,0,0,255,0,90,0,0,0,132,0,23,0,0,0,146,0,0,0,7,0,108,0,201,0,0,0,200,0,93,0,56,0,0,0,46,0,214,0,61,0,161,0,113,0,240,0,121,0,160,0,62,0,24,0,254,0,251,0,62,0,129,0,0,0,97,0,243,0,90,0,22,0,241,0,254,0,106,0,54,0,0,0,225,0,15,0,0,0,106,0,145,0,0,0,51,0,23,0,217,0,23,0,72,0,0,0,154,0,78,0,128,0,0,0,217,0,41,0);
signal scenario_full  : scenario_type := (186,31,223,31,223,30,240,31,240,30,252,31,220,31,171,31,111,31,36,31,169,31,108,31,175,31,98,31,98,30,15,31,81,31,81,30,120,31,38,31,234,31,176,31,252,31,7,31,7,30,241,31,172,31,112,31,112,30,112,29,83,31,50,31,157,31,197,31,27,31,219,31,229,31,229,30,223,31,125,31,183,31,95,31,71,31,182,31,182,30,45,31,4,31,4,30,173,31,173,30,13,31,16,31,235,31,118,31,118,30,118,29,71,31,76,31,7,31,29,31,11,31,100,31,68,31,43,31,95,31,132,31,83,31,24,31,24,30,233,31,119,31,91,31,199,31,199,30,23,31,23,30,87,31,107,31,192,31,205,31,154,31,59,31,127,31,81,31,81,30,209,31,171,31,251,31,78,31,78,30,78,29,148,31,250,31,153,31,180,31,55,31,123,31,78,31,78,30,180,31,218,31,205,31,48,31,212,31,212,30,17,31,162,31,233,31,213,31,213,30,168,31,129,31,101,31,78,31,148,31,194,31,126,31,249,31,179,31,4,31,4,30,26,31,187,31,89,31,47,31,47,30,132,31,214,31,214,30,83,31,69,31,219,31,60,31,134,31,134,30,63,31,63,30,108,31,108,30,23,31,31,31,52,31,245,31,46,31,37,31,214,31,169,31,199,31,31,31,199,31,42,31,28,31,141,31,131,31,168,31,206,31,32,31,50,31,50,30,50,29,14,31,14,30,43,31,229,31,82,31,206,31,206,30,206,29,206,28,206,27,250,31,51,31,51,30,134,31,134,30,192,31,125,31,174,31,32,31,101,31,101,30,239,31,177,31,118,31,117,31,185,31,185,30,13,31,13,30,13,29,241,31,80,31,92,31,75,31,75,30,32,31,86,31,167,31,166,31,141,31,144,31,131,31,46,31,46,30,46,29,60,31,60,30,13,31,54,31,31,31,47,31,4,31,225,31,225,30,44,31,112,31,80,31,126,31,126,30,95,31,95,30,196,31,63,31,83,31,105,31,145,31,145,30,145,29,145,28,21,31,58,31,31,31,79,31,206,31,151,31,131,31,227,31,227,30,244,31,244,30,244,29,208,31,28,31,151,31,216,31,249,31,120,31,212,31,212,30,169,31,67,31,221,31,241,31,100,31,146,31,18,31,108,31,108,30,108,29,59,31,97,31,11,31,144,31,105,31,23,31,23,30,23,29,207,31,55,31,55,30,55,29,87,31,151,31,63,31,85,31,163,31,252,31,242,31,143,31,13,31,61,31,38,31,106,31,231,31,104,31,34,31,160,31,157,31,5,31,5,30,5,29,149,31,82,31,82,30,29,31,29,30,186,31,70,31,243,31,231,31,231,30,77,31,77,30,232,31,161,31,212,31,249,31,216,31,216,30,1,31,54,31,247,31,99,31,87,31,58,31,214,31,214,30,4,31,213,31,2,31,7,31,162,31,176,31,9,31,244,31,244,30,200,31,200,30,168,31,124,31,124,30,157,31,157,30,90,31,228,31,192,31,200,31,200,30,13,31,18,31,18,30,222,31,247,31,200,31,121,31,239,31,21,31,135,31,125,31,76,31,27,31,27,30,27,29,27,28,104,31,104,30,237,31,193,31,51,31,51,30,17,31,17,30,196,31,196,30,167,31,146,31,174,31,64,31,158,31,95,31,27,31,113,31,150,31,150,30,104,31,157,31,157,30,157,29,48,31,13,31,84,31,180,31,45,31,181,31,80,31,168,31,162,31,214,31,168,31,54,31,81,31,174,31,174,30,105,31,51,31,245,31,245,30,245,29,235,31,75,31,41,31,63,31,177,31,177,30,177,29,213,31,110,31,239,31,177,31,71,31,168,31,206,31,80,31,156,31,14,31,14,30,104,31,104,30,104,29,156,31,156,30,145,31,226,31,163,31,163,30,34,31,5,31,41,31,18,31,127,31,253,31,253,31,147,31,147,30,24,31,213,31,177,31,165,31,129,31,129,30,171,31,35,31,23,31,23,30,56,31,201,31,211,31,14,31,58,31,110,31,104,31,8,31,161,31,161,30,195,31,227,31,110,31,241,31,241,30,85,31,207,31,196,31,108,31,227,31,58,31,125,31,115,31,44,31,44,31,44,30,139,31,248,31,124,31,67,31,79,31,97,31,205,31,178,31,152,31,245,31,27,31,77,31,77,30,129,31,232,31,187,31,134,31,34,31,34,30,45,31,23,31,23,30,203,31,221,31,197,31,93,31,24,31,76,31,173,31,106,31,202,31,247,31,247,30,203,31,120,31,225,31,225,30,64,31,161,31,161,30,153,31,227,31,224,31,165,31,165,30,66,31,221,31,106,31,209,31,40,31,40,30,24,31,27,31,227,31,80,31,247,31,101,31,179,31,116,31,46,31,46,30,63,31,63,30,63,29,92,31,161,31,215,31,157,31,192,31,37,31,8,31,104,31,204,31,137,31,21,31,91,31,228,31,94,31,8,31,170,31,170,30,157,31,188,31,152,31,149,31,139,31,139,30,105,31,105,30,169,31,121,31,47,31,14,31,14,30,184,31,184,30,228,31,89,31,198,31,24,31,203,31,249,31,192,31,206,31,206,30,157,31,244,31,202,31,60,31,28,31,55,31,103,31,83,31,228,31,83,31,44,31,125,31,108,31,108,30,108,29,158,31,158,30,228,31,36,31,83,31,123,31,126,31,47,31,181,31,58,31,8,31,93,31,93,30,187,31,111,31,111,30,221,31,124,31,190,31,149,31,142,31,142,30,214,31,15,31,15,30,152,31,146,31,155,31,155,30,155,29,106,31,49,31,49,30,49,29,49,28,150,31,248,31,82,31,113,31,135,31,135,30,135,29,25,31,214,31,180,31,148,31,49,31,69,31,199,31,218,31,218,30,218,29,191,31,202,31,42,31,120,31,120,30,120,29,175,31,203,31,8,31,8,30,144,31,239,31,239,30,24,31,154,31,154,30,241,31,241,30,5,31,5,30,5,29,110,31,162,31,220,31,51,31,76,31,76,30,103,31,168,31,168,30,243,31,67,31,142,31,242,31,104,31,113,31,113,30,142,31,44,31,166,31,166,30,148,31,124,31,230,31,9,31,175,31,19,31,219,31,29,31,197,31,79,31,79,30,53,31,53,30,25,31,180,31,16,31,97,31,97,30,37,31,101,31,67,31,67,30,67,29,61,31,130,31,106,31,28,31,188,31,193,31,140,31,140,30,129,31,214,31,248,31,248,30,1,31,1,30,158,31,158,30,242,31,124,31,106,31,17,31,151,31,151,30,151,29,168,31,45,31,202,31,125,31,125,30,90,31,90,30,90,29,13,31,119,31,153,31,201,31,117,31,173,31,185,31,196,31,222,31,156,31,95,31,139,31,193,31,68,31,217,31,63,31,71,31,126,31,192,31,157,31,42,31,75,31,209,31,209,30,109,31,109,30,147,31,206,31,112,31,154,31,211,31,57,31,179,31,165,31,165,30,72,31,210,31,100,31,192,31,26,31,51,31,174,31,219,31,165,31,165,30,127,31,232,31,190,31,252,31,131,31,110,31,110,30,159,31,110,31,110,30,105,31,173,31,173,30,173,29,100,31,138,31,138,30,142,31,141,31,78,31,50,31,50,30,171,31,105,31,105,30,8,31,71,31,231,31,231,30,85,31,21,31,21,30,159,31,135,31,119,31,119,30,55,31,171,31,78,31,185,31,240,31,211,31,132,31,101,31,14,31,115,31,115,30,241,31,125,31,73,31,187,31,210,31,97,31,200,31,20,31,20,30,13,31,74,31,74,30,74,29,198,31,165,31,38,31,248,31,133,31,118,31,2,31,229,31,229,30,132,31,251,31,251,30,129,31,152,31,152,30,255,31,90,31,90,30,132,31,23,31,23,30,146,31,146,30,7,31,108,31,201,31,201,30,200,31,93,31,56,31,56,30,46,31,214,31,61,31,161,31,113,31,240,31,121,31,160,31,62,31,24,31,254,31,251,31,62,31,129,31,129,30,97,31,243,31,90,31,22,31,241,31,254,31,106,31,54,31,54,30,225,31,15,31,15,30,106,31,145,31,145,30,51,31,23,31,217,31,23,31,72,31,72,30,154,31,78,31,128,31,128,30,217,31,41,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
