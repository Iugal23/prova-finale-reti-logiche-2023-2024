-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 644;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (8,0,0,0,29,0,64,0,106,0,20,0,0,0,228,0,70,0,34,0,168,0,41,0,122,0,0,0,88,0,17,0,0,0,49,0,72,0,136,0,2,0,211,0,225,0,133,0,0,0,73,0,54,0,238,0,129,0,90,0,113,0,148,0,81,0,0,0,175,0,34,0,203,0,25,0,22,0,0,0,124,0,0,0,210,0,68,0,139,0,0,0,227,0,45,0,70,0,0,0,57,0,0,0,94,0,0,0,0,0,98,0,147,0,210,0,141,0,87,0,190,0,211,0,0,0,0,0,232,0,113,0,8,0,0,0,0,0,129,0,176,0,243,0,241,0,218,0,49,0,153,0,176,0,23,0,171,0,0,0,122,0,49,0,62,0,143,0,214,0,220,0,118,0,157,0,38,0,208,0,181,0,56,0,204,0,99,0,0,0,188,0,209,0,193,0,137,0,249,0,168,0,205,0,224,0,156,0,122,0,144,0,3,0,222,0,79,0,239,0,20,0,177,0,107,0,127,0,193,0,145,0,3,0,116,0,222,0,54,0,171,0,20,0,242,0,201,0,10,0,225,0,217,0,87,0,28,0,210,0,109,0,107,0,105,0,97,0,0,0,219,0,105,0,46,0,77,0,198,0,0,0,91,0,193,0,32,0,251,0,241,0,0,0,0,0,0,0,0,0,59,0,184,0,172,0,118,0,126,0,11,0,0,0,120,0,218,0,78,0,0,0,105,0,230,0,223,0,25,0,0,0,209,0,0,0,209,0,0,0,185,0,170,0,173,0,97,0,113,0,13,0,0,0,75,0,212,0,169,0,20,0,100,0,63,0,57,0,82,0,156,0,136,0,105,0,192,0,141,0,204,0,0,0,0,0,32,0,148,0,0,0,87,0,31,0,213,0,84,0,0,0,0,0,35,0,8,0,200,0,80,0,216,0,155,0,221,0,197,0,74,0,164,0,0,0,188,0,18,0,216,0,223,0,170,0,162,0,82,0,0,0,217,0,121,0,236,0,2,0,11,0,50,0,187,0,58,0,0,0,0,0,165,0,232,0,0,0,51,0,128,0,0,0,0,0,17,0,0,0,158,0,75,0,2,0,175,0,189,0,123,0,0,0,0,0,0,0,181,0,4,0,0,0,162,0,3,0,0,0,86,0,133,0,0,0,3,0,58,0,52,0,223,0,235,0,214,0,0,0,110,0,81,0,210,0,37,0,0,0,208,0,0,0,170,0,0,0,7,0,195,0,206,0,0,0,218,0,0,0,24,0,109,0,217,0,0,0,95,0,13,0,80,0,0,0,0,0,137,0,102,0,128,0,20,0,0,0,0,0,68,0,108,0,0,0,66,0,15,0,0,0,131,0,166,0,103,0,180,0,238,0,165,0,187,0,96,0,0,0,133,0,8,0,125,0,0,0,0,0,93,0,0,0,0,0,0,0,57,0,181,0,113,0,238,0,244,0,20,0,2,0,89,0,208,0,23,0,0,0,111,0,213,0,230,0,0,0,0,0,226,0,180,0,241,0,72,0,0,0,0,0,23,0,210,0,235,0,223,0,98,0,146,0,0,0,216,0,91,0,148,0,91,0,100,0,237,0,0,0,130,0,75,0,0,0,0,0,0,0,204,0,33,0,11,0,10,0,162,0,166,0,142,0,89,0,19,0,128,0,34,0,224,0,199,0,181,0,146,0,50,0,180,0,1,0,52,0,223,0,0,0,219,0,113,0,207,0,76,0,146,0,245,0,140,0,49,0,0,0,0,0,60,0,0,0,0,0,0,0,20,0,31,0,39,0,239,0,136,0,4,0,232,0,58,0,203,0,133,0,210,0,180,0,0,0,86,0,0,0,97,0,230,0,26,0,0,0,141,0,199,0,98,0,93,0,41,0,185,0,174,0,0,0,255,0,157,0,75,0,24,0,197,0,37,0,228,0,91,0,58,0,255,0,249,0,183,0,31,0,0,0,167,0,218,0,103,0,0,0,229,0,16,0,6,0,233,0,93,0,147,0,218,0,0,0,57,0,0,0,0,0,70,0,187,0,102,0,249,0,77,0,50,0,94,0,142,0,214,0,142,0,27,0,132,0,0,0,45,0,0,0,212,0,215,0,0,0,226,0,49,0,191,0,0,0,186,0,81,0,73,0,67,0,91,0,0,0,10,0,90,0,0,0,233,0,29,0,137,0,23,0,185,0,196,0,223,0,99,0,216,0,44,0,236,0,77,0,170,0,214,0,215,0,98,0,0,0,156,0,28,0,0,0,70,0,236,0,72,0,174,0,38,0,83,0,6,0,116,0,208,0,108,0,23,0,76,0,88,0,0,0,33,0,0,0,138,0,0,0,117,0,105,0,0,0,0,0,193,0,168,0,56,0,190,0,240,0,213,0,159,0,0,0,27,0,0,0,192,0,0,0,0,0,72,0,182,0,113,0,52,0,112,0,245,0,146,0,12,0,162,0,25,0,226,0,77,0,145,0,245,0,13,0,0,0,0,0,0,0,128,0,181,0,67,0,159,0,224,0,175,0,31,0,167,0,101,0,0,0,94,0,7,0,195,0,75,0,120,0,119,0,14,0,10,0,0,0,25,0,0,0,0,0,48,0,229,0,158,0,0,0,241,0,7,0,90,0,0,0,36,0,47,0,248,0,226,0,211,0,228,0,124,0,55,0,68,0,0,0,48,0,100,0,0,0,71,0,75,0,93,0,107,0,125,0,0,0,155,0,82,0,0,0,126,0,0,0,158,0,132,0,209,0,220,0,0,0,130,0,200,0,208,0,248,0,187,0,0,0,225,0,194,0,56,0,233,0,0,0,96,0,0,0,216,0,251,0,0,0,88,0,165,0,0,0,151,0,0,0,0,0,113,0,112,0,153,0,19,0,0,0,6,0,119,0,41,0);
signal scenario_full  : scenario_type := (8,31,8,30,29,31,64,31,106,31,20,31,20,30,228,31,70,31,34,31,168,31,41,31,122,31,122,30,88,31,17,31,17,30,49,31,72,31,136,31,2,31,211,31,225,31,133,31,133,30,73,31,54,31,238,31,129,31,90,31,113,31,148,31,81,31,81,30,175,31,34,31,203,31,25,31,22,31,22,30,124,31,124,30,210,31,68,31,139,31,139,30,227,31,45,31,70,31,70,30,57,31,57,30,94,31,94,30,94,29,98,31,147,31,210,31,141,31,87,31,190,31,211,31,211,30,211,29,232,31,113,31,8,31,8,30,8,29,129,31,176,31,243,31,241,31,218,31,49,31,153,31,176,31,23,31,171,31,171,30,122,31,49,31,62,31,143,31,214,31,220,31,118,31,157,31,38,31,208,31,181,31,56,31,204,31,99,31,99,30,188,31,209,31,193,31,137,31,249,31,168,31,205,31,224,31,156,31,122,31,144,31,3,31,222,31,79,31,239,31,20,31,177,31,107,31,127,31,193,31,145,31,3,31,116,31,222,31,54,31,171,31,20,31,242,31,201,31,10,31,225,31,217,31,87,31,28,31,210,31,109,31,107,31,105,31,97,31,97,30,219,31,105,31,46,31,77,31,198,31,198,30,91,31,193,31,32,31,251,31,241,31,241,30,241,29,241,28,241,27,59,31,184,31,172,31,118,31,126,31,11,31,11,30,120,31,218,31,78,31,78,30,105,31,230,31,223,31,25,31,25,30,209,31,209,30,209,31,209,30,185,31,170,31,173,31,97,31,113,31,13,31,13,30,75,31,212,31,169,31,20,31,100,31,63,31,57,31,82,31,156,31,136,31,105,31,192,31,141,31,204,31,204,30,204,29,32,31,148,31,148,30,87,31,31,31,213,31,84,31,84,30,84,29,35,31,8,31,200,31,80,31,216,31,155,31,221,31,197,31,74,31,164,31,164,30,188,31,18,31,216,31,223,31,170,31,162,31,82,31,82,30,217,31,121,31,236,31,2,31,11,31,50,31,187,31,58,31,58,30,58,29,165,31,232,31,232,30,51,31,128,31,128,30,128,29,17,31,17,30,158,31,75,31,2,31,175,31,189,31,123,31,123,30,123,29,123,28,181,31,4,31,4,30,162,31,3,31,3,30,86,31,133,31,133,30,3,31,58,31,52,31,223,31,235,31,214,31,214,30,110,31,81,31,210,31,37,31,37,30,208,31,208,30,170,31,170,30,7,31,195,31,206,31,206,30,218,31,218,30,24,31,109,31,217,31,217,30,95,31,13,31,80,31,80,30,80,29,137,31,102,31,128,31,20,31,20,30,20,29,68,31,108,31,108,30,66,31,15,31,15,30,131,31,166,31,103,31,180,31,238,31,165,31,187,31,96,31,96,30,133,31,8,31,125,31,125,30,125,29,93,31,93,30,93,29,93,28,57,31,181,31,113,31,238,31,244,31,20,31,2,31,89,31,208,31,23,31,23,30,111,31,213,31,230,31,230,30,230,29,226,31,180,31,241,31,72,31,72,30,72,29,23,31,210,31,235,31,223,31,98,31,146,31,146,30,216,31,91,31,148,31,91,31,100,31,237,31,237,30,130,31,75,31,75,30,75,29,75,28,204,31,33,31,11,31,10,31,162,31,166,31,142,31,89,31,19,31,128,31,34,31,224,31,199,31,181,31,146,31,50,31,180,31,1,31,52,31,223,31,223,30,219,31,113,31,207,31,76,31,146,31,245,31,140,31,49,31,49,30,49,29,60,31,60,30,60,29,60,28,20,31,31,31,39,31,239,31,136,31,4,31,232,31,58,31,203,31,133,31,210,31,180,31,180,30,86,31,86,30,97,31,230,31,26,31,26,30,141,31,199,31,98,31,93,31,41,31,185,31,174,31,174,30,255,31,157,31,75,31,24,31,197,31,37,31,228,31,91,31,58,31,255,31,249,31,183,31,31,31,31,30,167,31,218,31,103,31,103,30,229,31,16,31,6,31,233,31,93,31,147,31,218,31,218,30,57,31,57,30,57,29,70,31,187,31,102,31,249,31,77,31,50,31,94,31,142,31,214,31,142,31,27,31,132,31,132,30,45,31,45,30,212,31,215,31,215,30,226,31,49,31,191,31,191,30,186,31,81,31,73,31,67,31,91,31,91,30,10,31,90,31,90,30,233,31,29,31,137,31,23,31,185,31,196,31,223,31,99,31,216,31,44,31,236,31,77,31,170,31,214,31,215,31,98,31,98,30,156,31,28,31,28,30,70,31,236,31,72,31,174,31,38,31,83,31,6,31,116,31,208,31,108,31,23,31,76,31,88,31,88,30,33,31,33,30,138,31,138,30,117,31,105,31,105,30,105,29,193,31,168,31,56,31,190,31,240,31,213,31,159,31,159,30,27,31,27,30,192,31,192,30,192,29,72,31,182,31,113,31,52,31,112,31,245,31,146,31,12,31,162,31,25,31,226,31,77,31,145,31,245,31,13,31,13,30,13,29,13,28,128,31,181,31,67,31,159,31,224,31,175,31,31,31,167,31,101,31,101,30,94,31,7,31,195,31,75,31,120,31,119,31,14,31,10,31,10,30,25,31,25,30,25,29,48,31,229,31,158,31,158,30,241,31,7,31,90,31,90,30,36,31,47,31,248,31,226,31,211,31,228,31,124,31,55,31,68,31,68,30,48,31,100,31,100,30,71,31,75,31,93,31,107,31,125,31,125,30,155,31,82,31,82,30,126,31,126,30,158,31,132,31,209,31,220,31,220,30,130,31,200,31,208,31,248,31,187,31,187,30,225,31,194,31,56,31,233,31,233,30,96,31,96,30,216,31,251,31,251,30,88,31,165,31,165,30,151,31,151,30,151,29,113,31,112,31,153,31,19,31,19,30,6,31,119,31,41,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
