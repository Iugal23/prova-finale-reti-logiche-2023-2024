-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_334 is
end project_tb_334;

architecture project_tb_arch_334 of project_tb_334 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 214;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (109,0,213,0,186,0,251,0,0,0,232,0,182,0,69,0,45,0,213,0,124,0,173,0,160,0,87,0,35,0,249,0,167,0,69,0,115,0,206,0,0,0,8,0,0,0,252,0,59,0,0,0,91,0,237,0,138,0,0,0,0,0,245,0,168,0,218,0,170,0,0,0,152,0,169,0,154,0,211,0,255,0,0,0,0,0,102,0,183,0,0,0,119,0,0,0,184,0,19,0,97,0,180,0,129,0,117,0,0,0,153,0,0,0,0,0,0,0,234,0,100,0,197,0,69,0,0,0,149,0,11,0,127,0,220,0,107,0,0,0,68,0,17,0,0,0,0,0,202,0,125,0,252,0,247,0,0,0,199,0,34,0,94,0,193,0,211,0,198,0,29,0,233,0,57,0,0,0,67,0,214,0,31,0,147,0,205,0,151,0,60,0,246,0,0,0,92,0,212,0,55,0,0,0,240,0,149,0,211,0,232,0,206,0,24,0,112,0,12,0,67,0,216,0,235,0,252,0,178,0,14,0,94,0,96,0,204,0,0,0,32,0,131,0,105,0,169,0,118,0,61,0,115,0,232,0,49,0,215,0,0,0,114,0,113,0,54,0,64,0,213,0,168,0,0,0,143,0,224,0,14,0,83,0,98,0,246,0,0,0,224,0,185,0,214,0,118,0,0,0,77,0,151,0,143,0,0,0,234,0,1,0,247,0,154,0,214,0,0,0,26,0,153,0,43,0,253,0,5,0,0,0,235,0,162,0,123,0,217,0,128,0,0,0,17,0,0,0,57,0,74,0,112,0,120,0,215,0,0,0,168,0,0,0,209,0,216,0,0,0,176,0,45,0,30,0,71,0,30,0,225,0,195,0,246,0,83,0,226,0,13,0,0,0,16,0,0,0,250,0,237,0,221,0,0,0,7,0,27,0,206,0,0,0,101,0,0,0,48,0,224,0,104,0,87,0,0,0);
signal scenario_full  : scenario_type := (109,31,213,31,186,31,251,31,251,30,232,31,182,31,69,31,45,31,213,31,124,31,173,31,160,31,87,31,35,31,249,31,167,31,69,31,115,31,206,31,206,30,8,31,8,30,252,31,59,31,59,30,91,31,237,31,138,31,138,30,138,29,245,31,168,31,218,31,170,31,170,30,152,31,169,31,154,31,211,31,255,31,255,30,255,29,102,31,183,31,183,30,119,31,119,30,184,31,19,31,97,31,180,31,129,31,117,31,117,30,153,31,153,30,153,29,153,28,234,31,100,31,197,31,69,31,69,30,149,31,11,31,127,31,220,31,107,31,107,30,68,31,17,31,17,30,17,29,202,31,125,31,252,31,247,31,247,30,199,31,34,31,94,31,193,31,211,31,198,31,29,31,233,31,57,31,57,30,67,31,214,31,31,31,147,31,205,31,151,31,60,31,246,31,246,30,92,31,212,31,55,31,55,30,240,31,149,31,211,31,232,31,206,31,24,31,112,31,12,31,67,31,216,31,235,31,252,31,178,31,14,31,94,31,96,31,204,31,204,30,32,31,131,31,105,31,169,31,118,31,61,31,115,31,232,31,49,31,215,31,215,30,114,31,113,31,54,31,64,31,213,31,168,31,168,30,143,31,224,31,14,31,83,31,98,31,246,31,246,30,224,31,185,31,214,31,118,31,118,30,77,31,151,31,143,31,143,30,234,31,1,31,247,31,154,31,214,31,214,30,26,31,153,31,43,31,253,31,5,31,5,30,235,31,162,31,123,31,217,31,128,31,128,30,17,31,17,30,57,31,74,31,112,31,120,31,215,31,215,30,168,31,168,30,209,31,216,31,216,30,176,31,45,31,30,31,71,31,30,31,225,31,195,31,246,31,83,31,226,31,13,31,13,30,16,31,16,30,250,31,237,31,221,31,221,30,7,31,27,31,206,31,206,30,101,31,101,30,48,31,224,31,104,31,87,31,87,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
