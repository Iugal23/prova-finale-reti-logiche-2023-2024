-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 397;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,138,0,10,0,0,0,0,0,2,0,101,0,214,0,0,0,192,0,40,0,120,0,0,0,141,0,0,0,0,0,22,0,230,0,173,0,29,0,134,0,46,0,0,0,149,0,0,0,194,0,252,0,185,0,149,0,6,0,248,0,56,0,249,0,0,0,0,0,181,0,15,0,0,0,0,0,0,0,137,0,37,0,230,0,172,0,0,0,0,0,204,0,126,0,246,0,0,0,91,0,72,0,62,0,73,0,8,0,65,0,199,0,99,0,0,0,0,0,39,0,0,0,141,0,54,0,62,0,0,0,0,0,23,0,217,0,224,0,153,0,0,0,114,0,0,0,24,0,39,0,2,0,87,0,45,0,155,0,0,0,0,0,0,0,110,0,189,0,91,0,0,0,97,0,195,0,50,0,87,0,158,0,230,0,222,0,35,0,251,0,145,0,141,0,50,0,250,0,0,0,0,0,3,0,204,0,207,0,0,0,4,0,12,0,173,0,114,0,119,0,236,0,126,0,0,0,203,0,25,0,0,0,19,0,228,0,0,0,0,0,215,0,100,0,224,0,103,0,165,0,0,0,150,0,6,0,0,0,208,0,51,0,141,0,144,0,159,0,0,0,0,0,205,0,6,0,98,0,0,0,69,0,198,0,0,0,0,0,242,0,0,0,193,0,203,0,0,0,45,0,235,0,129,0,128,0,170,0,147,0,0,0,180,0,155,0,0,0,194,0,200,0,23,0,202,0,178,0,57,0,211,0,231,0,3,0,0,0,59,0,245,0,102,0,11,0,136,0,216,0,193,0,78,0,0,0,177,0,249,0,56,0,7,0,83,0,40,0,53,0,29,0,238,0,21,0,0,0,0,0,207,0,238,0,184,0,201,0,0,0,107,0,166,0,180,0,43,0,97,0,21,0,161,0,0,0,54,0,156,0,56,0,208,0,0,0,0,0,235,0,238,0,196,0,31,0,197,0,224,0,0,0,0,0,240,0,0,0,51,0,129,0,81,0,85,0,0,0,0,0,0,0,236,0,113,0,182,0,142,0,17,0,182,0,177,0,25,0,65,0,176,0,159,0,67,0,33,0,0,0,17,0,0,0,0,0,72,0,94,0,148,0,149,0,206,0,27,0,2,0,0,0,70,0,52,0,99,0,248,0,56,0,101,0,149,0,120,0,155,0,231,0,103,0,231,0,130,0,0,0,34,0,0,0,0,0,0,0,34,0,0,0,237,0,69,0,12,0,207,0,250,0,109,0,227,0,153,0,219,0,126,0,213,0,0,0,159,0,225,0,162,0,113,0,106,0,0,0,52,0,204,0,198,0,23,0,135,0,0,0,96,0,224,0,249,0,92,0,204,0,239,0,60,0,0,0,196,0,59,0,255,0,8,0,0,0,147,0,0,0,26,0,162,0,202,0,156,0,0,0,10,0,150,0,121,0,0,0,118,0,3,0,0,0,0,0,30,0,43,0,173,0,0,0,8,0,0,0,25,0,119,0,54,0,173,0,109,0,182,0,174,0,102,0,0,0,24,0,0,0,0,0,0,0,128,0,217,0,78,0,78,0,0,0,16,0,234,0,0,0,0,0,155,0,31,0,64,0,73,0,245,0,33,0,142,0,45,0,128,0,27,0,150,0,212,0,146,0,167,0,49,0,248,0,210,0,58,0,0,0,95,0,219,0,143,0,125,0,197,0,89,0,123,0,108,0,88,0,197,0,116,0,36,0,110,0,106,0,19,0,83,0,191,0,198,0,55,0,129,0,117,0,0,0,166,0,245,0,254,0,147,0);
signal scenario_full  : scenario_type := (0,0,138,31,10,31,10,30,10,29,2,31,101,31,214,31,214,30,192,31,40,31,120,31,120,30,141,31,141,30,141,29,22,31,230,31,173,31,29,31,134,31,46,31,46,30,149,31,149,30,194,31,252,31,185,31,149,31,6,31,248,31,56,31,249,31,249,30,249,29,181,31,15,31,15,30,15,29,15,28,137,31,37,31,230,31,172,31,172,30,172,29,204,31,126,31,246,31,246,30,91,31,72,31,62,31,73,31,8,31,65,31,199,31,99,31,99,30,99,29,39,31,39,30,141,31,54,31,62,31,62,30,62,29,23,31,217,31,224,31,153,31,153,30,114,31,114,30,24,31,39,31,2,31,87,31,45,31,155,31,155,30,155,29,155,28,110,31,189,31,91,31,91,30,97,31,195,31,50,31,87,31,158,31,230,31,222,31,35,31,251,31,145,31,141,31,50,31,250,31,250,30,250,29,3,31,204,31,207,31,207,30,4,31,12,31,173,31,114,31,119,31,236,31,126,31,126,30,203,31,25,31,25,30,19,31,228,31,228,30,228,29,215,31,100,31,224,31,103,31,165,31,165,30,150,31,6,31,6,30,208,31,51,31,141,31,144,31,159,31,159,30,159,29,205,31,6,31,98,31,98,30,69,31,198,31,198,30,198,29,242,31,242,30,193,31,203,31,203,30,45,31,235,31,129,31,128,31,170,31,147,31,147,30,180,31,155,31,155,30,194,31,200,31,23,31,202,31,178,31,57,31,211,31,231,31,3,31,3,30,59,31,245,31,102,31,11,31,136,31,216,31,193,31,78,31,78,30,177,31,249,31,56,31,7,31,83,31,40,31,53,31,29,31,238,31,21,31,21,30,21,29,207,31,238,31,184,31,201,31,201,30,107,31,166,31,180,31,43,31,97,31,21,31,161,31,161,30,54,31,156,31,56,31,208,31,208,30,208,29,235,31,238,31,196,31,31,31,197,31,224,31,224,30,224,29,240,31,240,30,51,31,129,31,81,31,85,31,85,30,85,29,85,28,236,31,113,31,182,31,142,31,17,31,182,31,177,31,25,31,65,31,176,31,159,31,67,31,33,31,33,30,17,31,17,30,17,29,72,31,94,31,148,31,149,31,206,31,27,31,2,31,2,30,70,31,52,31,99,31,248,31,56,31,101,31,149,31,120,31,155,31,231,31,103,31,231,31,130,31,130,30,34,31,34,30,34,29,34,28,34,31,34,30,237,31,69,31,12,31,207,31,250,31,109,31,227,31,153,31,219,31,126,31,213,31,213,30,159,31,225,31,162,31,113,31,106,31,106,30,52,31,204,31,198,31,23,31,135,31,135,30,96,31,224,31,249,31,92,31,204,31,239,31,60,31,60,30,196,31,59,31,255,31,8,31,8,30,147,31,147,30,26,31,162,31,202,31,156,31,156,30,10,31,150,31,121,31,121,30,118,31,3,31,3,30,3,29,30,31,43,31,173,31,173,30,8,31,8,30,25,31,119,31,54,31,173,31,109,31,182,31,174,31,102,31,102,30,24,31,24,30,24,29,24,28,128,31,217,31,78,31,78,31,78,30,16,31,234,31,234,30,234,29,155,31,31,31,64,31,73,31,245,31,33,31,142,31,45,31,128,31,27,31,150,31,212,31,146,31,167,31,49,31,248,31,210,31,58,31,58,30,95,31,219,31,143,31,125,31,197,31,89,31,123,31,108,31,88,31,197,31,116,31,36,31,110,31,106,31,19,31,83,31,191,31,198,31,55,31,129,31,117,31,117,30,166,31,245,31,254,31,147,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
