-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 877;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (83,0,79,0,0,0,15,0,109,0,60,0,0,0,0,0,218,0,116,0,242,0,203,0,0,0,212,0,7,0,157,0,0,0,237,0,130,0,89,0,118,0,212,0,130,0,50,0,188,0,136,0,0,0,146,0,0,0,178,0,73,0,0,0,87,0,255,0,183,0,123,0,66,0,194,0,181,0,124,0,122,0,201,0,0,0,0,0,109,0,46,0,89,0,2,0,134,0,59,0,0,0,127,0,4,0,213,0,5,0,231,0,59,0,9,0,48,0,198,0,215,0,208,0,253,0,139,0,0,0,252,0,5,0,233,0,228,0,124,0,172,0,62,0,7,0,113,0,44,0,25,0,9,0,229,0,135,0,177,0,92,0,54,0,189,0,205,0,178,0,0,0,239,0,20,0,137,0,169,0,162,0,249,0,55,0,209,0,134,0,0,0,211,0,126,0,216,0,101,0,37,0,150,0,182,0,211,0,0,0,232,0,232,0,102,0,232,0,0,0,75,0,0,0,106,0,243,0,47,0,0,0,157,0,12,0,97,0,71,0,119,0,55,0,125,0,145,0,60,0,0,0,157,0,125,0,215,0,50,0,210,0,56,0,0,0,204,0,95,0,105,0,13,0,223,0,0,0,35,0,184,0,0,0,72,0,222,0,0,0,0,0,71,0,52,0,0,0,117,0,83,0,0,0,144,0,250,0,60,0,0,0,139,0,131,0,79,0,97,0,0,0,248,0,219,0,182,0,59,0,223,0,140,0,0,0,49,0,65,0,0,0,80,0,106,0,107,0,20,0,138,0,185,0,109,0,240,0,4,0,33,0,157,0,220,0,0,0,59,0,86,0,0,0,44,0,191,0,227,0,56,0,0,0,89,0,150,0,177,0,0,0,240,0,221,0,206,0,130,0,60,0,241,0,22,0,241,0,0,0,178,0,84,0,74,0,27,0,0,0,72,0,132,0,0,0,157,0,243,0,0,0,11,0,204,0,228,0,199,0,33,0,0,0,143,0,0,0,10,0,225,0,189,0,119,0,0,0,239,0,148,0,188,0,130,0,110,0,245,0,0,0,19,0,31,0,0,0,37,0,117,0,129,0,23,0,154,0,0,0,46,0,72,0,0,0,153,0,201,0,224,0,13,0,0,0,218,0,4,0,140,0,0,0,5,0,0,0,239,0,10,0,74,0,0,0,5,0,128,0,76,0,0,0,135,0,130,0,0,0,255,0,25,0,7,0,65,0,157,0,0,0,90,0,157,0,121,0,182,0,249,0,0,0,152,0,185,0,107,0,124,0,164,0,183,0,210,0,0,0,0,0,135,0,244,0,0,0,248,0,23,0,37,0,159,0,12,0,184,0,208,0,165,0,45,0,113,0,127,0,230,0,42,0,23,0,0,0,96,0,77,0,195,0,82,0,205,0,113,0,138,0,157,0,0,0,152,0,231,0,130,0,168,0,133,0,152,0,0,0,114,0,0,0,0,0,188,0,0,0,0,0,165,0,108,0,6,0,79,0,74,0,25,0,46,0,0,0,196,0,193,0,227,0,193,0,199,0,139,0,0,0,80,0,94,0,238,0,0,0,199,0,176,0,125,0,241,0,140,0,124,0,217,0,209,0,15,0,62,0,0,0,0,0,25,0,205,0,189,0,80,0,174,0,198,0,115,0,133,0,136,0,40,0,0,0,181,0,0,0,0,0,0,0,29,0,4,0,236,0,202,0,206,0,73,0,254,0,0,0,204,0,192,0,0,0,113,0,45,0,0,0,108,0,182,0,198,0,16,0,0,0,16,0,0,0,0,0,0,0,153,0,181,0,235,0,205,0,255,0,11,0,67,0,86,0,103,0,0,0,171,0,10,0,0,0,91,0,139,0,72,0,108,0,219,0,27,0,197,0,71,0,239,0,20,0,233,0,242,0,224,0,138,0,199,0,0,0,0,0,185,0,230,0,15,0,61,0,61,0,11,0,42,0,68,0,218,0,72,0,214,0,252,0,35,0,104,0,87,0,196,0,24,0,0,0,137,0,12,0,104,0,37,0,70,0,163,0,104,0,192,0,179,0,197,0,146,0,139,0,136,0,191,0,0,0,135,0,245,0,64,0,85,0,100,0,220,0,120,0,0,0,0,0,0,0,33,0,47,0,143,0,123,0,158,0,85,0,94,0,0,0,3,0,48,0,0,0,63,0,98,0,140,0,0,0,0,0,0,0,20,0,17,0,248,0,0,0,92,0,181,0,80,0,0,0,64,0,108,0,0,0,20,0,0,0,208,0,198,0,181,0,172,0,0,0,164,0,242,0,225,0,219,0,215,0,246,0,69,0,167,0,203,0,101,0,252,0,51,0,39,0,163,0,198,0,157,0,149,0,79,0,52,0,0,0,210,0,0,0,159,0,54,0,31,0,118,0,224,0,205,0,0,0,219,0,252,0,160,0,248,0,103,0,182,0,0,0,37,0,0,0,53,0,248,0,104,0,134,0,238,0,0,0,235,0,228,0,236,0,219,0,61,0,0,0,0,0,67,0,230,0,166,0,250,0,0,0,32,0,2,0,175,0,236,0,0,0,124,0,30,0,0,0,0,0,140,0,122,0,124,0,0,0,151,0,86,0,162,0,83,0,12,0,109,0,185,0,139,0,32,0,21,0,0,0,213,0,89,0,223,0,0,0,37,0,163,0,27,0,49,0,0,0,0,0,34,0,31,0,20,0,0,0,52,0,120,0,0,0,62,0,38,0,167,0,0,0,186,0,3,0,153,0,201,0,251,0,126,0,0,0,0,0,235,0,71,0,15,0,31,0,0,0,43,0,244,0,65,0,0,0,96,0,34,0,125,0,0,0,80,0,0,0,83,0,156,0,47,0,88,0,44,0,165,0,196,0,0,0,160,0,155,0,21,0,17,0,97,0,211,0,0,0,53,0,245,0,158,0,3,0,78,0,0,0,13,0,0,0,152,0,42,0,229,0,215,0,0,0,213,0,0,0,4,0,223,0,238,0,0,0,81,0,0,0,82,0,47,0,93,0,135,0,223,0,0,0,0,0,3,0,201,0,84,0,39,0,47,0,77,0,0,0,143,0,116,0,236,0,109,0,18,0,162,0,49,0,170,0,182,0,184,0,56,0,42,0,0,0,254,0,199,0,154,0,43,0,210,0,242,0,117,0,0,0,121,0,44,0,136,0,8,0,123,0,13,0,108,0,136,0,72,0,99,0,16,0,191,0,9,0,195,0,253,0,77,0,40,0,140,0,0,0,206,0,52,0,114,0,38,0,178,0,195,0,54,0,1,0,74,0,160,0,117,0,178,0,235,0,58,0,135,0,0,0,100,0,246,0,136,0,0,0,8,0,242,0,0,0,74,0,98,0,69,0,163,0,2,0,0,0,5,0,193,0,95,0,0,0,64,0,160,0,0,0,140,0,173,0,0,0,78,0,233,0,114,0,10,0,0,0,151,0,35,0,219,0,0,0,0,0,0,0,0,0,0,0,185,0,215,0,0,0,0,0,219,0,11,0,172,0,71,0,109,0,106,0,73,0,105,0,134,0,146,0,27,0,31,0,146,0,195,0,246,0,84,0,227,0,108,0,55,0,38,0,140,0,223,0,146,0,212,0,0,0,237,0,186,0,238,0,0,0,13,0,104,0,196,0,221,0,130,0,12,0,0,0,114,0,66,0,0,0,196,0,148,0,69,0,98,0,229,0,161,0,209,0,0,0,198,0,146,0,0,0,0,0,13,0,91,0,0,0,123,0,172,0,182,0,118,0,0,0,182,0,212,0,138,0,20,0,237,0,238,0,201,0,32,0,133,0,198,0,220,0,81,0,32,0,161,0,211,0,10,0,0,0,79,0,169,0,0,0,19,0,0,0,0,0,0,0,82,0,141,0,174,0,192,0,82,0,30,0,52,0,0,0,94,0,45,0,0,0,0,0,218,0,95,0,0,0,0,0);
signal scenario_full  : scenario_type := (83,31,79,31,79,30,15,31,109,31,60,31,60,30,60,29,218,31,116,31,242,31,203,31,203,30,212,31,7,31,157,31,157,30,237,31,130,31,89,31,118,31,212,31,130,31,50,31,188,31,136,31,136,30,146,31,146,30,178,31,73,31,73,30,87,31,255,31,183,31,123,31,66,31,194,31,181,31,124,31,122,31,201,31,201,30,201,29,109,31,46,31,89,31,2,31,134,31,59,31,59,30,127,31,4,31,213,31,5,31,231,31,59,31,9,31,48,31,198,31,215,31,208,31,253,31,139,31,139,30,252,31,5,31,233,31,228,31,124,31,172,31,62,31,7,31,113,31,44,31,25,31,9,31,229,31,135,31,177,31,92,31,54,31,189,31,205,31,178,31,178,30,239,31,20,31,137,31,169,31,162,31,249,31,55,31,209,31,134,31,134,30,211,31,126,31,216,31,101,31,37,31,150,31,182,31,211,31,211,30,232,31,232,31,102,31,232,31,232,30,75,31,75,30,106,31,243,31,47,31,47,30,157,31,12,31,97,31,71,31,119,31,55,31,125,31,145,31,60,31,60,30,157,31,125,31,215,31,50,31,210,31,56,31,56,30,204,31,95,31,105,31,13,31,223,31,223,30,35,31,184,31,184,30,72,31,222,31,222,30,222,29,71,31,52,31,52,30,117,31,83,31,83,30,144,31,250,31,60,31,60,30,139,31,131,31,79,31,97,31,97,30,248,31,219,31,182,31,59,31,223,31,140,31,140,30,49,31,65,31,65,30,80,31,106,31,107,31,20,31,138,31,185,31,109,31,240,31,4,31,33,31,157,31,220,31,220,30,59,31,86,31,86,30,44,31,191,31,227,31,56,31,56,30,89,31,150,31,177,31,177,30,240,31,221,31,206,31,130,31,60,31,241,31,22,31,241,31,241,30,178,31,84,31,74,31,27,31,27,30,72,31,132,31,132,30,157,31,243,31,243,30,11,31,204,31,228,31,199,31,33,31,33,30,143,31,143,30,10,31,225,31,189,31,119,31,119,30,239,31,148,31,188,31,130,31,110,31,245,31,245,30,19,31,31,31,31,30,37,31,117,31,129,31,23,31,154,31,154,30,46,31,72,31,72,30,153,31,201,31,224,31,13,31,13,30,218,31,4,31,140,31,140,30,5,31,5,30,239,31,10,31,74,31,74,30,5,31,128,31,76,31,76,30,135,31,130,31,130,30,255,31,25,31,7,31,65,31,157,31,157,30,90,31,157,31,121,31,182,31,249,31,249,30,152,31,185,31,107,31,124,31,164,31,183,31,210,31,210,30,210,29,135,31,244,31,244,30,248,31,23,31,37,31,159,31,12,31,184,31,208,31,165,31,45,31,113,31,127,31,230,31,42,31,23,31,23,30,96,31,77,31,195,31,82,31,205,31,113,31,138,31,157,31,157,30,152,31,231,31,130,31,168,31,133,31,152,31,152,30,114,31,114,30,114,29,188,31,188,30,188,29,165,31,108,31,6,31,79,31,74,31,25,31,46,31,46,30,196,31,193,31,227,31,193,31,199,31,139,31,139,30,80,31,94,31,238,31,238,30,199,31,176,31,125,31,241,31,140,31,124,31,217,31,209,31,15,31,62,31,62,30,62,29,25,31,205,31,189,31,80,31,174,31,198,31,115,31,133,31,136,31,40,31,40,30,181,31,181,30,181,29,181,28,29,31,4,31,236,31,202,31,206,31,73,31,254,31,254,30,204,31,192,31,192,30,113,31,45,31,45,30,108,31,182,31,198,31,16,31,16,30,16,31,16,30,16,29,16,28,153,31,181,31,235,31,205,31,255,31,11,31,67,31,86,31,103,31,103,30,171,31,10,31,10,30,91,31,139,31,72,31,108,31,219,31,27,31,197,31,71,31,239,31,20,31,233,31,242,31,224,31,138,31,199,31,199,30,199,29,185,31,230,31,15,31,61,31,61,31,11,31,42,31,68,31,218,31,72,31,214,31,252,31,35,31,104,31,87,31,196,31,24,31,24,30,137,31,12,31,104,31,37,31,70,31,163,31,104,31,192,31,179,31,197,31,146,31,139,31,136,31,191,31,191,30,135,31,245,31,64,31,85,31,100,31,220,31,120,31,120,30,120,29,120,28,33,31,47,31,143,31,123,31,158,31,85,31,94,31,94,30,3,31,48,31,48,30,63,31,98,31,140,31,140,30,140,29,140,28,20,31,17,31,248,31,248,30,92,31,181,31,80,31,80,30,64,31,108,31,108,30,20,31,20,30,208,31,198,31,181,31,172,31,172,30,164,31,242,31,225,31,219,31,215,31,246,31,69,31,167,31,203,31,101,31,252,31,51,31,39,31,163,31,198,31,157,31,149,31,79,31,52,31,52,30,210,31,210,30,159,31,54,31,31,31,118,31,224,31,205,31,205,30,219,31,252,31,160,31,248,31,103,31,182,31,182,30,37,31,37,30,53,31,248,31,104,31,134,31,238,31,238,30,235,31,228,31,236,31,219,31,61,31,61,30,61,29,67,31,230,31,166,31,250,31,250,30,32,31,2,31,175,31,236,31,236,30,124,31,30,31,30,30,30,29,140,31,122,31,124,31,124,30,151,31,86,31,162,31,83,31,12,31,109,31,185,31,139,31,32,31,21,31,21,30,213,31,89,31,223,31,223,30,37,31,163,31,27,31,49,31,49,30,49,29,34,31,31,31,20,31,20,30,52,31,120,31,120,30,62,31,38,31,167,31,167,30,186,31,3,31,153,31,201,31,251,31,126,31,126,30,126,29,235,31,71,31,15,31,31,31,31,30,43,31,244,31,65,31,65,30,96,31,34,31,125,31,125,30,80,31,80,30,83,31,156,31,47,31,88,31,44,31,165,31,196,31,196,30,160,31,155,31,21,31,17,31,97,31,211,31,211,30,53,31,245,31,158,31,3,31,78,31,78,30,13,31,13,30,152,31,42,31,229,31,215,31,215,30,213,31,213,30,4,31,223,31,238,31,238,30,81,31,81,30,82,31,47,31,93,31,135,31,223,31,223,30,223,29,3,31,201,31,84,31,39,31,47,31,77,31,77,30,143,31,116,31,236,31,109,31,18,31,162,31,49,31,170,31,182,31,184,31,56,31,42,31,42,30,254,31,199,31,154,31,43,31,210,31,242,31,117,31,117,30,121,31,44,31,136,31,8,31,123,31,13,31,108,31,136,31,72,31,99,31,16,31,191,31,9,31,195,31,253,31,77,31,40,31,140,31,140,30,206,31,52,31,114,31,38,31,178,31,195,31,54,31,1,31,74,31,160,31,117,31,178,31,235,31,58,31,135,31,135,30,100,31,246,31,136,31,136,30,8,31,242,31,242,30,74,31,98,31,69,31,163,31,2,31,2,30,5,31,193,31,95,31,95,30,64,31,160,31,160,30,140,31,173,31,173,30,78,31,233,31,114,31,10,31,10,30,151,31,35,31,219,31,219,30,219,29,219,28,219,27,219,26,185,31,215,31,215,30,215,29,219,31,11,31,172,31,71,31,109,31,106,31,73,31,105,31,134,31,146,31,27,31,31,31,146,31,195,31,246,31,84,31,227,31,108,31,55,31,38,31,140,31,223,31,146,31,212,31,212,30,237,31,186,31,238,31,238,30,13,31,104,31,196,31,221,31,130,31,12,31,12,30,114,31,66,31,66,30,196,31,148,31,69,31,98,31,229,31,161,31,209,31,209,30,198,31,146,31,146,30,146,29,13,31,91,31,91,30,123,31,172,31,182,31,118,31,118,30,182,31,212,31,138,31,20,31,237,31,238,31,201,31,32,31,133,31,198,31,220,31,81,31,32,31,161,31,211,31,10,31,10,30,79,31,169,31,169,30,19,31,19,30,19,29,19,28,82,31,141,31,174,31,192,31,82,31,30,31,52,31,52,30,94,31,45,31,45,30,45,29,218,31,95,31,95,30,95,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
