-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 605;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,149,0,243,0,48,0,246,0,103,0,19,0,0,0,142,0,228,0,49,0,146,0,223,0,10,0,124,0,105,0,189,0,92,0,151,0,91,0,8,0,0,0,176,0,181,0,1,0,72,0,3,0,1,0,196,0,224,0,59,0,223,0,206,0,132,0,195,0,149,0,58,0,254,0,0,0,0,0,0,0,207,0,240,0,104,0,163,0,88,0,63,0,28,0,73,0,115,0,144,0,153,0,0,0,63,0,12,0,255,0,40,0,51,0,74,0,18,0,152,0,0,0,0,0,0,0,46,0,104,0,129,0,0,0,102,0,129,0,177,0,226,0,236,0,48,0,94,0,0,0,3,0,0,0,63,0,218,0,85,0,155,0,44,0,48,0,165,0,164,0,202,0,176,0,167,0,148,0,251,0,23,0,24,0,91,0,222,0,68,0,162,0,239,0,229,0,0,0,120,0,221,0,209,0,79,0,245,0,0,0,47,0,62,0,78,0,201,0,29,0,0,0,226,0,132,0,125,0,139,0,115,0,212,0,0,0,246,0,68,0,0,0,0,0,227,0,50,0,89,0,70,0,95,0,208,0,122,0,67,0,172,0,225,0,95,0,95,0,189,0,0,0,2,0,131,0,232,0,0,0,104,0,0,0,128,0,122,0,56,0,0,0,113,0,0,0,68,0,135,0,145,0,96,0,15,0,104,0,0,0,97,0,212,0,69,0,0,0,232,0,80,0,0,0,37,0,13,0,0,0,0,0,49,0,81,0,200,0,0,0,248,0,40,0,116,0,0,0,226,0,243,0,98,0,220,0,161,0,71,0,241,0,220,0,73,0,20,0,13,0,174,0,10,0,220,0,82,0,3,0,0,0,254,0,0,0,127,0,150,0,37,0,215,0,52,0,0,0,3,0,118,0,99,0,182,0,0,0,0,0,0,0,0,0,174,0,125,0,205,0,161,0,167,0,210,0,242,0,31,0,0,0,0,0,123,0,78,0,0,0,74,0,230,0,160,0,40,0,178,0,0,0,174,0,157,0,249,0,37,0,97,0,48,0,0,0,0,0,228,0,236,0,197,0,25,0,81,0,132,0,241,0,239,0,0,0,28,0,255,0,92,0,76,0,181,0,41,0,166,0,108,0,183,0,94,0,33,0,254,0,239,0,228,0,150,0,104,0,190,0,215,0,48,0,136,0,0,0,124,0,163,0,180,0,82,0,173,0,224,0,211,0,0,0,0,0,227,0,0,0,128,0,111,0,242,0,86,0,154,0,191,0,99,0,204,0,22,0,152,0,83,0,175,0,192,0,73,0,0,0,93,0,82,0,23,0,174,0,154,0,38,0,211,0,57,0,126,0,27,0,187,0,163,0,207,0,0,0,89,0,131,0,0,0,193,0,0,0,96,0,103,0,253,0,0,0,0,0,181,0,43,0,0,0,171,0,135,0,33,0,11,0,134,0,152,0,0,0,12,0,154,0,7,0,181,0,71,0,135,0,252,0,39,0,0,0,26,0,190,0,156,0,22,0,22,0,0,0,215,0,0,0,134,0,169,0,69,0,0,0,0,0,0,0,0,0,190,0,230,0,175,0,61,0,215,0,50,0,248,0,138,0,159,0,190,0,9,0,96,0,0,0,180,0,196,0,0,0,6,0,83,0,198,0,134,0,203,0,176,0,76,0,0,0,231,0,65,0,141,0,0,0,100,0,127,0,233,0,62,0,0,0,78,0,100,0,122,0,0,0,66,0,0,0,128,0,131,0,59,0,30,0,124,0,227,0,73,0,234,0,52,0,0,0,112,0,0,0,0,0,0,0,146,0,46,0,0,0,112,0,132,0,231,0,0,0,120,0,18,0,186,0,8,0,139,0,213,0,1,0,211,0,210,0,23,0,0,0,89,0,6,0,223,0,23,0,80,0,101,0,214,0,0,0,106,0,55,0,158,0,0,0,0,0,231,0,21,0,41,0,117,0,26,0,118,0,222,0,233,0,0,0,172,0,105,0,242,0,222,0,223,0,0,0,40,0,85,0,64,0,0,0,184,0,0,0,249,0,164,0,92,0,177,0,7,0,95,0,2,0,0,0,111,0,122,0,135,0,22,0,214,0,138,0,0,0,0,0,226,0,113,0,93,0,0,0,0,0,0,0,0,0,2,0,0,0,0,0,114,0,101,0,30,0,0,0,187,0,87,0,0,0,170,0,0,0,183,0,180,0,247,0,249,0,0,0,83,0,27,0,41,0,60,0,59,0,53,0,167,0,140,0,206,0,218,0,178,0,126,0,11,0,0,0,209,0,218,0,170,0,21,0,39,0,136,0,181,0,36,0,46,0,50,0,158,0,139,0,84,0,247,0,0,0,79,0,124,0,0,0,136,0,89,0,246,0,109,0,163,0,0,0,11,0,0,0,136,0,32,0,0,0,11,0,108,0,103,0,0,0,0,0,0,0,56,0,96,0,0,0,250,0,56,0,167,0,0,0,178,0,16,0,5,0,97,0,193,0,86,0,199,0,0,0,0,0,0,0,0,0,174,0,103,0,109,0,71,0,107,0,89,0,167,0,0,0,130,0,10,0,0,0,216,0,239,0,123,0,97,0,0,0,16,0,113,0,54,0,222,0,0,0,151,0,72,0,139,0,235,0,0,0,28,0,0,0,208,0,17,0,0,0,167,0,222,0,173,0,55,0,15,0,75,0,137,0,190,0,236,0,55,0,0,0,75,0,16,0);
signal scenario_full  : scenario_type := (0,0,149,31,243,31,48,31,246,31,103,31,19,31,19,30,142,31,228,31,49,31,146,31,223,31,10,31,124,31,105,31,189,31,92,31,151,31,91,31,8,31,8,30,176,31,181,31,1,31,72,31,3,31,1,31,196,31,224,31,59,31,223,31,206,31,132,31,195,31,149,31,58,31,254,31,254,30,254,29,254,28,207,31,240,31,104,31,163,31,88,31,63,31,28,31,73,31,115,31,144,31,153,31,153,30,63,31,12,31,255,31,40,31,51,31,74,31,18,31,152,31,152,30,152,29,152,28,46,31,104,31,129,31,129,30,102,31,129,31,177,31,226,31,236,31,48,31,94,31,94,30,3,31,3,30,63,31,218,31,85,31,155,31,44,31,48,31,165,31,164,31,202,31,176,31,167,31,148,31,251,31,23,31,24,31,91,31,222,31,68,31,162,31,239,31,229,31,229,30,120,31,221,31,209,31,79,31,245,31,245,30,47,31,62,31,78,31,201,31,29,31,29,30,226,31,132,31,125,31,139,31,115,31,212,31,212,30,246,31,68,31,68,30,68,29,227,31,50,31,89,31,70,31,95,31,208,31,122,31,67,31,172,31,225,31,95,31,95,31,189,31,189,30,2,31,131,31,232,31,232,30,104,31,104,30,128,31,122,31,56,31,56,30,113,31,113,30,68,31,135,31,145,31,96,31,15,31,104,31,104,30,97,31,212,31,69,31,69,30,232,31,80,31,80,30,37,31,13,31,13,30,13,29,49,31,81,31,200,31,200,30,248,31,40,31,116,31,116,30,226,31,243,31,98,31,220,31,161,31,71,31,241,31,220,31,73,31,20,31,13,31,174,31,10,31,220,31,82,31,3,31,3,30,254,31,254,30,127,31,150,31,37,31,215,31,52,31,52,30,3,31,118,31,99,31,182,31,182,30,182,29,182,28,182,27,174,31,125,31,205,31,161,31,167,31,210,31,242,31,31,31,31,30,31,29,123,31,78,31,78,30,74,31,230,31,160,31,40,31,178,31,178,30,174,31,157,31,249,31,37,31,97,31,48,31,48,30,48,29,228,31,236,31,197,31,25,31,81,31,132,31,241,31,239,31,239,30,28,31,255,31,92,31,76,31,181,31,41,31,166,31,108,31,183,31,94,31,33,31,254,31,239,31,228,31,150,31,104,31,190,31,215,31,48,31,136,31,136,30,124,31,163,31,180,31,82,31,173,31,224,31,211,31,211,30,211,29,227,31,227,30,128,31,111,31,242,31,86,31,154,31,191,31,99,31,204,31,22,31,152,31,83,31,175,31,192,31,73,31,73,30,93,31,82,31,23,31,174,31,154,31,38,31,211,31,57,31,126,31,27,31,187,31,163,31,207,31,207,30,89,31,131,31,131,30,193,31,193,30,96,31,103,31,253,31,253,30,253,29,181,31,43,31,43,30,171,31,135,31,33,31,11,31,134,31,152,31,152,30,12,31,154,31,7,31,181,31,71,31,135,31,252,31,39,31,39,30,26,31,190,31,156,31,22,31,22,31,22,30,215,31,215,30,134,31,169,31,69,31,69,30,69,29,69,28,69,27,190,31,230,31,175,31,61,31,215,31,50,31,248,31,138,31,159,31,190,31,9,31,96,31,96,30,180,31,196,31,196,30,6,31,83,31,198,31,134,31,203,31,176,31,76,31,76,30,231,31,65,31,141,31,141,30,100,31,127,31,233,31,62,31,62,30,78,31,100,31,122,31,122,30,66,31,66,30,128,31,131,31,59,31,30,31,124,31,227,31,73,31,234,31,52,31,52,30,112,31,112,30,112,29,112,28,146,31,46,31,46,30,112,31,132,31,231,31,231,30,120,31,18,31,186,31,8,31,139,31,213,31,1,31,211,31,210,31,23,31,23,30,89,31,6,31,223,31,23,31,80,31,101,31,214,31,214,30,106,31,55,31,158,31,158,30,158,29,231,31,21,31,41,31,117,31,26,31,118,31,222,31,233,31,233,30,172,31,105,31,242,31,222,31,223,31,223,30,40,31,85,31,64,31,64,30,184,31,184,30,249,31,164,31,92,31,177,31,7,31,95,31,2,31,2,30,111,31,122,31,135,31,22,31,214,31,138,31,138,30,138,29,226,31,113,31,93,31,93,30,93,29,93,28,93,27,2,31,2,30,2,29,114,31,101,31,30,31,30,30,187,31,87,31,87,30,170,31,170,30,183,31,180,31,247,31,249,31,249,30,83,31,27,31,41,31,60,31,59,31,53,31,167,31,140,31,206,31,218,31,178,31,126,31,11,31,11,30,209,31,218,31,170,31,21,31,39,31,136,31,181,31,36,31,46,31,50,31,158,31,139,31,84,31,247,31,247,30,79,31,124,31,124,30,136,31,89,31,246,31,109,31,163,31,163,30,11,31,11,30,136,31,32,31,32,30,11,31,108,31,103,31,103,30,103,29,103,28,56,31,96,31,96,30,250,31,56,31,167,31,167,30,178,31,16,31,5,31,97,31,193,31,86,31,199,31,199,30,199,29,199,28,199,27,174,31,103,31,109,31,71,31,107,31,89,31,167,31,167,30,130,31,10,31,10,30,216,31,239,31,123,31,97,31,97,30,16,31,113,31,54,31,222,31,222,30,151,31,72,31,139,31,235,31,235,30,28,31,28,30,208,31,17,31,17,30,167,31,222,31,173,31,55,31,15,31,75,31,137,31,190,31,236,31,55,31,55,30,75,31,16,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
