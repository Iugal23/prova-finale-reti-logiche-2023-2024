-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_846 is
end project_tb_846;

architecture project_tb_arch_846 of project_tb_846 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 346;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (104,0,23,0,102,0,0,0,248,0,80,0,0,0,137,0,245,0,250,0,123,0,117,0,0,0,161,0,228,0,62,0,145,0,104,0,152,0,129,0,218,0,64,0,134,0,78,0,142,0,0,0,1,0,44,0,8,0,0,0,76,0,30,0,184,0,123,0,199,0,0,0,0,0,102,0,102,0,173,0,73,0,0,0,0,0,0,0,0,0,148,0,136,0,198,0,214,0,89,0,50,0,94,0,26,0,3,0,0,0,214,0,169,0,0,0,11,0,33,0,0,0,0,0,242,0,0,0,149,0,190,0,0,0,0,0,215,0,232,0,36,0,0,0,0,0,202,0,235,0,159,0,6,0,45,0,16,0,0,0,163,0,134,0,0,0,19,0,9,0,0,0,37,0,115,0,147,0,0,0,221,0,156,0,111,0,125,0,179,0,60,0,109,0,32,0,203,0,135,0,168,0,177,0,22,0,0,0,0,0,101,0,239,0,155,0,0,0,70,0,115,0,225,0,98,0,35,0,194,0,0,0,4,0,34,0,144,0,56,0,93,0,30,0,77,0,17,0,110,0,230,0,197,0,25,0,85,0,130,0,181,0,201,0,224,0,0,0,43,0,156,0,101,0,212,0,127,0,186,0,14,0,236,0,0,0,7,0,172,0,0,0,179,0,8,0,0,0,191,0,189,0,226,0,248,0,0,0,167,0,98,0,184,0,0,0,36,0,189,0,146,0,162,0,154,0,131,0,249,0,19,0,0,0,118,0,153,0,230,0,0,0,49,0,0,0,178,0,251,0,135,0,197,0,4,0,114,0,161,0,234,0,75,0,6,0,185,0,246,0,50,0,196,0,0,0,0,0,19,0,244,0,94,0,83,0,19,0,201,0,25,0,31,0,30,0,79,0,0,0,0,0,239,0,0,0,0,0,11,0,0,0,134,0,75,0,24,0,124,0,0,0,167,0,254,0,159,0,100,0,11,0,55,0,43,0,0,0,219,0,81,0,110,0,219,0,186,0,71,0,185,0,127,0,0,0,0,0,9,0,12,0,229,0,41,0,0,0,20,0,35,0,166,0,85,0,81,0,51,0,79,0,190,0,176,0,0,0,242,0,36,0,0,0,0,0,0,0,167,0,0,0,92,0,4,0,99,0,18,0,26,0,5,0,101,0,190,0,206,0,53,0,126,0,59,0,0,0,96,0,168,0,239,0,221,0,253,0,76,0,186,0,0,0,33,0,0,0,98,0,0,0,17,0,89,0,251,0,33,0,177,0,64,0,180,0,98,0,243,0,215,0,165,0,242,0,0,0,165,0,187,0,20,0,0,0,47,0,102,0,114,0,0,0,83,0,88,0,44,0,117,0,57,0,0,0,118,0,189,0,35,0,23,0,204,0,18,0,98,0,203,0,26,0,74,0,0,0,102,0,41,0,0,0,177,0,61,0,88,0,107,0,226,0,161,0,9,0,185,0,204,0,253,0,253,0,176,0,140,0,0,0,224,0,247,0,57,0,27,0,18,0,23,0,230,0,72,0,179,0,90,0,153,0,105,0,0,0,107,0,88,0);
signal scenario_full  : scenario_type := (104,31,23,31,102,31,102,30,248,31,80,31,80,30,137,31,245,31,250,31,123,31,117,31,117,30,161,31,228,31,62,31,145,31,104,31,152,31,129,31,218,31,64,31,134,31,78,31,142,31,142,30,1,31,44,31,8,31,8,30,76,31,30,31,184,31,123,31,199,31,199,30,199,29,102,31,102,31,173,31,73,31,73,30,73,29,73,28,73,27,148,31,136,31,198,31,214,31,89,31,50,31,94,31,26,31,3,31,3,30,214,31,169,31,169,30,11,31,33,31,33,30,33,29,242,31,242,30,149,31,190,31,190,30,190,29,215,31,232,31,36,31,36,30,36,29,202,31,235,31,159,31,6,31,45,31,16,31,16,30,163,31,134,31,134,30,19,31,9,31,9,30,37,31,115,31,147,31,147,30,221,31,156,31,111,31,125,31,179,31,60,31,109,31,32,31,203,31,135,31,168,31,177,31,22,31,22,30,22,29,101,31,239,31,155,31,155,30,70,31,115,31,225,31,98,31,35,31,194,31,194,30,4,31,34,31,144,31,56,31,93,31,30,31,77,31,17,31,110,31,230,31,197,31,25,31,85,31,130,31,181,31,201,31,224,31,224,30,43,31,156,31,101,31,212,31,127,31,186,31,14,31,236,31,236,30,7,31,172,31,172,30,179,31,8,31,8,30,191,31,189,31,226,31,248,31,248,30,167,31,98,31,184,31,184,30,36,31,189,31,146,31,162,31,154,31,131,31,249,31,19,31,19,30,118,31,153,31,230,31,230,30,49,31,49,30,178,31,251,31,135,31,197,31,4,31,114,31,161,31,234,31,75,31,6,31,185,31,246,31,50,31,196,31,196,30,196,29,19,31,244,31,94,31,83,31,19,31,201,31,25,31,31,31,30,31,79,31,79,30,79,29,239,31,239,30,239,29,11,31,11,30,134,31,75,31,24,31,124,31,124,30,167,31,254,31,159,31,100,31,11,31,55,31,43,31,43,30,219,31,81,31,110,31,219,31,186,31,71,31,185,31,127,31,127,30,127,29,9,31,12,31,229,31,41,31,41,30,20,31,35,31,166,31,85,31,81,31,51,31,79,31,190,31,176,31,176,30,242,31,36,31,36,30,36,29,36,28,167,31,167,30,92,31,4,31,99,31,18,31,26,31,5,31,101,31,190,31,206,31,53,31,126,31,59,31,59,30,96,31,168,31,239,31,221,31,253,31,76,31,186,31,186,30,33,31,33,30,98,31,98,30,17,31,89,31,251,31,33,31,177,31,64,31,180,31,98,31,243,31,215,31,165,31,242,31,242,30,165,31,187,31,20,31,20,30,47,31,102,31,114,31,114,30,83,31,88,31,44,31,117,31,57,31,57,30,118,31,189,31,35,31,23,31,204,31,18,31,98,31,203,31,26,31,74,31,74,30,102,31,41,31,41,30,177,31,61,31,88,31,107,31,226,31,161,31,9,31,185,31,204,31,253,31,253,31,176,31,140,31,140,30,224,31,247,31,57,31,27,31,18,31,23,31,230,31,72,31,179,31,90,31,153,31,105,31,105,30,107,31,88,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
