-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_967 is
end project_tb_967;

architecture project_tb_arch_967 of project_tb_967 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 340;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (218,0,190,0,175,0,61,0,176,0,57,0,232,0,104,0,255,0,23,0,86,0,47,0,0,0,0,0,76,0,14,0,78,0,168,0,0,0,88,0,22,0,45,0,148,0,239,0,54,0,176,0,73,0,14,0,0,0,0,0,127,0,233,0,211,0,222,0,0,0,71,0,80,0,113,0,221,0,188,0,116,0,0,0,213,0,117,0,93,0,0,0,231,0,166,0,143,0,0,0,0,0,30,0,231,0,209,0,247,0,25,0,198,0,243,0,223,0,124,0,236,0,34,0,189,0,255,0,131,0,198,0,0,0,148,0,172,0,29,0,29,0,122,0,10,0,0,0,36,0,73,0,4,0,114,0,99,0,23,0,185,0,69,0,234,0,228,0,158,0,238,0,97,0,225,0,0,0,238,0,127,0,122,0,221,0,140,0,0,0,206,0,17,0,222,0,18,0,130,0,164,0,55,0,45,0,148,0,41,0,160,0,0,0,248,0,0,0,229,0,254,0,0,0,252,0,152,0,227,0,157,0,176,0,79,0,113,0,219,0,13,0,225,0,104,0,68,0,159,0,235,0,163,0,198,0,175,0,16,0,215,0,43,0,241,0,225,0,150,0,0,0,137,0,58,0,161,0,68,0,45,0,234,0,165,0,82,0,173,0,246,0,83,0,212,0,16,0,0,0,35,0,168,0,0,0,27,0,71,0,106,0,227,0,85,0,115,0,0,0,117,0,0,0,202,0,4,0,0,0,0,0,93,0,12,0,252,0,144,0,0,0,0,0,122,0,54,0,15,0,174,0,167,0,79,0,150,0,37,0,244,0,6,0,0,0,231,0,246,0,133,0,170,0,135,0,66,0,0,0,0,0,171,0,119,0,229,0,102,0,123,0,152,0,0,0,0,0,37,0,215,0,120,0,185,0,61,0,196,0,112,0,116,0,0,0,0,0,202,0,74,0,178,0,0,0,82,0,85,0,220,0,229,0,187,0,149,0,239,0,0,0,152,0,0,0,191,0,0,0,0,0,0,0,0,0,23,0,0,0,15,0,250,0,248,0,80,0,27,0,70,0,177,0,0,0,0,0,17,0,117,0,11,0,0,0,0,0,145,0,133,0,41,0,223,0,215,0,91,0,0,0,211,0,95,0,148,0,0,0,184,0,0,0,65,0,0,0,16,0,16,0,93,0,0,0,94,0,0,0,41,0,101,0,110,0,167,0,133,0,98,0,0,0,95,0,92,0,32,0,51,0,0,0,93,0,82,0,116,0,39,0,69,0,46,0,0,0,198,0,231,0,170,0,156,0,143,0,53,0,203,0,22,0,215,0,84,0,145,0,0,0,154,0,43,0,11,0,225,0,248,0,0,0,174,0,0,0,66,0,108,0,15,0,200,0,3,0,168,0,0,0,23,0,126,0,6,0,27,0,27,0,4,0,217,0,47,0,122,0,253,0,216,0,182,0,253,0,75,0,142,0,232,0,148,0,18,0,165,0,118,0,102,0,243,0,87,0,32,0,197,0,106,0,139,0,31,0,155,0);
signal scenario_full  : scenario_type := (218,31,190,31,175,31,61,31,176,31,57,31,232,31,104,31,255,31,23,31,86,31,47,31,47,30,47,29,76,31,14,31,78,31,168,31,168,30,88,31,22,31,45,31,148,31,239,31,54,31,176,31,73,31,14,31,14,30,14,29,127,31,233,31,211,31,222,31,222,30,71,31,80,31,113,31,221,31,188,31,116,31,116,30,213,31,117,31,93,31,93,30,231,31,166,31,143,31,143,30,143,29,30,31,231,31,209,31,247,31,25,31,198,31,243,31,223,31,124,31,236,31,34,31,189,31,255,31,131,31,198,31,198,30,148,31,172,31,29,31,29,31,122,31,10,31,10,30,36,31,73,31,4,31,114,31,99,31,23,31,185,31,69,31,234,31,228,31,158,31,238,31,97,31,225,31,225,30,238,31,127,31,122,31,221,31,140,31,140,30,206,31,17,31,222,31,18,31,130,31,164,31,55,31,45,31,148,31,41,31,160,31,160,30,248,31,248,30,229,31,254,31,254,30,252,31,152,31,227,31,157,31,176,31,79,31,113,31,219,31,13,31,225,31,104,31,68,31,159,31,235,31,163,31,198,31,175,31,16,31,215,31,43,31,241,31,225,31,150,31,150,30,137,31,58,31,161,31,68,31,45,31,234,31,165,31,82,31,173,31,246,31,83,31,212,31,16,31,16,30,35,31,168,31,168,30,27,31,71,31,106,31,227,31,85,31,115,31,115,30,117,31,117,30,202,31,4,31,4,30,4,29,93,31,12,31,252,31,144,31,144,30,144,29,122,31,54,31,15,31,174,31,167,31,79,31,150,31,37,31,244,31,6,31,6,30,231,31,246,31,133,31,170,31,135,31,66,31,66,30,66,29,171,31,119,31,229,31,102,31,123,31,152,31,152,30,152,29,37,31,215,31,120,31,185,31,61,31,196,31,112,31,116,31,116,30,116,29,202,31,74,31,178,31,178,30,82,31,85,31,220,31,229,31,187,31,149,31,239,31,239,30,152,31,152,30,191,31,191,30,191,29,191,28,191,27,23,31,23,30,15,31,250,31,248,31,80,31,27,31,70,31,177,31,177,30,177,29,17,31,117,31,11,31,11,30,11,29,145,31,133,31,41,31,223,31,215,31,91,31,91,30,211,31,95,31,148,31,148,30,184,31,184,30,65,31,65,30,16,31,16,31,93,31,93,30,94,31,94,30,41,31,101,31,110,31,167,31,133,31,98,31,98,30,95,31,92,31,32,31,51,31,51,30,93,31,82,31,116,31,39,31,69,31,46,31,46,30,198,31,231,31,170,31,156,31,143,31,53,31,203,31,22,31,215,31,84,31,145,31,145,30,154,31,43,31,11,31,225,31,248,31,248,30,174,31,174,30,66,31,108,31,15,31,200,31,3,31,168,31,168,30,23,31,126,31,6,31,27,31,27,31,4,31,217,31,47,31,122,31,253,31,216,31,182,31,253,31,75,31,142,31,232,31,148,31,18,31,165,31,118,31,102,31,243,31,87,31,32,31,197,31,106,31,139,31,31,31,155,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
