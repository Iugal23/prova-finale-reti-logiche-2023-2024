-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 666;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (82,0,0,0,60,0,0,0,35,0,173,0,170,0,215,0,187,0,37,0,38,0,250,0,171,0,140,0,0,0,172,0,6,0,209,0,0,0,186,0,185,0,0,0,8,0,0,0,153,0,198,0,0,0,0,0,76,0,209,0,144,0,40,0,215,0,104,0,31,0,0,0,252,0,215,0,106,0,216,0,150,0,231,0,0,0,13,0,100,0,0,0,147,0,239,0,180,0,125,0,13,0,4,0,0,0,178,0,30,0,0,0,183,0,128,0,7,0,0,0,240,0,101,0,48,0,40,0,151,0,90,0,5,0,232,0,0,0,0,0,110,0,4,0,168,0,143,0,147,0,11,0,231,0,105,0,178,0,24,0,104,0,38,0,163,0,82,0,129,0,0,0,103,0,107,0,226,0,77,0,0,0,16,0,115,0,155,0,127,0,233,0,213,0,11,0,17,0,148,0,100,0,203,0,134,0,138,0,0,0,0,0,0,0,53,0,160,0,242,0,238,0,192,0,0,0,97,0,243,0,0,0,244,0,85,0,99,0,184,0,74,0,172,0,0,0,2,0,0,0,170,0,0,0,183,0,0,0,0,0,40,0,146,0,78,0,0,0,2,0,16,0,0,0,196,0,46,0,1,0,8,0,0,0,69,0,150,0,202,0,126,0,203,0,194,0,185,0,234,0,89,0,220,0,35,0,42,0,225,0,71,0,79,0,193,0,21,0,145,0,173,0,145,0,86,0,214,0,202,0,65,0,53,0,46,0,0,0,143,0,0,0,30,0,89,0,122,0,177,0,161,0,27,0,0,0,41,0,15,0,114,0,77,0,139,0,96,0,0,0,246,0,150,0,137,0,138,0,132,0,0,0,46,0,178,0,0,0,89,0,226,0,246,0,203,0,211,0,208,0,144,0,178,0,46,0,249,0,160,0,67,0,47,0,12,0,250,0,161,0,241,0,178,0,20,0,0,0,0,0,0,0,9,0,203,0,71,0,0,0,66,0,222,0,127,0,79,0,200,0,0,0,86,0,0,0,180,0,0,0,112,0,67,0,0,0,33,0,23,0,178,0,59,0,97,0,249,0,98,0,65,0,0,0,0,0,7,0,52,0,85,0,127,0,0,0,41,0,118,0,0,0,41,0,138,0,227,0,64,0,78,0,21,0,155,0,213,0,226,0,0,0,100,0,235,0,70,0,108,0,189,0,181,0,0,0,19,0,239,0,160,0,165,0,77,0,173,0,238,0,142,0,212,0,9,0,110,0,158,0,0,0,0,0,0,0,78,0,0,0,77,0,52,0,0,0,75,0,98,0,86,0,0,0,0,0,0,0,190,0,51,0,142,0,71,0,63,0,0,0,0,0,170,0,28,0,175,0,110,0,0,0,159,0,0,0,32,0,0,0,200,0,229,0,126,0,101,0,248,0,37,0,185,0,159,0,51,0,117,0,18,0,203,0,70,0,148,0,149,0,132,0,0,0,18,0,111,0,212,0,156,0,100,0,36,0,26,0,120,0,0,0,249,0,77,0,0,0,0,0,14,0,243,0,0,0,219,0,87,0,109,0,253,0,32,0,15,0,251,0,0,0,228,0,236,0,210,0,195,0,229,0,0,0,106,0,0,0,227,0,24,0,129,0,204,0,255,0,98,0,96,0,131,0,166,0,134,0,223,0,0,0,30,0,168,0,78,0,166,0,122,0,0,0,46,0,181,0,23,0,0,0,0,0,109,0,0,0,229,0,112,0,20,0,87,0,134,0,142,0,101,0,128,0,117,0,33,0,79,0,0,0,0,0,193,0,214,0,148,0,86,0,89,0,0,0,250,0,0,0,34,0,0,0,51,0,149,0,0,0,144,0,142,0,0,0,229,0,233,0,0,0,197,0,68,0,231,0,165,0,228,0,11,0,0,0,255,0,31,0,223,0,0,0,46,0,133,0,213,0,97,0,190,0,0,0,54,0,3,0,0,0,253,0,34,0,104,0,235,0,173,0,205,0,0,0,239,0,96,0,90,0,225,0,36,0,107,0,38,0,116,0,216,0,214,0,106,0,131,0,0,0,245,0,202,0,209,0,72,0,199,0,180,0,12,0,225,0,27,0,75,0,106,0,250,0,34,0,83,0,0,0,180,0,223,0,0,0,17,0,147,0,131,0,126,0,147,0,139,0,168,0,84,0,189,0,161,0,0,0,0,0,110,0,180,0,179,0,225,0,121,0,171,0,0,0,0,0,127,0,81,0,114,0,248,0,0,0,51,0,157,0,235,0,95,0,173,0,142,0,17,0,83,0,216,0,65,0,163,0,138,0,153,0,43,0,0,0,37,0,159,0,162,0,178,0,56,0,178,0,110,0,202,0,21,0,0,0,0,0,64,0,141,0,201,0,0,0,191,0,59,0,64,0,27,0,145,0,24,0,68,0,181,0,228,0,56,0,107,0,124,0,0,0,46,0,246,0,58,0,220,0,0,0,57,0,52,0,90,0,0,0,87,0,170,0,0,0,0,0,228,0,4,0,4,0,3,0,0,0,18,0,103,0,183,0,27,0,29,0,102,0,241,0,0,0,160,0,167,0,48,0,65,0,0,0,0,0,0,0,22,0,50,0,169,0,0,0,228,0,186,0,2,0,87,0,44,0,115,0,65,0,224,0,30,0,124,0,219,0,0,0,9,0,0,0,14,0,66,0,0,0,225,0,104,0,255,0,0,0,95,0,16,0,215,0,193,0,165,0,47,0,72,0,28,0,0,0,163,0,236,0,0,0,184,0,34,0,133,0,81,0,0,0,191,0,0,0,91,0,228,0,247,0,131,0,97,0,240,0,84,0,188,0,170,0,0,0,233,0,166,0,0,0,83,0,134,0,56,0,7,0,113,0,0,0,208,0,205,0,217,0,0,0,221,0,44,0,112,0,128,0,65,0,183,0,44,0,0,0,238,0,47,0,83,0,87,0,157,0,34,0,58,0,174,0,0,0,197,0,8,0,168,0,53,0,206,0,43,0,231,0);
signal scenario_full  : scenario_type := (82,31,82,30,60,31,60,30,35,31,173,31,170,31,215,31,187,31,37,31,38,31,250,31,171,31,140,31,140,30,172,31,6,31,209,31,209,30,186,31,185,31,185,30,8,31,8,30,153,31,198,31,198,30,198,29,76,31,209,31,144,31,40,31,215,31,104,31,31,31,31,30,252,31,215,31,106,31,216,31,150,31,231,31,231,30,13,31,100,31,100,30,147,31,239,31,180,31,125,31,13,31,4,31,4,30,178,31,30,31,30,30,183,31,128,31,7,31,7,30,240,31,101,31,48,31,40,31,151,31,90,31,5,31,232,31,232,30,232,29,110,31,4,31,168,31,143,31,147,31,11,31,231,31,105,31,178,31,24,31,104,31,38,31,163,31,82,31,129,31,129,30,103,31,107,31,226,31,77,31,77,30,16,31,115,31,155,31,127,31,233,31,213,31,11,31,17,31,148,31,100,31,203,31,134,31,138,31,138,30,138,29,138,28,53,31,160,31,242,31,238,31,192,31,192,30,97,31,243,31,243,30,244,31,85,31,99,31,184,31,74,31,172,31,172,30,2,31,2,30,170,31,170,30,183,31,183,30,183,29,40,31,146,31,78,31,78,30,2,31,16,31,16,30,196,31,46,31,1,31,8,31,8,30,69,31,150,31,202,31,126,31,203,31,194,31,185,31,234,31,89,31,220,31,35,31,42,31,225,31,71,31,79,31,193,31,21,31,145,31,173,31,145,31,86,31,214,31,202,31,65,31,53,31,46,31,46,30,143,31,143,30,30,31,89,31,122,31,177,31,161,31,27,31,27,30,41,31,15,31,114,31,77,31,139,31,96,31,96,30,246,31,150,31,137,31,138,31,132,31,132,30,46,31,178,31,178,30,89,31,226,31,246,31,203,31,211,31,208,31,144,31,178,31,46,31,249,31,160,31,67,31,47,31,12,31,250,31,161,31,241,31,178,31,20,31,20,30,20,29,20,28,9,31,203,31,71,31,71,30,66,31,222,31,127,31,79,31,200,31,200,30,86,31,86,30,180,31,180,30,112,31,67,31,67,30,33,31,23,31,178,31,59,31,97,31,249,31,98,31,65,31,65,30,65,29,7,31,52,31,85,31,127,31,127,30,41,31,118,31,118,30,41,31,138,31,227,31,64,31,78,31,21,31,155,31,213,31,226,31,226,30,100,31,235,31,70,31,108,31,189,31,181,31,181,30,19,31,239,31,160,31,165,31,77,31,173,31,238,31,142,31,212,31,9,31,110,31,158,31,158,30,158,29,158,28,78,31,78,30,77,31,52,31,52,30,75,31,98,31,86,31,86,30,86,29,86,28,190,31,51,31,142,31,71,31,63,31,63,30,63,29,170,31,28,31,175,31,110,31,110,30,159,31,159,30,32,31,32,30,200,31,229,31,126,31,101,31,248,31,37,31,185,31,159,31,51,31,117,31,18,31,203,31,70,31,148,31,149,31,132,31,132,30,18,31,111,31,212,31,156,31,100,31,36,31,26,31,120,31,120,30,249,31,77,31,77,30,77,29,14,31,243,31,243,30,219,31,87,31,109,31,253,31,32,31,15,31,251,31,251,30,228,31,236,31,210,31,195,31,229,31,229,30,106,31,106,30,227,31,24,31,129,31,204,31,255,31,98,31,96,31,131,31,166,31,134,31,223,31,223,30,30,31,168,31,78,31,166,31,122,31,122,30,46,31,181,31,23,31,23,30,23,29,109,31,109,30,229,31,112,31,20,31,87,31,134,31,142,31,101,31,128,31,117,31,33,31,79,31,79,30,79,29,193,31,214,31,148,31,86,31,89,31,89,30,250,31,250,30,34,31,34,30,51,31,149,31,149,30,144,31,142,31,142,30,229,31,233,31,233,30,197,31,68,31,231,31,165,31,228,31,11,31,11,30,255,31,31,31,223,31,223,30,46,31,133,31,213,31,97,31,190,31,190,30,54,31,3,31,3,30,253,31,34,31,104,31,235,31,173,31,205,31,205,30,239,31,96,31,90,31,225,31,36,31,107,31,38,31,116,31,216,31,214,31,106,31,131,31,131,30,245,31,202,31,209,31,72,31,199,31,180,31,12,31,225,31,27,31,75,31,106,31,250,31,34,31,83,31,83,30,180,31,223,31,223,30,17,31,147,31,131,31,126,31,147,31,139,31,168,31,84,31,189,31,161,31,161,30,161,29,110,31,180,31,179,31,225,31,121,31,171,31,171,30,171,29,127,31,81,31,114,31,248,31,248,30,51,31,157,31,235,31,95,31,173,31,142,31,17,31,83,31,216,31,65,31,163,31,138,31,153,31,43,31,43,30,37,31,159,31,162,31,178,31,56,31,178,31,110,31,202,31,21,31,21,30,21,29,64,31,141,31,201,31,201,30,191,31,59,31,64,31,27,31,145,31,24,31,68,31,181,31,228,31,56,31,107,31,124,31,124,30,46,31,246,31,58,31,220,31,220,30,57,31,52,31,90,31,90,30,87,31,170,31,170,30,170,29,228,31,4,31,4,31,3,31,3,30,18,31,103,31,183,31,27,31,29,31,102,31,241,31,241,30,160,31,167,31,48,31,65,31,65,30,65,29,65,28,22,31,50,31,169,31,169,30,228,31,186,31,2,31,87,31,44,31,115,31,65,31,224,31,30,31,124,31,219,31,219,30,9,31,9,30,14,31,66,31,66,30,225,31,104,31,255,31,255,30,95,31,16,31,215,31,193,31,165,31,47,31,72,31,28,31,28,30,163,31,236,31,236,30,184,31,34,31,133,31,81,31,81,30,191,31,191,30,91,31,228,31,247,31,131,31,97,31,240,31,84,31,188,31,170,31,170,30,233,31,166,31,166,30,83,31,134,31,56,31,7,31,113,31,113,30,208,31,205,31,217,31,217,30,221,31,44,31,112,31,128,31,65,31,183,31,44,31,44,30,238,31,47,31,83,31,87,31,157,31,34,31,58,31,174,31,174,30,197,31,8,31,168,31,53,31,206,31,43,31,231,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
