-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 966;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (69,0,204,0,0,0,242,0,0,0,59,0,0,0,171,0,67,0,20,0,102,0,246,0,0,0,39,0,215,0,15,0,173,0,0,0,90,0,83,0,217,0,18,0,0,0,207,0,226,0,161,0,47,0,204,0,189,0,204,0,36,0,42,0,45,0,177,0,143,0,219,0,129,0,247,0,0,0,145,0,0,0,208,0,177,0,0,0,134,0,152,0,0,0,0,0,138,0,244,0,100,0,0,0,171,0,232,0,168,0,109,0,33,0,85,0,133,0,31,0,152,0,60,0,189,0,63,0,190,0,8,0,0,0,0,0,81,0,0,0,120,0,231,0,103,0,172,0,255,0,209,0,0,0,4,0,61,0,80,0,200,0,58,0,0,0,127,0,80,0,0,0,0,0,238,0,111,0,233,0,48,0,200,0,253,0,169,0,160,0,54,0,188,0,0,0,232,0,222,0,134,0,104,0,215,0,143,0,0,0,75,0,56,0,229,0,86,0,0,0,246,0,102,0,25,0,3,0,117,0,83,0,82,0,0,0,194,0,250,0,156,0,25,0,179,0,68,0,140,0,96,0,0,0,238,0,151,0,36,0,113,0,114,0,0,0,223,0,83,0,117,0,225,0,72,0,0,0,77,0,0,0,165,0,0,0,0,0,149,0,157,0,82,0,208,0,0,0,195,0,247,0,28,0,1,0,135,0,233,0,34,0,79,0,15,0,0,0,118,0,0,0,157,0,184,0,170,0,223,0,230,0,120,0,2,0,96,0,0,0,0,0,0,0,0,0,196,0,32,0,71,0,0,0,29,0,227,0,183,0,169,0,26,0,51,0,137,0,40,0,5,0,52,0,0,0,127,0,153,0,186,0,244,0,187,0,107,0,0,0,0,0,115,0,200,0,10,0,37,0,128,0,49,0,0,0,200,0,210,0,0,0,247,0,237,0,247,0,154,0,111,0,0,0,108,0,8,0,192,0,33,0,112,0,85,0,81,0,170,0,157,0,187,0,182,0,186,0,70,0,230,0,207,0,240,0,52,0,105,0,167,0,0,0,58,0,64,0,205,0,87,0,128,0,48,0,217,0,44,0,177,0,52,0,139,0,70,0,219,0,209,0,82,0,65,0,220,0,0,0,0,0,243,0,32,0,0,0,167,0,60,0,184,0,192,0,183,0,250,0,242,0,143,0,109,0,77,0,4,0,54,0,31,0,25,0,69,0,186,0,79,0,192,0,181,0,0,0,233,0,128,0,225,0,93,0,65,0,0,0,159,0,185,0,217,0,0,0,248,0,237,0,19,0,101,0,0,0,0,0,0,0,0,0,160,0,209,0,241,0,86,0,197,0,242,0,0,0,78,0,248,0,57,0,0,0,10,0,125,0,104,0,20,0,112,0,11,0,190,0,0,0,199,0,192,0,36,0,85,0,177,0,253,0,0,0,47,0,214,0,125,0,0,0,95,0,113,0,82,0,166,0,70,0,160,0,204,0,4,0,66,0,0,0,253,0,116,0,56,0,168,0,101,0,84,0,204,0,79,0,200,0,0,0,92,0,166,0,251,0,195,0,197,0,97,0,138,0,25,0,217,0,0,0,54,0,253,0,0,0,0,0,183,0,50,0,178,0,251,0,82,0,167,0,39,0,0,0,30,0,0,0,99,0,0,0,141,0,147,0,0,0,240,0,42,0,114,0,175,0,175,0,208,0,211,0,0,0,0,0,24,0,207,0,32,0,123,0,61,0,177,0,165,0,6,0,0,0,53,0,169,0,50,0,128,0,75,0,202,0,0,0,4,0,0,0,15,0,87,0,87,0,34,0,201,0,220,0,212,0,125,0,39,0,207,0,211,0,205,0,16,0,46,0,78,0,1,0,25,0,232,0,0,0,25,0,242,0,0,0,110,0,107,0,99,0,12,0,0,0,248,0,140,0,90,0,26,0,21,0,145,0,86,0,114,0,254,0,206,0,163,0,248,0,202,0,193,0,175,0,0,0,255,0,243,0,0,0,10,0,11,0,83,0,51,0,203,0,0,0,126,0,108,0,183,0,0,0,232,0,213,0,17,0,227,0,108,0,0,0,0,0,0,0,202,0,67,0,212,0,0,0,81,0,4,0,239,0,204,0,183,0,20,0,251,0,109,0,0,0,83,0,0,0,0,0,54,0,48,0,37,0,141,0,188,0,0,0,151,0,0,0,65,0,176,0,0,0,104,0,227,0,185,0,182,0,47,0,0,0,102,0,0,0,143,0,0,0,0,0,146,0,107,0,158,0,121,0,207,0,15,0,229,0,7,0,0,0,167,0,214,0,9,0,139,0,152,0,0,0,0,0,107,0,207,0,224,0,103,0,150,0,65,0,148,0,53,0,45,0,182,0,186,0,192,0,183,0,0,0,105,0,0,0,0,0,0,0,125,0,0,0,0,0,197,0,0,0,149,0,0,0,21,0,100,0,1,0,21,0,143,0,184,0,123,0,209,0,33,0,199,0,21,0,47,0,127,0,190,0,116,0,166,0,232,0,132,0,101,0,0,0,89,0,0,0,152,0,18,0,116,0,0,0,206,0,239,0,114,0,0,0,149,0,0,0,53,0,0,0,184,0,162,0,241,0,14,0,77,0,243,0,168,0,58,0,176,0,0,0,234,0,197,0,80,0,252,0,0,0,84,0,30,0,0,0,85,0,115,0,41,0,193,0,6,0,185,0,150,0,28,0,0,0,214,0,55,0,69,0,13,0,180,0,120,0,192,0,0,0,0,0,0,0,165,0,193,0,136,0,174,0,0,0,0,0,170,0,173,0,254,0,208,0,206,0,11,0,80,0,0,0,174,0,60,0,136,0,63,0,0,0,74,0,49,0,132,0,22,0,0,0,123,0,0,0,82,0,0,0,254,0,24,0,0,0,218,0,180,0,0,0,74,0,151,0,6,0,176,0,49,0,160,0,30,0,0,0,173,0,0,0,0,0,0,0,120,0,118,0,233,0,69,0,150,0,101,0,0,0,218,0,0,0,0,0,184,0,159,0,76,0,71,0,246,0,82,0,84,0,174,0,124,0,203,0,61,0,231,0,245,0,112,0,123,0,0,0,82,0,0,0,0,0,205,0,242,0,108,0,92,0,99,0,53,0,184,0,47,0,19,0,249,0,197,0,155,0,165,0,240,0,129,0,121,0,56,0,79,0,4,0,143,0,38,0,0,0,143,0,92,0,208,0,98,0,237,0,46,0,97,0,0,0,172,0,178,0,0,0,137,0,231,0,0,0,94,0,0,0,246,0,159,0,30,0,0,0,0,0,230,0,42,0,216,0,60,0,207,0,47,0,0,0,69,0,224,0,44,0,137,0,46,0,188,0,0,0,126,0,79,0,144,0,0,0,0,0,126,0,209,0,76,0,250,0,0,0,166,0,26,0,251,0,0,0,236,0,0,0,132,0,167,0,2,0,114,0,101,0,155,0,218,0,126,0,238,0,104,0,0,0,38,0,44,0,79,0,209,0,81,0,18,0,248,0,87,0,168,0,0,0,19,0,0,0,94,0,211,0,0,0,239,0,69,0,0,0,44,0,114,0,230,0,247,0,0,0,0,0,162,0,53,0,0,0,96,0,93,0,59,0,105,0,198,0,30,0,69,0,0,0,237,0,0,0,100,0,201,0,82,0,0,0,46,0,166,0,215,0,0,0,53,0,80,0,194,0,8,0,79,0,6,0,125,0,85,0,8,0,98,0,0,0,225,0,110,0,251,0,51,0,0,0,131,0,112,0,128,0,153,0,10,0,182,0,80,0,207,0,173,0,122,0,171,0,0,0,235,0,49,0,0,0,76,0,185,0,189,0,0,0,0,0,0,0,158,0,0,0,225,0,206,0,48,0,205,0,171,0,250,0,184,0,8,0,177,0,78,0,181,0,0,0,36,0,43,0,101,0,188,0,233,0,163,0,124,0,236,0,13,0,196,0,0,0,0,0,95,0,91,0,207,0,48,0,135,0,34,0,0,0,0,0,0,0,107,0,9,0,225,0,34,0,171,0,29,0,0,0,133,0,74,0,0,0,160,0,28,0,225,0,186,0,0,0,46,0,241,0,224,0,92,0,22,0,113,0,0,0,21,0,176,0,140,0,77,0,161,0,81,0,45,0,48,0,5,0,64,0,140,0,181,0,0,0,234,0,1,0,41,0,0,0,219,0,95,0,30,0,10,0,149,0,202,0,141,0,0,0,203,0,45,0,44,0,250,0,251,0,101,0,70,0,78,0,0,0,253,0,233,0,228,0,97,0,112,0,174,0,145,0,0,0,141,0,224,0,231,0,0,0,140,0,115,0,167,0,190,0,96,0,254,0,0,0,244,0,135,0,131,0);
signal scenario_full  : scenario_type := (69,31,204,31,204,30,242,31,242,30,59,31,59,30,171,31,67,31,20,31,102,31,246,31,246,30,39,31,215,31,15,31,173,31,173,30,90,31,83,31,217,31,18,31,18,30,207,31,226,31,161,31,47,31,204,31,189,31,204,31,36,31,42,31,45,31,177,31,143,31,219,31,129,31,247,31,247,30,145,31,145,30,208,31,177,31,177,30,134,31,152,31,152,30,152,29,138,31,244,31,100,31,100,30,171,31,232,31,168,31,109,31,33,31,85,31,133,31,31,31,152,31,60,31,189,31,63,31,190,31,8,31,8,30,8,29,81,31,81,30,120,31,231,31,103,31,172,31,255,31,209,31,209,30,4,31,61,31,80,31,200,31,58,31,58,30,127,31,80,31,80,30,80,29,238,31,111,31,233,31,48,31,200,31,253,31,169,31,160,31,54,31,188,31,188,30,232,31,222,31,134,31,104,31,215,31,143,31,143,30,75,31,56,31,229,31,86,31,86,30,246,31,102,31,25,31,3,31,117,31,83,31,82,31,82,30,194,31,250,31,156,31,25,31,179,31,68,31,140,31,96,31,96,30,238,31,151,31,36,31,113,31,114,31,114,30,223,31,83,31,117,31,225,31,72,31,72,30,77,31,77,30,165,31,165,30,165,29,149,31,157,31,82,31,208,31,208,30,195,31,247,31,28,31,1,31,135,31,233,31,34,31,79,31,15,31,15,30,118,31,118,30,157,31,184,31,170,31,223,31,230,31,120,31,2,31,96,31,96,30,96,29,96,28,96,27,196,31,32,31,71,31,71,30,29,31,227,31,183,31,169,31,26,31,51,31,137,31,40,31,5,31,52,31,52,30,127,31,153,31,186,31,244,31,187,31,107,31,107,30,107,29,115,31,200,31,10,31,37,31,128,31,49,31,49,30,200,31,210,31,210,30,247,31,237,31,247,31,154,31,111,31,111,30,108,31,8,31,192,31,33,31,112,31,85,31,81,31,170,31,157,31,187,31,182,31,186,31,70,31,230,31,207,31,240,31,52,31,105,31,167,31,167,30,58,31,64,31,205,31,87,31,128,31,48,31,217,31,44,31,177,31,52,31,139,31,70,31,219,31,209,31,82,31,65,31,220,31,220,30,220,29,243,31,32,31,32,30,167,31,60,31,184,31,192,31,183,31,250,31,242,31,143,31,109,31,77,31,4,31,54,31,31,31,25,31,69,31,186,31,79,31,192,31,181,31,181,30,233,31,128,31,225,31,93,31,65,31,65,30,159,31,185,31,217,31,217,30,248,31,237,31,19,31,101,31,101,30,101,29,101,28,101,27,160,31,209,31,241,31,86,31,197,31,242,31,242,30,78,31,248,31,57,31,57,30,10,31,125,31,104,31,20,31,112,31,11,31,190,31,190,30,199,31,192,31,36,31,85,31,177,31,253,31,253,30,47,31,214,31,125,31,125,30,95,31,113,31,82,31,166,31,70,31,160,31,204,31,4,31,66,31,66,30,253,31,116,31,56,31,168,31,101,31,84,31,204,31,79,31,200,31,200,30,92,31,166,31,251,31,195,31,197,31,97,31,138,31,25,31,217,31,217,30,54,31,253,31,253,30,253,29,183,31,50,31,178,31,251,31,82,31,167,31,39,31,39,30,30,31,30,30,99,31,99,30,141,31,147,31,147,30,240,31,42,31,114,31,175,31,175,31,208,31,211,31,211,30,211,29,24,31,207,31,32,31,123,31,61,31,177,31,165,31,6,31,6,30,53,31,169,31,50,31,128,31,75,31,202,31,202,30,4,31,4,30,15,31,87,31,87,31,34,31,201,31,220,31,212,31,125,31,39,31,207,31,211,31,205,31,16,31,46,31,78,31,1,31,25,31,232,31,232,30,25,31,242,31,242,30,110,31,107,31,99,31,12,31,12,30,248,31,140,31,90,31,26,31,21,31,145,31,86,31,114,31,254,31,206,31,163,31,248,31,202,31,193,31,175,31,175,30,255,31,243,31,243,30,10,31,11,31,83,31,51,31,203,31,203,30,126,31,108,31,183,31,183,30,232,31,213,31,17,31,227,31,108,31,108,30,108,29,108,28,202,31,67,31,212,31,212,30,81,31,4,31,239,31,204,31,183,31,20,31,251,31,109,31,109,30,83,31,83,30,83,29,54,31,48,31,37,31,141,31,188,31,188,30,151,31,151,30,65,31,176,31,176,30,104,31,227,31,185,31,182,31,47,31,47,30,102,31,102,30,143,31,143,30,143,29,146,31,107,31,158,31,121,31,207,31,15,31,229,31,7,31,7,30,167,31,214,31,9,31,139,31,152,31,152,30,152,29,107,31,207,31,224,31,103,31,150,31,65,31,148,31,53,31,45,31,182,31,186,31,192,31,183,31,183,30,105,31,105,30,105,29,105,28,125,31,125,30,125,29,197,31,197,30,149,31,149,30,21,31,100,31,1,31,21,31,143,31,184,31,123,31,209,31,33,31,199,31,21,31,47,31,127,31,190,31,116,31,166,31,232,31,132,31,101,31,101,30,89,31,89,30,152,31,18,31,116,31,116,30,206,31,239,31,114,31,114,30,149,31,149,30,53,31,53,30,184,31,162,31,241,31,14,31,77,31,243,31,168,31,58,31,176,31,176,30,234,31,197,31,80,31,252,31,252,30,84,31,30,31,30,30,85,31,115,31,41,31,193,31,6,31,185,31,150,31,28,31,28,30,214,31,55,31,69,31,13,31,180,31,120,31,192,31,192,30,192,29,192,28,165,31,193,31,136,31,174,31,174,30,174,29,170,31,173,31,254,31,208,31,206,31,11,31,80,31,80,30,174,31,60,31,136,31,63,31,63,30,74,31,49,31,132,31,22,31,22,30,123,31,123,30,82,31,82,30,254,31,24,31,24,30,218,31,180,31,180,30,74,31,151,31,6,31,176,31,49,31,160,31,30,31,30,30,173,31,173,30,173,29,173,28,120,31,118,31,233,31,69,31,150,31,101,31,101,30,218,31,218,30,218,29,184,31,159,31,76,31,71,31,246,31,82,31,84,31,174,31,124,31,203,31,61,31,231,31,245,31,112,31,123,31,123,30,82,31,82,30,82,29,205,31,242,31,108,31,92,31,99,31,53,31,184,31,47,31,19,31,249,31,197,31,155,31,165,31,240,31,129,31,121,31,56,31,79,31,4,31,143,31,38,31,38,30,143,31,92,31,208,31,98,31,237,31,46,31,97,31,97,30,172,31,178,31,178,30,137,31,231,31,231,30,94,31,94,30,246,31,159,31,30,31,30,30,30,29,230,31,42,31,216,31,60,31,207,31,47,31,47,30,69,31,224,31,44,31,137,31,46,31,188,31,188,30,126,31,79,31,144,31,144,30,144,29,126,31,209,31,76,31,250,31,250,30,166,31,26,31,251,31,251,30,236,31,236,30,132,31,167,31,2,31,114,31,101,31,155,31,218,31,126,31,238,31,104,31,104,30,38,31,44,31,79,31,209,31,81,31,18,31,248,31,87,31,168,31,168,30,19,31,19,30,94,31,211,31,211,30,239,31,69,31,69,30,44,31,114,31,230,31,247,31,247,30,247,29,162,31,53,31,53,30,96,31,93,31,59,31,105,31,198,31,30,31,69,31,69,30,237,31,237,30,100,31,201,31,82,31,82,30,46,31,166,31,215,31,215,30,53,31,80,31,194,31,8,31,79,31,6,31,125,31,85,31,8,31,98,31,98,30,225,31,110,31,251,31,51,31,51,30,131,31,112,31,128,31,153,31,10,31,182,31,80,31,207,31,173,31,122,31,171,31,171,30,235,31,49,31,49,30,76,31,185,31,189,31,189,30,189,29,189,28,158,31,158,30,225,31,206,31,48,31,205,31,171,31,250,31,184,31,8,31,177,31,78,31,181,31,181,30,36,31,43,31,101,31,188,31,233,31,163,31,124,31,236,31,13,31,196,31,196,30,196,29,95,31,91,31,207,31,48,31,135,31,34,31,34,30,34,29,34,28,107,31,9,31,225,31,34,31,171,31,29,31,29,30,133,31,74,31,74,30,160,31,28,31,225,31,186,31,186,30,46,31,241,31,224,31,92,31,22,31,113,31,113,30,21,31,176,31,140,31,77,31,161,31,81,31,45,31,48,31,5,31,64,31,140,31,181,31,181,30,234,31,1,31,41,31,41,30,219,31,95,31,30,31,10,31,149,31,202,31,141,31,141,30,203,31,45,31,44,31,250,31,251,31,101,31,70,31,78,31,78,30,253,31,233,31,228,31,97,31,112,31,174,31,145,31,145,30,141,31,224,31,231,31,231,30,140,31,115,31,167,31,190,31,96,31,254,31,254,30,244,31,135,31,131,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
