-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 979;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (223,0,17,0,85,0,209,0,106,0,42,0,172,0,254,0,181,0,0,0,185,0,71,0,113,0,48,0,0,0,111,0,0,0,0,0,140,0,241,0,4,0,155,0,79,0,233,0,45,0,0,0,0,0,0,0,163,0,0,0,121,0,17,0,0,0,50,0,131,0,66,0,215,0,0,0,85,0,186,0,182,0,56,0,210,0,229,0,63,0,178,0,237,0,31,0,11,0,244,0,149,0,0,0,172,0,200,0,150,0,187,0,0,0,143,0,121,0,0,0,141,0,208,0,38,0,135,0,205,0,167,0,0,0,137,0,21,0,118,0,108,0,52,0,184,0,0,0,0,0,214,0,238,0,13,0,82,0,0,0,189,0,58,0,0,0,39,0,79,0,163,0,162,0,117,0,0,0,250,0,221,0,4,0,69,0,161,0,41,0,169,0,241,0,35,0,45,0,158,0,45,0,14,0,168,0,85,0,0,0,89,0,5,0,103,0,124,0,0,0,195,0,151,0,17,0,234,0,0,0,182,0,211,0,183,0,124,0,197,0,0,0,165,0,241,0,98,0,96,0,0,0,132,0,221,0,178,0,192,0,166,0,88,0,0,0,161,0,238,0,0,0,17,0,10,0,97,0,44,0,90,0,177,0,43,0,9,0,173,0,29,0,167,0,0,0,65,0,0,0,219,0,42,0,43,0,174,0,54,0,46,0,21,0,12,0,0,0,85,0,12,0,0,0,93,0,221,0,160,0,1,0,172,0,46,0,0,0,77,0,28,0,0,0,60,0,0,0,178,0,251,0,0,0,0,0,146,0,116,0,0,0,189,0,180,0,0,0,17,0,237,0,177,0,162,0,0,0,170,0,131,0,0,0,161,0,92,0,82,0,9,0,162,0,174,0,117,0,44,0,30,0,156,0,107,0,243,0,41,0,95,0,33,0,0,0,0,0,225,0,137,0,130,0,0,0,0,0,120,0,87,0,85,0,15,0,120,0,215,0,237,0,103,0,0,0,85,0,152,0,141,0,0,0,0,0,137,0,245,0,230,0,191,0,163,0,18,0,220,0,128,0,98,0,0,0,243,0,74,0,24,0,0,0,158,0,252,0,99,0,15,0,0,0,232,0,161,0,41,0,247,0,225,0,94,0,0,0,124,0,56,0,242,0,215,0,0,0,230,0,8,0,221,0,194,0,89,0,253,0,164,0,77,0,0,0,106,0,74,0,176,0,69,0,138,0,109,0,228,0,179,0,156,0,0,0,101,0,0,0,177,0,0,0,81,0,226,0,0,0,171,0,157,0,126,0,0,0,0,0,163,0,210,0,51,0,0,0,0,0,42,0,37,0,152,0,159,0,215,0,7,0,63,0,0,0,210,0,122,0,97,0,0,0,228,0,220,0,208,0,0,0,0,0,125,0,176,0,0,0,153,0,17,0,86,0,184,0,0,0,202,0,0,0,104,0,8,0,42,0,44,0,0,0,155,0,152,0,26,0,112,0,183,0,120,0,80,0,124,0,189,0,158,0,208,0,19,0,46,0,111,0,79,0,201,0,0,0,140,0,245,0,59,0,124,0,43,0,10,0,180,0,122,0,0,0,136,0,67,0,187,0,7,0,0,0,45,0,81,0,207,0,0,0,55,0,0,0,0,0,219,0,0,0,233,0,91,0,237,0,0,0,184,0,66,0,0,0,79,0,196,0,34,0,0,0,141,0,100,0,140,0,39,0,109,0,0,0,251,0,58,0,0,0,217,0,212,0,0,0,0,0,177,0,213,0,49,0,185,0,0,0,67,0,119,0,0,0,96,0,9,0,15,0,49,0,0,0,0,0,127,0,149,0,0,0,184,0,0,0,0,0,72,0,0,0,145,0,239,0,27,0,186,0,30,0,209,0,185,0,149,0,0,0,0,0,226,0,119,0,219,0,0,0,213,0,233,0,163,0,77,0,187,0,132,0,82,0,0,0,160,0,0,0,101,0,4,0,36,0,134,0,166,0,75,0,196,0,0,0,202,0,57,0,32,0,7,0,184,0,7,0,56,0,0,0,0,0,186,0,2,0,3,0,0,0,0,0,86,0,70,0,179,0,128,0,37,0,21,0,148,0,0,0,0,0,191,0,159,0,36,0,0,0,237,0,252,0,188,0,61,0,0,0,7,0,200,0,167,0,0,0,154,0,61,0,6,0,0,0,158,0,110,0,0,0,243,0,228,0,243,0,183,0,83,0,8,0,193,0,0,0,74,0,126,0,216,0,242,0,0,0,116,0,0,0,0,0,79,0,171,0,206,0,7,0,8,0,140,0,71,0,15,0,29,0,148,0,77,0,116,0,0,0,50,0,0,0,199,0,107,0,0,0,213,0,106,0,48,0,150,0,102,0,182,0,31,0,174,0,32,0,180,0,27,0,8,0,64,0,0,0,221,0,0,0,31,0,45,0,0,0,0,0,58,0,191,0,75,0,39,0,36,0,133,0,138,0,31,0,0,0,199,0,11,0,252,0,58,0,182,0,176,0,47,0,89,0,170,0,91,0,223,0,0,0,78,0,80,0,19,0,159,0,96,0,228,0,55,0,36,0,154,0,0,0,20,0,0,0,0,0,47,0,118,0,11,0,222,0,0,0,189,0,150,0,5,0,233,0,73,0,213,0,35,0,36,0,2,0,8,0,205,0,0,0,100,0,86,0,178,0,0,0,17,0,47,0,159,0,111,0,196,0,117,0,0,0,185,0,0,0,223,0,146,0,21,0,0,0,10,0,0,0,251,0,5,0,35,0,36,0,118,0,0,0,142,0,0,0,216,0,0,0,129,0,103,0,40,0,75,0,199,0,20,0,241,0,125,0,107,0,31,0,48,0,183,0,189,0,130,0,196,0,243,0,53,0,144,0,171,0,159,0,208,0,249,0,135,0,249,0,151,0,77,0,0,0,242,0,0,0,0,0,253,0,114,0,110,0,237,0,0,0,0,0,0,0,105,0,215,0,252,0,24,0,0,0,92,0,54,0,136,0,154,0,22,0,255,0,175,0,220,0,145,0,103,0,251,0,186,0,233,0,244,0,111,0,23,0,217,0,161,0,212,0,92,0,156,0,103,0,0,0,0,0,124,0,90,0,0,0,14,0,57,0,0,0,214,0,2,0,159,0,45,0,197,0,143,0,135,0,0,0,136,0,255,0,0,0,41,0,0,0,194,0,170,0,166,0,175,0,76,0,179,0,99,0,33,0,227,0,0,0,65,0,45,0,120,0,88,0,150,0,214,0,243,0,13,0,0,0,231,0,183,0,0,0,0,0,234,0,16,0,7,0,13,0,0,0,245,0,242,0,53,0,172,0,50,0,18,0,235,0,192,0,212,0,156,0,27,0,98,0,0,0,16,0,129,0,127,0,49,0,115,0,18,0,0,0,4,0,253,0,49,0,162,0,0,0,168,0,149,0,0,0,23,0,205,0,236,0,79,0,93,0,29,0,74,0,66,0,189,0,162,0,144,0,87,0,15,0,91,0,22,0,90,0,175,0,201,0,87,0,72,0,234,0,242,0,243,0,201,0,135,0,0,0,86,0,0,0,217,0,0,0,113,0,0,0,97,0,75,0,174,0,167,0,238,0,177,0,0,0,117,0,117,0,110,0,132,0,61,0,29,0,242,0,47,0,0,0,0,0,117,0,62,0,244,0,0,0,0,0,112,0,50,0,0,0,174,0,18,0,36,0,185,0,168,0,59,0,189,0,64,0,0,0,38,0,237,0,53,0,24,0,0,0,82,0,0,0,0,0,121,0,114,0,128,0,152,0,95,0,90,0,71,0,0,0,123,0,0,0,202,0,26,0,179,0,218,0,0,0,0,0,0,0,169,0,209,0,46,0,62,0,251,0,50,0,0,0,43,0,0,0,104,0,35,0,196,0,71,0,204,0,225,0,138,0,222,0,12,0,204,0,65,0,93,0,85,0,0,0,0,0,65,0,36,0,94,0,249,0,42,0,196,0,33,0,161,0,122,0,168,0,0,0,104,0,137,0,126,0,69,0,9,0,161,0,194,0,142,0,146,0,0,0,101,0,49,0,224,0,165,0,0,0,74,0,107,0,106,0,0,0,192,0,154,0,0,0,103,0,0,0,103,0,0,0,124,0,16,0,227,0,151,0,178,0,188,0,48,0,64,0,10,0,240,0,45,0,195,0,32,0,77,0,191,0,37,0,0,0,172,0,130,0,132,0,35,0,54,0,233,0,0,0,39,0,206,0,235,0,0,0,113,0,209,0,0,0,5,0,14,0,0,0,0,0,96,0,207,0,0,0,192,0,92,0,55,0,239,0,254,0,135,0,123,0,176,0,0,0,146,0,101,0,4,0,21,0,0,0,246,0,168,0,60,0,0,0,0,0,239,0,221,0,235,0,254,0,47,0,155,0,232,0);
signal scenario_full  : scenario_type := (223,31,17,31,85,31,209,31,106,31,42,31,172,31,254,31,181,31,181,30,185,31,71,31,113,31,48,31,48,30,111,31,111,30,111,29,140,31,241,31,4,31,155,31,79,31,233,31,45,31,45,30,45,29,45,28,163,31,163,30,121,31,17,31,17,30,50,31,131,31,66,31,215,31,215,30,85,31,186,31,182,31,56,31,210,31,229,31,63,31,178,31,237,31,31,31,11,31,244,31,149,31,149,30,172,31,200,31,150,31,187,31,187,30,143,31,121,31,121,30,141,31,208,31,38,31,135,31,205,31,167,31,167,30,137,31,21,31,118,31,108,31,52,31,184,31,184,30,184,29,214,31,238,31,13,31,82,31,82,30,189,31,58,31,58,30,39,31,79,31,163,31,162,31,117,31,117,30,250,31,221,31,4,31,69,31,161,31,41,31,169,31,241,31,35,31,45,31,158,31,45,31,14,31,168,31,85,31,85,30,89,31,5,31,103,31,124,31,124,30,195,31,151,31,17,31,234,31,234,30,182,31,211,31,183,31,124,31,197,31,197,30,165,31,241,31,98,31,96,31,96,30,132,31,221,31,178,31,192,31,166,31,88,31,88,30,161,31,238,31,238,30,17,31,10,31,97,31,44,31,90,31,177,31,43,31,9,31,173,31,29,31,167,31,167,30,65,31,65,30,219,31,42,31,43,31,174,31,54,31,46,31,21,31,12,31,12,30,85,31,12,31,12,30,93,31,221,31,160,31,1,31,172,31,46,31,46,30,77,31,28,31,28,30,60,31,60,30,178,31,251,31,251,30,251,29,146,31,116,31,116,30,189,31,180,31,180,30,17,31,237,31,177,31,162,31,162,30,170,31,131,31,131,30,161,31,92,31,82,31,9,31,162,31,174,31,117,31,44,31,30,31,156,31,107,31,243,31,41,31,95,31,33,31,33,30,33,29,225,31,137,31,130,31,130,30,130,29,120,31,87,31,85,31,15,31,120,31,215,31,237,31,103,31,103,30,85,31,152,31,141,31,141,30,141,29,137,31,245,31,230,31,191,31,163,31,18,31,220,31,128,31,98,31,98,30,243,31,74,31,24,31,24,30,158,31,252,31,99,31,15,31,15,30,232,31,161,31,41,31,247,31,225,31,94,31,94,30,124,31,56,31,242,31,215,31,215,30,230,31,8,31,221,31,194,31,89,31,253,31,164,31,77,31,77,30,106,31,74,31,176,31,69,31,138,31,109,31,228,31,179,31,156,31,156,30,101,31,101,30,177,31,177,30,81,31,226,31,226,30,171,31,157,31,126,31,126,30,126,29,163,31,210,31,51,31,51,30,51,29,42,31,37,31,152,31,159,31,215,31,7,31,63,31,63,30,210,31,122,31,97,31,97,30,228,31,220,31,208,31,208,30,208,29,125,31,176,31,176,30,153,31,17,31,86,31,184,31,184,30,202,31,202,30,104,31,8,31,42,31,44,31,44,30,155,31,152,31,26,31,112,31,183,31,120,31,80,31,124,31,189,31,158,31,208,31,19,31,46,31,111,31,79,31,201,31,201,30,140,31,245,31,59,31,124,31,43,31,10,31,180,31,122,31,122,30,136,31,67,31,187,31,7,31,7,30,45,31,81,31,207,31,207,30,55,31,55,30,55,29,219,31,219,30,233,31,91,31,237,31,237,30,184,31,66,31,66,30,79,31,196,31,34,31,34,30,141,31,100,31,140,31,39,31,109,31,109,30,251,31,58,31,58,30,217,31,212,31,212,30,212,29,177,31,213,31,49,31,185,31,185,30,67,31,119,31,119,30,96,31,9,31,15,31,49,31,49,30,49,29,127,31,149,31,149,30,184,31,184,30,184,29,72,31,72,30,145,31,239,31,27,31,186,31,30,31,209,31,185,31,149,31,149,30,149,29,226,31,119,31,219,31,219,30,213,31,233,31,163,31,77,31,187,31,132,31,82,31,82,30,160,31,160,30,101,31,4,31,36,31,134,31,166,31,75,31,196,31,196,30,202,31,57,31,32,31,7,31,184,31,7,31,56,31,56,30,56,29,186,31,2,31,3,31,3,30,3,29,86,31,70,31,179,31,128,31,37,31,21,31,148,31,148,30,148,29,191,31,159,31,36,31,36,30,237,31,252,31,188,31,61,31,61,30,7,31,200,31,167,31,167,30,154,31,61,31,6,31,6,30,158,31,110,31,110,30,243,31,228,31,243,31,183,31,83,31,8,31,193,31,193,30,74,31,126,31,216,31,242,31,242,30,116,31,116,30,116,29,79,31,171,31,206,31,7,31,8,31,140,31,71,31,15,31,29,31,148,31,77,31,116,31,116,30,50,31,50,30,199,31,107,31,107,30,213,31,106,31,48,31,150,31,102,31,182,31,31,31,174,31,32,31,180,31,27,31,8,31,64,31,64,30,221,31,221,30,31,31,45,31,45,30,45,29,58,31,191,31,75,31,39,31,36,31,133,31,138,31,31,31,31,30,199,31,11,31,252,31,58,31,182,31,176,31,47,31,89,31,170,31,91,31,223,31,223,30,78,31,80,31,19,31,159,31,96,31,228,31,55,31,36,31,154,31,154,30,20,31,20,30,20,29,47,31,118,31,11,31,222,31,222,30,189,31,150,31,5,31,233,31,73,31,213,31,35,31,36,31,2,31,8,31,205,31,205,30,100,31,86,31,178,31,178,30,17,31,47,31,159,31,111,31,196,31,117,31,117,30,185,31,185,30,223,31,146,31,21,31,21,30,10,31,10,30,251,31,5,31,35,31,36,31,118,31,118,30,142,31,142,30,216,31,216,30,129,31,103,31,40,31,75,31,199,31,20,31,241,31,125,31,107,31,31,31,48,31,183,31,189,31,130,31,196,31,243,31,53,31,144,31,171,31,159,31,208,31,249,31,135,31,249,31,151,31,77,31,77,30,242,31,242,30,242,29,253,31,114,31,110,31,237,31,237,30,237,29,237,28,105,31,215,31,252,31,24,31,24,30,92,31,54,31,136,31,154,31,22,31,255,31,175,31,220,31,145,31,103,31,251,31,186,31,233,31,244,31,111,31,23,31,217,31,161,31,212,31,92,31,156,31,103,31,103,30,103,29,124,31,90,31,90,30,14,31,57,31,57,30,214,31,2,31,159,31,45,31,197,31,143,31,135,31,135,30,136,31,255,31,255,30,41,31,41,30,194,31,170,31,166,31,175,31,76,31,179,31,99,31,33,31,227,31,227,30,65,31,45,31,120,31,88,31,150,31,214,31,243,31,13,31,13,30,231,31,183,31,183,30,183,29,234,31,16,31,7,31,13,31,13,30,245,31,242,31,53,31,172,31,50,31,18,31,235,31,192,31,212,31,156,31,27,31,98,31,98,30,16,31,129,31,127,31,49,31,115,31,18,31,18,30,4,31,253,31,49,31,162,31,162,30,168,31,149,31,149,30,23,31,205,31,236,31,79,31,93,31,29,31,74,31,66,31,189,31,162,31,144,31,87,31,15,31,91,31,22,31,90,31,175,31,201,31,87,31,72,31,234,31,242,31,243,31,201,31,135,31,135,30,86,31,86,30,217,31,217,30,113,31,113,30,97,31,75,31,174,31,167,31,238,31,177,31,177,30,117,31,117,31,110,31,132,31,61,31,29,31,242,31,47,31,47,30,47,29,117,31,62,31,244,31,244,30,244,29,112,31,50,31,50,30,174,31,18,31,36,31,185,31,168,31,59,31,189,31,64,31,64,30,38,31,237,31,53,31,24,31,24,30,82,31,82,30,82,29,121,31,114,31,128,31,152,31,95,31,90,31,71,31,71,30,123,31,123,30,202,31,26,31,179,31,218,31,218,30,218,29,218,28,169,31,209,31,46,31,62,31,251,31,50,31,50,30,43,31,43,30,104,31,35,31,196,31,71,31,204,31,225,31,138,31,222,31,12,31,204,31,65,31,93,31,85,31,85,30,85,29,65,31,36,31,94,31,249,31,42,31,196,31,33,31,161,31,122,31,168,31,168,30,104,31,137,31,126,31,69,31,9,31,161,31,194,31,142,31,146,31,146,30,101,31,49,31,224,31,165,31,165,30,74,31,107,31,106,31,106,30,192,31,154,31,154,30,103,31,103,30,103,31,103,30,124,31,16,31,227,31,151,31,178,31,188,31,48,31,64,31,10,31,240,31,45,31,195,31,32,31,77,31,191,31,37,31,37,30,172,31,130,31,132,31,35,31,54,31,233,31,233,30,39,31,206,31,235,31,235,30,113,31,209,31,209,30,5,31,14,31,14,30,14,29,96,31,207,31,207,30,192,31,92,31,55,31,239,31,254,31,135,31,123,31,176,31,176,30,146,31,101,31,4,31,21,31,21,30,246,31,168,31,60,31,60,30,60,29,239,31,221,31,235,31,254,31,47,31,155,31,232,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
