-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 566;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (78,0,0,0,104,0,1,0,15,0,0,0,0,0,67,0,0,0,83,0,227,0,120,0,0,0,59,0,216,0,158,0,0,0,161,0,0,0,76,0,57,0,0,0,0,0,122,0,185,0,64,0,189,0,150,0,114,0,66,0,0,0,43,0,253,0,134,0,163,0,0,0,228,0,232,0,224,0,89,0,94,0,38,0,68,0,0,0,0,0,9,0,25,0,207,0,52,0,217,0,54,0,0,0,0,0,0,0,172,0,0,0,147,0,182,0,84,0,238,0,175,0,144,0,199,0,0,0,186,0,0,0,155,0,0,0,128,0,122,0,125,0,104,0,241,0,147,0,72,0,218,0,175,0,222,0,253,0,213,0,135,0,41,0,178,0,222,0,41,0,0,0,21,0,230,0,61,0,113,0,0,0,114,0,71,0,94,0,97,0,141,0,0,0,38,0,182,0,152,0,0,0,92,0,0,0,0,0,133,0,182,0,231,0,178,0,181,0,76,0,51,0,176,0,0,0,95,0,0,0,31,0,160,0,200,0,216,0,40,0,163,0,54,0,18,0,158,0,33,0,55,0,30,0,64,0,130,0,103,0,152,0,119,0,234,0,12,0,0,0,210,0,0,0,159,0,194,0,24,0,134,0,0,0,0,0,63,0,78,0,35,0,77,0,48,0,78,0,139,0,240,0,106,0,191,0,159,0,40,0,0,0,83,0,125,0,68,0,18,0,127,0,204,0,43,0,107,0,0,0,81,0,232,0,219,0,132,0,0,0,154,0,0,0,214,0,16,0,220,0,104,0,0,0,237,0,47,0,231,0,62,0,219,0,78,0,217,0,4,0,98,0,51,0,0,0,179,0,92,0,80,0,125,0,0,0,232,0,41,0,124,0,81,0,149,0,46,0,209,0,0,0,92,0,168,0,0,0,53,0,65,0,93,0,0,0,66,0,178,0,0,0,103,0,0,0,0,0,32,0,9,0,27,0,164,0,231,0,42,0,66,0,117,0,193,0,180,0,0,0,61,0,133,0,74,0,34,0,120,0,0,0,34,0,62,0,5,0,252,0,120,0,201,0,108,0,169,0,0,0,33,0,0,0,204,0,111,0,146,0,23,0,17,0,201,0,30,0,89,0,81,0,27,0,0,0,0,0,213,0,28,0,174,0,184,0,0,0,36,0,158,0,199,0,254,0,0,0,146,0,27,0,186,0,51,0,113,0,0,0,17,0,163,0,248,0,120,0,249,0,216,0,12,0,218,0,60,0,21,0,0,0,0,0,70,0,141,0,0,0,54,0,46,0,0,0,143,0,0,0,210,0,117,0,249,0,0,0,96,0,217,0,247,0,152,0,239,0,231,0,23,0,3,0,37,0,71,0,123,0,0,0,73,0,134,0,100,0,130,0,147,0,187,0,169,0,104,0,112,0,127,0,30,0,85,0,248,0,247,0,211,0,103,0,0,0,92,0,0,0,27,0,1,0,70,0,85,0,150,0,86,0,116,0,196,0,213,0,0,0,204,0,101,0,57,0,128,0,202,0,0,0,202,0,0,0,158,0,95,0,60,0,0,0,60,0,0,0,191,0,22,0,236,0,0,0,243,0,197,0,147,0,167,0,0,0,150,0,61,0,0,0,0,0,0,0,221,0,126,0,0,0,174,0,43,0,0,0,4,0,0,0,189,0,82,0,143,0,236,0,0,0,2,0,71,0,30,0,168,0,0,0,215,0,153,0,157,0,89,0,164,0,72,0,79,0,0,0,0,0,105,0,218,0,0,0,205,0,179,0,187,0,78,0,164,0,212,0,191,0,0,0,65,0,214,0,222,0,85,0,0,0,170,0,139,0,176,0,168,0,77,0,0,0,160,0,101,0,0,0,229,0,224,0,161,0,86,0,246,0,113,0,137,0,188,0,172,0,31,0,0,0,80,0,151,0,56,0,144,0,35,0,225,0,0,0,121,0,69,0,0,0,0,0,187,0,0,0,109,0,0,0,167,0,0,0,23,0,85,0,119,0,114,0,113,0,155,0,137,0,102,0,188,0,26,0,67,0,177,0,51,0,0,0,0,0,38,0,75,0,101,0,249,0,3,0,0,0,193,0,250,0,0,0,173,0,170,0,42,0,0,0,135,0,0,0,170,0,132,0,121,0,174,0,196,0,0,0,76,0,17,0,0,0,8,0,145,0,8,0,96,0,68,0,31,0,85,0,149,0,250,0,255,0,118,0,173,0,109,0,0,0,165,0,100,0,0,0,0,0,205,0,6,0,63,0,146,0,26,0,170,0,199,0,163,0,0,0,229,0,0,0,14,0,130,0,54,0,87,0,86,0,0,0,224,0,255,0,0,0,176,0,0,0,246,0,165,0,184,0,201,0,20,0,0,0,146,0,44,0,97,0,0,0,212,0,106,0,205,0,4,0,0,0,251,0,24,0,24,0,74,0,65,0,79,0,187,0,202,0,0,0,224,0,159,0,243,0,185,0,203,0,0,0,47,0,0,0,0,0,235,0,193,0,53,0,0,0,150,0,25,0,147,0,96,0,0,0,53,0,230,0);
signal scenario_full  : scenario_type := (78,31,78,30,104,31,1,31,15,31,15,30,15,29,67,31,67,30,83,31,227,31,120,31,120,30,59,31,216,31,158,31,158,30,161,31,161,30,76,31,57,31,57,30,57,29,122,31,185,31,64,31,189,31,150,31,114,31,66,31,66,30,43,31,253,31,134,31,163,31,163,30,228,31,232,31,224,31,89,31,94,31,38,31,68,31,68,30,68,29,9,31,25,31,207,31,52,31,217,31,54,31,54,30,54,29,54,28,172,31,172,30,147,31,182,31,84,31,238,31,175,31,144,31,199,31,199,30,186,31,186,30,155,31,155,30,128,31,122,31,125,31,104,31,241,31,147,31,72,31,218,31,175,31,222,31,253,31,213,31,135,31,41,31,178,31,222,31,41,31,41,30,21,31,230,31,61,31,113,31,113,30,114,31,71,31,94,31,97,31,141,31,141,30,38,31,182,31,152,31,152,30,92,31,92,30,92,29,133,31,182,31,231,31,178,31,181,31,76,31,51,31,176,31,176,30,95,31,95,30,31,31,160,31,200,31,216,31,40,31,163,31,54,31,18,31,158,31,33,31,55,31,30,31,64,31,130,31,103,31,152,31,119,31,234,31,12,31,12,30,210,31,210,30,159,31,194,31,24,31,134,31,134,30,134,29,63,31,78,31,35,31,77,31,48,31,78,31,139,31,240,31,106,31,191,31,159,31,40,31,40,30,83,31,125,31,68,31,18,31,127,31,204,31,43,31,107,31,107,30,81,31,232,31,219,31,132,31,132,30,154,31,154,30,214,31,16,31,220,31,104,31,104,30,237,31,47,31,231,31,62,31,219,31,78,31,217,31,4,31,98,31,51,31,51,30,179,31,92,31,80,31,125,31,125,30,232,31,41,31,124,31,81,31,149,31,46,31,209,31,209,30,92,31,168,31,168,30,53,31,65,31,93,31,93,30,66,31,178,31,178,30,103,31,103,30,103,29,32,31,9,31,27,31,164,31,231,31,42,31,66,31,117,31,193,31,180,31,180,30,61,31,133,31,74,31,34,31,120,31,120,30,34,31,62,31,5,31,252,31,120,31,201,31,108,31,169,31,169,30,33,31,33,30,204,31,111,31,146,31,23,31,17,31,201,31,30,31,89,31,81,31,27,31,27,30,27,29,213,31,28,31,174,31,184,31,184,30,36,31,158,31,199,31,254,31,254,30,146,31,27,31,186,31,51,31,113,31,113,30,17,31,163,31,248,31,120,31,249,31,216,31,12,31,218,31,60,31,21,31,21,30,21,29,70,31,141,31,141,30,54,31,46,31,46,30,143,31,143,30,210,31,117,31,249,31,249,30,96,31,217,31,247,31,152,31,239,31,231,31,23,31,3,31,37,31,71,31,123,31,123,30,73,31,134,31,100,31,130,31,147,31,187,31,169,31,104,31,112,31,127,31,30,31,85,31,248,31,247,31,211,31,103,31,103,30,92,31,92,30,27,31,1,31,70,31,85,31,150,31,86,31,116,31,196,31,213,31,213,30,204,31,101,31,57,31,128,31,202,31,202,30,202,31,202,30,158,31,95,31,60,31,60,30,60,31,60,30,191,31,22,31,236,31,236,30,243,31,197,31,147,31,167,31,167,30,150,31,61,31,61,30,61,29,61,28,221,31,126,31,126,30,174,31,43,31,43,30,4,31,4,30,189,31,82,31,143,31,236,31,236,30,2,31,71,31,30,31,168,31,168,30,215,31,153,31,157,31,89,31,164,31,72,31,79,31,79,30,79,29,105,31,218,31,218,30,205,31,179,31,187,31,78,31,164,31,212,31,191,31,191,30,65,31,214,31,222,31,85,31,85,30,170,31,139,31,176,31,168,31,77,31,77,30,160,31,101,31,101,30,229,31,224,31,161,31,86,31,246,31,113,31,137,31,188,31,172,31,31,31,31,30,80,31,151,31,56,31,144,31,35,31,225,31,225,30,121,31,69,31,69,30,69,29,187,31,187,30,109,31,109,30,167,31,167,30,23,31,85,31,119,31,114,31,113,31,155,31,137,31,102,31,188,31,26,31,67,31,177,31,51,31,51,30,51,29,38,31,75,31,101,31,249,31,3,31,3,30,193,31,250,31,250,30,173,31,170,31,42,31,42,30,135,31,135,30,170,31,132,31,121,31,174,31,196,31,196,30,76,31,17,31,17,30,8,31,145,31,8,31,96,31,68,31,31,31,85,31,149,31,250,31,255,31,118,31,173,31,109,31,109,30,165,31,100,31,100,30,100,29,205,31,6,31,63,31,146,31,26,31,170,31,199,31,163,31,163,30,229,31,229,30,14,31,130,31,54,31,87,31,86,31,86,30,224,31,255,31,255,30,176,31,176,30,246,31,165,31,184,31,201,31,20,31,20,30,146,31,44,31,97,31,97,30,212,31,106,31,205,31,4,31,4,30,251,31,24,31,24,31,74,31,65,31,79,31,187,31,202,31,202,30,224,31,159,31,243,31,185,31,203,31,203,30,47,31,47,30,47,29,235,31,193,31,53,31,53,30,150,31,25,31,147,31,96,31,96,30,53,31,230,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
