-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_34 is
end project_tb_34;

architecture project_tb_arch_34 of project_tb_34 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 815;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (104,0,224,0,122,0,77,0,235,0,252,0,210,0,50,0,118,0,227,0,170,0,6,0,202,0,0,0,74,0,222,0,57,0,248,0,164,0,157,0,241,0,89,0,0,0,138,0,24,0,188,0,121,0,60,0,147,0,177,0,112,0,0,0,0,0,78,0,48,0,49,0,184,0,0,0,18,0,245,0,0,0,0,0,0,0,0,0,0,0,234,0,70,0,136,0,214,0,0,0,240,0,65,0,251,0,183,0,144,0,0,0,149,0,0,0,100,0,0,0,242,0,141,0,53,0,140,0,0,0,3,0,245,0,0,0,32,0,244,0,19,0,0,0,51,0,144,0,134,0,152,0,206,0,57,0,0,0,164,0,45,0,162,0,12,0,104,0,170,0,0,0,214,0,49,0,50,0,28,0,0,0,0,0,59,0,18,0,0,0,163,0,127,0,52,0,231,0,34,0,168,0,239,0,54,0,26,0,252,0,64,0,108,0,27,0,81,0,212,0,0,0,133,0,181,0,159,0,0,0,158,0,9,0,0,0,2,0,0,0,112,0,224,0,171,0,84,0,115,0,131,0,0,0,191,0,205,0,225,0,129,0,31,0,0,0,105,0,96,0,52,0,89,0,238,0,97,0,246,0,29,0,88,0,61,0,0,0,144,0,0,0,0,0,237,0,151,0,0,0,154,0,172,0,0,0,96,0,162,0,31,0,29,0,60,0,95,0,109,0,90,0,0,0,0,0,78,0,138,0,10,0,178,0,241,0,35,0,2,0,2,0,35,0,173,0,0,0,162,0,112,0,176,0,111,0,0,0,134,0,0,0,150,0,247,0,195,0,177,0,92,0,55,0,136,0,0,0,97,0,28,0,21,0,214,0,56,0,75,0,9,0,241,0,109,0,137,0,14,0,71,0,0,0,0,0,0,0,220,0,62,0,72,0,110,0,94,0,211,0,57,0,59,0,93,0,54,0,0,0,125,0,32,0,150,0,0,0,177,0,0,0,253,0,185,0,0,0,39,0,0,0,69,0,11,0,49,0,149,0,69,0,129,0,0,0,166,0,176,0,29,0,181,0,0,0,66,0,0,0,7,0,202,0,2,0,161,0,42,0,167,0,162,0,237,0,36,0,57,0,171,0,0,0,214,0,38,0,0,0,142,0,235,0,50,0,0,0,212,0,251,0,140,0,145,0,186,0,52,0,170,0,104,0,94,0,62,0,75,0,187,0,0,0,132,0,0,0,0,0,248,0,180,0,90,0,191,0,196,0,127,0,14,0,234,0,201,0,177,0,213,0,162,0,207,0,171,0,146,0,0,0,0,0,236,0,0,0,231,0,99,0,31,0,83,0,127,0,0,0,3,0,115,0,231,0,0,0,119,0,0,0,0,0,0,0,158,0,35,0,0,0,179,0,217,0,0,0,201,0,19,0,44,0,0,0,0,0,89,0,0,0,254,0,189,0,24,0,87,0,126,0,248,0,98,0,99,0,249,0,14,0,0,0,80,0,154,0,144,0,110,0,89,0,0,0,181,0,0,0,130,0,97,0,83,0,83,0,71,0,206,0,199,0,42,0,31,0,0,0,0,0,14,0,0,0,127,0,0,0,63,0,0,0,0,0,250,0,166,0,95,0,8,0,0,0,60,0,212,0,137,0,0,0,42,0,0,0,174,0,97,0,219,0,25,0,0,0,158,0,238,0,0,0,57,0,169,0,0,0,102,0,118,0,113,0,0,0,41,0,0,0,0,0,61,0,130,0,0,0,21,0,13,0,0,0,60,0,178,0,0,0,242,0,137,0,0,0,0,0,0,0,174,0,51,0,65,0,12,0,206,0,135,0,161,0,228,0,0,0,83,0,137,0,154,0,25,0,147,0,0,0,71,0,79,0,9,0,119,0,215,0,0,0,105,0,65,0,0,0,115,0,133,0,240,0,223,0,133,0,4,0,15,0,216,0,0,0,203,0,54,0,28,0,164,0,137,0,108,0,0,0,213,0,33,0,145,0,238,0,0,0,66,0,162,0,206,0,0,0,205,0,227,0,68,0,231,0,5,0,28,0,79,0,252,0,28,0,255,0,146,0,89,0,45,0,0,0,46,0,0,0,90,0,58,0,4,0,0,0,74,0,108,0,135,0,165,0,159,0,90,0,177,0,181,0,215,0,186,0,207,0,251,0,131,0,100,0,193,0,0,0,0,0,80,0,100,0,144,0,0,0,222,0,210,0,0,0,36,0,88,0,250,0,115,0,103,0,96,0,0,0,126,0,0,0,210,0,215,0,132,0,103,0,115,0,0,0,255,0,238,0,84,0,55,0,123,0,0,0,83,0,109,0,63,0,16,0,110,0,13,0,60,0,138,0,162,0,164,0,188,0,183,0,239,0,81,0,0,0,45,0,10,0,84,0,82,0,71,0,25,0,197,0,209,0,0,0,155,0,211,0,0,0,201,0,0,0,185,0,0,0,42,0,178,0,120,0,91,0,205,0,0,0,10,0,55,0,92,0,138,0,211,0,0,0,152,0,51,0,207,0,122,0,134,0,0,0,233,0,110,0,225,0,210,0,24,0,0,0,4,0,104,0,116,0,6,0,140,0,6,0,134,0,0,0,100,0,142,0,0,0,184,0,174,0,46,0,169,0,48,0,0,0,94,0,93,0,85,0,0,0,165,0,24,0,233,0,0,0,90,0,195,0,5,0,0,0,87,0,244,0,217,0,183,0,46,0,0,0,229,0,172,0,90,0,0,0,205,0,195,0,224,0,69,0,180,0,44,0,241,0,162,0,52,0,13,0,0,0,35,0,0,0,154,0,118,0,113,0,0,0,117,0,204,0,0,0,190,0,50,0,195,0,220,0,243,0,77,0,77,0,171,0,159,0,60,0,121,0,26,0,240,0,221,0,187,0,79,0,87,0,225,0,231,0,220,0,0,0,69,0,66,0,29,0,0,0,119,0,90,0,0,0,23,0,227,0,29,0,0,0,7,0,187,0,204,0,144,0,203,0,56,0,60,0,167,0,83,0,0,0,210,0,29,0,40,0,64,0,0,0,234,0,14,0,83,0,227,0,0,0,71,0,75,0,163,0,94,0,128,0,188,0,250,0,138,0,0,0,218,0,0,0,174,0,79,0,236,0,145,0,46,0,0,0,203,0,0,0,138,0,97,0,128,0,163,0,151,0,0,0,204,0,109,0,168,0,0,0,53,0,210,0,211,0,120,0,0,0,196,0,72,0,124,0,117,0,50,0,71,0,17,0,203,0,18,0,59,0,0,0,151,0,5,0,43,0,39,0,217,0,0,0,189,0,232,0,0,0,249,0,250,0,0,0,232,0,60,0,92,0,220,0,0,0,71,0,16,0,112,0,19,0,102,0,241,0,45,0,232,0,208,0,10,0,191,0,240,0,124,0,51,0,156,0,240,0,197,0,250,0,216,0,1,0,139,0,84,0,253,0,137,0,12,0,242,0,88,0,171,0,228,0,0,0,231,0,235,0,0,0,66,0,121,0,181,0,44,0,169,0,62,0,0,0,239,0,199,0,0,0,0,0,70,0,0,0,217,0,184,0,247,0,152,0,89,0,241,0,0,0,227,0,38,0,134,0,56,0,0,0,56,0,20,0,113,0,104,0,9,0,193,0,0,0,56,0,147,0,235,0,244,0,91,0,84,0,105,0);
signal scenario_full  : scenario_type := (104,31,224,31,122,31,77,31,235,31,252,31,210,31,50,31,118,31,227,31,170,31,6,31,202,31,202,30,74,31,222,31,57,31,248,31,164,31,157,31,241,31,89,31,89,30,138,31,24,31,188,31,121,31,60,31,147,31,177,31,112,31,112,30,112,29,78,31,48,31,49,31,184,31,184,30,18,31,245,31,245,30,245,29,245,28,245,27,245,26,234,31,70,31,136,31,214,31,214,30,240,31,65,31,251,31,183,31,144,31,144,30,149,31,149,30,100,31,100,30,242,31,141,31,53,31,140,31,140,30,3,31,245,31,245,30,32,31,244,31,19,31,19,30,51,31,144,31,134,31,152,31,206,31,57,31,57,30,164,31,45,31,162,31,12,31,104,31,170,31,170,30,214,31,49,31,50,31,28,31,28,30,28,29,59,31,18,31,18,30,163,31,127,31,52,31,231,31,34,31,168,31,239,31,54,31,26,31,252,31,64,31,108,31,27,31,81,31,212,31,212,30,133,31,181,31,159,31,159,30,158,31,9,31,9,30,2,31,2,30,112,31,224,31,171,31,84,31,115,31,131,31,131,30,191,31,205,31,225,31,129,31,31,31,31,30,105,31,96,31,52,31,89,31,238,31,97,31,246,31,29,31,88,31,61,31,61,30,144,31,144,30,144,29,237,31,151,31,151,30,154,31,172,31,172,30,96,31,162,31,31,31,29,31,60,31,95,31,109,31,90,31,90,30,90,29,78,31,138,31,10,31,178,31,241,31,35,31,2,31,2,31,35,31,173,31,173,30,162,31,112,31,176,31,111,31,111,30,134,31,134,30,150,31,247,31,195,31,177,31,92,31,55,31,136,31,136,30,97,31,28,31,21,31,214,31,56,31,75,31,9,31,241,31,109,31,137,31,14,31,71,31,71,30,71,29,71,28,220,31,62,31,72,31,110,31,94,31,211,31,57,31,59,31,93,31,54,31,54,30,125,31,32,31,150,31,150,30,177,31,177,30,253,31,185,31,185,30,39,31,39,30,69,31,11,31,49,31,149,31,69,31,129,31,129,30,166,31,176,31,29,31,181,31,181,30,66,31,66,30,7,31,202,31,2,31,161,31,42,31,167,31,162,31,237,31,36,31,57,31,171,31,171,30,214,31,38,31,38,30,142,31,235,31,50,31,50,30,212,31,251,31,140,31,145,31,186,31,52,31,170,31,104,31,94,31,62,31,75,31,187,31,187,30,132,31,132,30,132,29,248,31,180,31,90,31,191,31,196,31,127,31,14,31,234,31,201,31,177,31,213,31,162,31,207,31,171,31,146,31,146,30,146,29,236,31,236,30,231,31,99,31,31,31,83,31,127,31,127,30,3,31,115,31,231,31,231,30,119,31,119,30,119,29,119,28,158,31,35,31,35,30,179,31,217,31,217,30,201,31,19,31,44,31,44,30,44,29,89,31,89,30,254,31,189,31,24,31,87,31,126,31,248,31,98,31,99,31,249,31,14,31,14,30,80,31,154,31,144,31,110,31,89,31,89,30,181,31,181,30,130,31,97,31,83,31,83,31,71,31,206,31,199,31,42,31,31,31,31,30,31,29,14,31,14,30,127,31,127,30,63,31,63,30,63,29,250,31,166,31,95,31,8,31,8,30,60,31,212,31,137,31,137,30,42,31,42,30,174,31,97,31,219,31,25,31,25,30,158,31,238,31,238,30,57,31,169,31,169,30,102,31,118,31,113,31,113,30,41,31,41,30,41,29,61,31,130,31,130,30,21,31,13,31,13,30,60,31,178,31,178,30,242,31,137,31,137,30,137,29,137,28,174,31,51,31,65,31,12,31,206,31,135,31,161,31,228,31,228,30,83,31,137,31,154,31,25,31,147,31,147,30,71,31,79,31,9,31,119,31,215,31,215,30,105,31,65,31,65,30,115,31,133,31,240,31,223,31,133,31,4,31,15,31,216,31,216,30,203,31,54,31,28,31,164,31,137,31,108,31,108,30,213,31,33,31,145,31,238,31,238,30,66,31,162,31,206,31,206,30,205,31,227,31,68,31,231,31,5,31,28,31,79,31,252,31,28,31,255,31,146,31,89,31,45,31,45,30,46,31,46,30,90,31,58,31,4,31,4,30,74,31,108,31,135,31,165,31,159,31,90,31,177,31,181,31,215,31,186,31,207,31,251,31,131,31,100,31,193,31,193,30,193,29,80,31,100,31,144,31,144,30,222,31,210,31,210,30,36,31,88,31,250,31,115,31,103,31,96,31,96,30,126,31,126,30,210,31,215,31,132,31,103,31,115,31,115,30,255,31,238,31,84,31,55,31,123,31,123,30,83,31,109,31,63,31,16,31,110,31,13,31,60,31,138,31,162,31,164,31,188,31,183,31,239,31,81,31,81,30,45,31,10,31,84,31,82,31,71,31,25,31,197,31,209,31,209,30,155,31,211,31,211,30,201,31,201,30,185,31,185,30,42,31,178,31,120,31,91,31,205,31,205,30,10,31,55,31,92,31,138,31,211,31,211,30,152,31,51,31,207,31,122,31,134,31,134,30,233,31,110,31,225,31,210,31,24,31,24,30,4,31,104,31,116,31,6,31,140,31,6,31,134,31,134,30,100,31,142,31,142,30,184,31,174,31,46,31,169,31,48,31,48,30,94,31,93,31,85,31,85,30,165,31,24,31,233,31,233,30,90,31,195,31,5,31,5,30,87,31,244,31,217,31,183,31,46,31,46,30,229,31,172,31,90,31,90,30,205,31,195,31,224,31,69,31,180,31,44,31,241,31,162,31,52,31,13,31,13,30,35,31,35,30,154,31,118,31,113,31,113,30,117,31,204,31,204,30,190,31,50,31,195,31,220,31,243,31,77,31,77,31,171,31,159,31,60,31,121,31,26,31,240,31,221,31,187,31,79,31,87,31,225,31,231,31,220,31,220,30,69,31,66,31,29,31,29,30,119,31,90,31,90,30,23,31,227,31,29,31,29,30,7,31,187,31,204,31,144,31,203,31,56,31,60,31,167,31,83,31,83,30,210,31,29,31,40,31,64,31,64,30,234,31,14,31,83,31,227,31,227,30,71,31,75,31,163,31,94,31,128,31,188,31,250,31,138,31,138,30,218,31,218,30,174,31,79,31,236,31,145,31,46,31,46,30,203,31,203,30,138,31,97,31,128,31,163,31,151,31,151,30,204,31,109,31,168,31,168,30,53,31,210,31,211,31,120,31,120,30,196,31,72,31,124,31,117,31,50,31,71,31,17,31,203,31,18,31,59,31,59,30,151,31,5,31,43,31,39,31,217,31,217,30,189,31,232,31,232,30,249,31,250,31,250,30,232,31,60,31,92,31,220,31,220,30,71,31,16,31,112,31,19,31,102,31,241,31,45,31,232,31,208,31,10,31,191,31,240,31,124,31,51,31,156,31,240,31,197,31,250,31,216,31,1,31,139,31,84,31,253,31,137,31,12,31,242,31,88,31,171,31,228,31,228,30,231,31,235,31,235,30,66,31,121,31,181,31,44,31,169,31,62,31,62,30,239,31,199,31,199,30,199,29,70,31,70,30,217,31,184,31,247,31,152,31,89,31,241,31,241,30,227,31,38,31,134,31,56,31,56,30,56,31,20,31,113,31,104,31,9,31,193,31,193,30,56,31,147,31,235,31,244,31,91,31,84,31,105,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
