-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 285;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (199,0,101,0,247,0,234,0,75,0,15,0,94,0,114,0,211,0,0,0,184,0,18,0,39,0,167,0,232,0,161,0,151,0,0,0,0,0,4,0,69,0,52,0,1,0,14,0,202,0,168,0,46,0,252,0,245,0,162,0,122,0,50,0,1,0,104,0,0,0,0,0,0,0,159,0,114,0,111,0,253,0,147,0,255,0,236,0,14,0,94,0,130,0,0,0,0,0,62,0,104,0,227,0,254,0,131,0,34,0,251,0,72,0,0,0,126,0,104,0,17,0,204,0,137,0,112,0,46,0,32,0,157,0,0,0,0,0,198,0,229,0,0,0,61,0,228,0,126,0,66,0,20,0,0,0,228,0,37,0,107,0,0,0,63,0,6,0,9,0,0,0,0,0,226,0,82,0,92,0,159,0,191,0,128,0,68,0,63,0,0,0,210,0,100,0,93,0,0,0,203,0,240,0,111,0,152,0,169,0,157,0,0,0,184,0,14,0,125,0,180,0,208,0,0,0,0,0,211,0,136,0,202,0,0,0,44,0,181,0,0,0,205,0,0,0,207,0,226,0,253,0,0,0,128,0,53,0,163,0,0,0,209,0,194,0,0,0,107,0,140,0,160,0,229,0,110,0,61,0,29,0,7,0,172,0,170,0,0,0,0,0,177,0,208,0,93,0,13,0,135,0,7,0,249,0,29,0,73,0,230,0,195,0,200,0,60,0,0,0,195,0,133,0,0,0,0,0,71,0,15,0,125,0,39,0,113,0,63,0,0,0,192,0,53,0,132,0,251,0,55,0,220,0,236,0,225,0,41,0,185,0,0,0,167,0,196,0,112,0,181,0,89,0,110,0,222,0,0,0,0,0,0,0,136,0,0,0,23,0,1,0,28,0,55,0,134,0,104,0,69,0,7,0,17,0,0,0,185,0,23,0,174,0,227,0,133,0,89,0,233,0,233,0,57,0,54,0,32,0,37,0,0,0,0,0,0,0,204,0,0,0,112,0,0,0,51,0,28,0,39,0,4,0,133,0,237,0,242,0,222,0,178,0,186,0,51,0,80,0,107,0,71,0,252,0,135,0,6,0,105,0,97,0,66,0,193,0,0,0,56,0,201,0,0,0,0,0,0,0,92,0,212,0,110,0,0,0,165,0,105,0,0,0,39,0,112,0,0,0,3,0,193,0,0,0,77,0,66,0,8,0,233,0,37,0,85,0,75,0,141,0,0,0,80,0,235,0,0,0,0,0,92,0,144,0,0,0,0,0,170,0,192,0,148,0,109,0,230,0);
signal scenario_full  : scenario_type := (199,31,101,31,247,31,234,31,75,31,15,31,94,31,114,31,211,31,211,30,184,31,18,31,39,31,167,31,232,31,161,31,151,31,151,30,151,29,4,31,69,31,52,31,1,31,14,31,202,31,168,31,46,31,252,31,245,31,162,31,122,31,50,31,1,31,104,31,104,30,104,29,104,28,159,31,114,31,111,31,253,31,147,31,255,31,236,31,14,31,94,31,130,31,130,30,130,29,62,31,104,31,227,31,254,31,131,31,34,31,251,31,72,31,72,30,126,31,104,31,17,31,204,31,137,31,112,31,46,31,32,31,157,31,157,30,157,29,198,31,229,31,229,30,61,31,228,31,126,31,66,31,20,31,20,30,228,31,37,31,107,31,107,30,63,31,6,31,9,31,9,30,9,29,226,31,82,31,92,31,159,31,191,31,128,31,68,31,63,31,63,30,210,31,100,31,93,31,93,30,203,31,240,31,111,31,152,31,169,31,157,31,157,30,184,31,14,31,125,31,180,31,208,31,208,30,208,29,211,31,136,31,202,31,202,30,44,31,181,31,181,30,205,31,205,30,207,31,226,31,253,31,253,30,128,31,53,31,163,31,163,30,209,31,194,31,194,30,107,31,140,31,160,31,229,31,110,31,61,31,29,31,7,31,172,31,170,31,170,30,170,29,177,31,208,31,93,31,13,31,135,31,7,31,249,31,29,31,73,31,230,31,195,31,200,31,60,31,60,30,195,31,133,31,133,30,133,29,71,31,15,31,125,31,39,31,113,31,63,31,63,30,192,31,53,31,132,31,251,31,55,31,220,31,236,31,225,31,41,31,185,31,185,30,167,31,196,31,112,31,181,31,89,31,110,31,222,31,222,30,222,29,222,28,136,31,136,30,23,31,1,31,28,31,55,31,134,31,104,31,69,31,7,31,17,31,17,30,185,31,23,31,174,31,227,31,133,31,89,31,233,31,233,31,57,31,54,31,32,31,37,31,37,30,37,29,37,28,204,31,204,30,112,31,112,30,51,31,28,31,39,31,4,31,133,31,237,31,242,31,222,31,178,31,186,31,51,31,80,31,107,31,71,31,252,31,135,31,6,31,105,31,97,31,66,31,193,31,193,30,56,31,201,31,201,30,201,29,201,28,92,31,212,31,110,31,110,30,165,31,105,31,105,30,39,31,112,31,112,30,3,31,193,31,193,30,77,31,66,31,8,31,233,31,37,31,85,31,75,31,141,31,141,30,80,31,235,31,235,30,235,29,92,31,144,31,144,30,144,29,170,31,192,31,148,31,109,31,230,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
