-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_973 is
end project_tb_973;

architecture project_tb_arch_973 of project_tb_973 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 985;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (40,0,234,0,59,0,172,0,97,0,133,0,228,0,0,0,0,0,162,0,66,0,7,0,90,0,7,0,0,0,0,0,0,0,78,0,0,0,32,0,126,0,113,0,118,0,120,0,0,0,0,0,125,0,11,0,0,0,223,0,99,0,32,0,51,0,0,0,91,0,0,0,44,0,48,0,0,0,48,0,23,0,157,0,125,0,85,0,55,0,0,0,160,0,123,0,89,0,44,0,64,0,0,0,186,0,255,0,18,0,126,0,0,0,0,0,140,0,214,0,115,0,195,0,170,0,0,0,249,0,227,0,28,0,104,0,49,0,0,0,221,0,0,0,253,0,78,0,163,0,44,0,87,0,0,0,251,0,119,0,212,0,71,0,223,0,57,0,0,0,97,0,114,0,183,0,184,0,0,0,164,0,42,0,248,0,0,0,170,0,0,0,229,0,22,0,83,0,168,0,0,0,151,0,0,0,0,0,0,0,0,0,229,0,0,0,163,0,166,0,203,0,0,0,218,0,113,0,109,0,0,0,0,0,236,0,152,0,104,0,68,0,79,0,90,0,196,0,0,0,10,0,50,0,190,0,0,0,146,0,129,0,182,0,221,0,247,0,0,0,237,0,0,0,44,0,0,0,53,0,247,0,216,0,250,0,235,0,128,0,187,0,0,0,11,0,73,0,0,0,97,0,246,0,105,0,0,0,210,0,93,0,145,0,81,0,35,0,0,0,0,0,137,0,138,0,197,0,149,0,26,0,0,0,3,0,177,0,0,0,187,0,117,0,141,0,138,0,115,0,139,0,63,0,1,0,50,0,158,0,87,0,0,0,252,0,0,0,178,0,123,0,247,0,70,0,34,0,86,0,149,0,0,0,0,0,0,0,89,0,82,0,254,0,16,0,193,0,161,0,228,0,0,0,0,0,234,0,164,0,14,0,0,0,21,0,158,0,107,0,193,0,0,0,0,0,12,0,169,0,0,0,0,0,0,0,173,0,29,0,143,0,236,0,155,0,0,0,85,0,38,0,174,0,214,0,114,0,38,0,0,0,0,0,41,0,75,0,3,0,177,0,94,0,106,0,165,0,46,0,0,0,200,0,179,0,108,0,98,0,0,0,0,0,1,0,0,0,110,0,215,0,206,0,165,0,56,0,21,0,119,0,242,0,2,0,0,0,180,0,254,0,128,0,121,0,155,0,95,0,224,0,53,0,228,0,22,0,192,0,0,0,83,0,0,0,13,0,114,0,231,0,224,0,43,0,238,0,0,0,81,0,0,0,186,0,112,0,0,0,165,0,0,0,0,0,17,0,55,0,22,0,106,0,110,0,183,0,0,0,0,0,144,0,3,0,94,0,0,0,183,0,0,0,84,0,169,0,105,0,165,0,124,0,238,0,178,0,4,0,0,0,251,0,50,0,95,0,167,0,0,0,57,0,0,0,164,0,29,0,103,0,0,0,153,0,209,0,193,0,23,0,121,0,190,0,242,0,0,0,129,0,0,0,121,0,44,0,0,0,37,0,85,0,235,0,232,0,103,0,159,0,6,0,215,0,81,0,236,0,175,0,92,0,31,0,35,0,70,0,0,0,49,0,16,0,193,0,92,0,1,0,116,0,117,0,198,0,222,0,177,0,159,0,113,0,98,0,217,0,0,0,148,0,128,0,47,0,159,0,0,0,74,0,163,0,0,0,245,0,56,0,45,0,252,0,158,0,39,0,0,0,108,0,66,0,83,0,143,0,216,0,143,0,198,0,99,0,155,0,193,0,134,0,0,0,191,0,40,0,0,0,228,0,203,0,103,0,96,0,236,0,169,0,0,0,0,0,80,0,0,0,202,0,248,0,87,0,0,0,89,0,0,0,0,0,88,0,76,0,217,0,149,0,71,0,10,0,47,0,220,0,127,0,181,0,225,0,9,0,0,0,110,0,181,0,218,0,67,0,79,0,102,0,0,0,159,0,124,0,157,0,37,0,61,0,93,0,122,0,91,0,164,0,247,0,125,0,142,0,99,0,74,0,44,0,170,0,230,0,139,0,189,0,35,0,63,0,202,0,0,0,37,0,120,0,0,0,148,0,135,0,249,0,155,0,183,0,47,0,214,0,32,0,47,0,242,0,132,0,180,0,140,0,0,0,19,0,156,0,146,0,129,0,0,0,0,0,73,0,245,0,215,0,180,0,132,0,0,0,186,0,5,0,0,0,53,0,127,0,250,0,0,0,126,0,0,0,229,0,129,0,0,0,168,0,127,0,0,0,162,0,0,0,216,0,0,0,0,0,155,0,249,0,68,0,202,0,52,0,103,0,185,0,87,0,0,0,184,0,238,0,0,0,166,0,193,0,75,0,160,0,20,0,100,0,71,0,60,0,134,0,0,0,0,0,234,0,135,0,159,0,0,0,225,0,144,0,203,0,116,0,95,0,124,0,0,0,237,0,166,0,29,0,112,0,140,0,78,0,164,0,0,0,188,0,231,0,0,0,217,0,71,0,0,0,103,0,139,0,120,0,33,0,117,0,209,0,131,0,0,0,25,0,111,0,44,0,66,0,79,0,51,0,231,0,127,0,13,0,0,0,0,0,106,0,0,0,91,0,92,0,11,0,245,0,213,0,0,0,129,0,183,0,0,0,28,0,43,0,0,0,0,0,100,0,145,0,96,0,238,0,247,0,176,0,215,0,52,0,37,0,52,0,117,0,255,0,1,0,146,0,229,0,73,0,58,0,0,0,180,0,171,0,149,0,73,0,181,0,0,0,155,0,167,0,0,0,231,0,0,0,0,0,90,0,249,0,107,0,18,0,40,0,0,0,188,0,0,0,234,0,171,0,12,0,27,0,102,0,175,0,59,0,183,0,195,0,0,0,0,0,246,0,83,0,135,0,0,0,72,0,0,0,200,0,133,0,0,0,128,0,138,0,13,0,0,0,7,0,176,0,217,0,36,0,8,0,0,0,250,0,0,0,0,0,0,0,167,0,0,0,36,0,191,0,65,0,28,0,200,0,163,0,43,0,89,0,28,0,101,0,163,0,1,0,20,0,213,0,67,0,135,0,120,0,193,0,0,0,5,0,217,0,148,0,206,0,216,0,131,0,164,0,242,0,3,0,249,0,163,0,32,0,73,0,0,0,161,0,71,0,93,0,0,0,213,0,34,0,0,0,15,0,238,0,229,0,90,0,209,0,10,0,0,0,17,0,130,0,192,0,72,0,0,0,74,0,0,0,70,0,142,0,210,0,34,0,148,0,0,0,37,0,205,0,15,0,164,0,107,0,252,0,146,0,60,0,22,0,191,0,0,0,167,0,0,0,209,0,205,0,0,0,189,0,178,0,24,0,175,0,182,0,135,0,236,0,139,0,0,0,48,0,156,0,235,0,0,0,0,0,206,0,194,0,232,0,224,0,63,0,35,0,194,0,94,0,251,0,228,0,55,0,202,0,148,0,62,0,0,0,78,0,134,0,106,0,95,0,81,0,72,0,17,0,191,0,26,0,100,0,186,0,22,0,0,0,200,0,0,0,20,0,237,0,146,0,68,0,91,0,19,0,202,0,41,0,73,0,161,0,208,0,147,0,0,0,39,0,0,0,166,0,47,0,83,0,214,0,0,0,15,0,0,0,57,0,171,0,0,0,38,0,133,0,133,0,255,0,223,0,0,0,0,0,147,0,175,0,199,0,0,0,13,0,150,0,55,0,0,0,156,0,181,0,18,0,166,0,125,0,229,0,146,0,238,0,195,0,0,0,25,0,0,0,13,0,93,0,160,0,76,0,23,0,198,0,0,0,170,0,0,0,0,0,162,0,137,0,29,0,242,0,0,0,13,0,44,0,100,0,32,0,233,0,82,0,50,0,195,0,0,0,224,0,57,0,135,0,86,0,31,0,0,0,63,0,97,0,248,0,72,0,172,0,175,0,184,0,103,0,69,0,191,0,47,0,0,0,230,0,0,0,133,0,67,0,103,0,115,0,139,0,208,0,65,0,54,0,138,0,205,0,27,0,203,0,69,0,253,0,0,0,53,0,79,0,145,0,63,0,0,0,174,0,150,0,79,0,250,0,31,0,149,0,119,0,228,0,117,0,93,0,126,0,244,0,113,0,190,0,0,0,127,0,156,0,0,0,66,0,195,0,230,0,164,0,0,0,237,0,116,0,155,0,0,0,92,0,220,0,146,0,0,0,115,0,0,0,191,0,0,0,3,0,0,0,108,0,162,0,137,0,62,0,21,0,203,0,107,0,187,0,0,0,137,0,212,0,139,0,197,0,0,0,0,0,213,0,9,0,92,0,182,0,0,0,83,0,57,0,153,0,115,0,175,0,20,0,222,0,0,0,117,0,186,0,81,0,0,0,0,0,0,0,121,0,154,0,137,0,0,0,5,0,145,0,0,0,166,0,52,0,91,0,213,0,106,0,230,0,58,0,101,0,6,0,53,0);
signal scenario_full  : scenario_type := (40,31,234,31,59,31,172,31,97,31,133,31,228,31,228,30,228,29,162,31,66,31,7,31,90,31,7,31,7,30,7,29,7,28,78,31,78,30,32,31,126,31,113,31,118,31,120,31,120,30,120,29,125,31,11,31,11,30,223,31,99,31,32,31,51,31,51,30,91,31,91,30,44,31,48,31,48,30,48,31,23,31,157,31,125,31,85,31,55,31,55,30,160,31,123,31,89,31,44,31,64,31,64,30,186,31,255,31,18,31,126,31,126,30,126,29,140,31,214,31,115,31,195,31,170,31,170,30,249,31,227,31,28,31,104,31,49,31,49,30,221,31,221,30,253,31,78,31,163,31,44,31,87,31,87,30,251,31,119,31,212,31,71,31,223,31,57,31,57,30,97,31,114,31,183,31,184,31,184,30,164,31,42,31,248,31,248,30,170,31,170,30,229,31,22,31,83,31,168,31,168,30,151,31,151,30,151,29,151,28,151,27,229,31,229,30,163,31,166,31,203,31,203,30,218,31,113,31,109,31,109,30,109,29,236,31,152,31,104,31,68,31,79,31,90,31,196,31,196,30,10,31,50,31,190,31,190,30,146,31,129,31,182,31,221,31,247,31,247,30,237,31,237,30,44,31,44,30,53,31,247,31,216,31,250,31,235,31,128,31,187,31,187,30,11,31,73,31,73,30,97,31,246,31,105,31,105,30,210,31,93,31,145,31,81,31,35,31,35,30,35,29,137,31,138,31,197,31,149,31,26,31,26,30,3,31,177,31,177,30,187,31,117,31,141,31,138,31,115,31,139,31,63,31,1,31,50,31,158,31,87,31,87,30,252,31,252,30,178,31,123,31,247,31,70,31,34,31,86,31,149,31,149,30,149,29,149,28,89,31,82,31,254,31,16,31,193,31,161,31,228,31,228,30,228,29,234,31,164,31,14,31,14,30,21,31,158,31,107,31,193,31,193,30,193,29,12,31,169,31,169,30,169,29,169,28,173,31,29,31,143,31,236,31,155,31,155,30,85,31,38,31,174,31,214,31,114,31,38,31,38,30,38,29,41,31,75,31,3,31,177,31,94,31,106,31,165,31,46,31,46,30,200,31,179,31,108,31,98,31,98,30,98,29,1,31,1,30,110,31,215,31,206,31,165,31,56,31,21,31,119,31,242,31,2,31,2,30,180,31,254,31,128,31,121,31,155,31,95,31,224,31,53,31,228,31,22,31,192,31,192,30,83,31,83,30,13,31,114,31,231,31,224,31,43,31,238,31,238,30,81,31,81,30,186,31,112,31,112,30,165,31,165,30,165,29,17,31,55,31,22,31,106,31,110,31,183,31,183,30,183,29,144,31,3,31,94,31,94,30,183,31,183,30,84,31,169,31,105,31,165,31,124,31,238,31,178,31,4,31,4,30,251,31,50,31,95,31,167,31,167,30,57,31,57,30,164,31,29,31,103,31,103,30,153,31,209,31,193,31,23,31,121,31,190,31,242,31,242,30,129,31,129,30,121,31,44,31,44,30,37,31,85,31,235,31,232,31,103,31,159,31,6,31,215,31,81,31,236,31,175,31,92,31,31,31,35,31,70,31,70,30,49,31,16,31,193,31,92,31,1,31,116,31,117,31,198,31,222,31,177,31,159,31,113,31,98,31,217,31,217,30,148,31,128,31,47,31,159,31,159,30,74,31,163,31,163,30,245,31,56,31,45,31,252,31,158,31,39,31,39,30,108,31,66,31,83,31,143,31,216,31,143,31,198,31,99,31,155,31,193,31,134,31,134,30,191,31,40,31,40,30,228,31,203,31,103,31,96,31,236,31,169,31,169,30,169,29,80,31,80,30,202,31,248,31,87,31,87,30,89,31,89,30,89,29,88,31,76,31,217,31,149,31,71,31,10,31,47,31,220,31,127,31,181,31,225,31,9,31,9,30,110,31,181,31,218,31,67,31,79,31,102,31,102,30,159,31,124,31,157,31,37,31,61,31,93,31,122,31,91,31,164,31,247,31,125,31,142,31,99,31,74,31,44,31,170,31,230,31,139,31,189,31,35,31,63,31,202,31,202,30,37,31,120,31,120,30,148,31,135,31,249,31,155,31,183,31,47,31,214,31,32,31,47,31,242,31,132,31,180,31,140,31,140,30,19,31,156,31,146,31,129,31,129,30,129,29,73,31,245,31,215,31,180,31,132,31,132,30,186,31,5,31,5,30,53,31,127,31,250,31,250,30,126,31,126,30,229,31,129,31,129,30,168,31,127,31,127,30,162,31,162,30,216,31,216,30,216,29,155,31,249,31,68,31,202,31,52,31,103,31,185,31,87,31,87,30,184,31,238,31,238,30,166,31,193,31,75,31,160,31,20,31,100,31,71,31,60,31,134,31,134,30,134,29,234,31,135,31,159,31,159,30,225,31,144,31,203,31,116,31,95,31,124,31,124,30,237,31,166,31,29,31,112,31,140,31,78,31,164,31,164,30,188,31,231,31,231,30,217,31,71,31,71,30,103,31,139,31,120,31,33,31,117,31,209,31,131,31,131,30,25,31,111,31,44,31,66,31,79,31,51,31,231,31,127,31,13,31,13,30,13,29,106,31,106,30,91,31,92,31,11,31,245,31,213,31,213,30,129,31,183,31,183,30,28,31,43,31,43,30,43,29,100,31,145,31,96,31,238,31,247,31,176,31,215,31,52,31,37,31,52,31,117,31,255,31,1,31,146,31,229,31,73,31,58,31,58,30,180,31,171,31,149,31,73,31,181,31,181,30,155,31,167,31,167,30,231,31,231,30,231,29,90,31,249,31,107,31,18,31,40,31,40,30,188,31,188,30,234,31,171,31,12,31,27,31,102,31,175,31,59,31,183,31,195,31,195,30,195,29,246,31,83,31,135,31,135,30,72,31,72,30,200,31,133,31,133,30,128,31,138,31,13,31,13,30,7,31,176,31,217,31,36,31,8,31,8,30,250,31,250,30,250,29,250,28,167,31,167,30,36,31,191,31,65,31,28,31,200,31,163,31,43,31,89,31,28,31,101,31,163,31,1,31,20,31,213,31,67,31,135,31,120,31,193,31,193,30,5,31,217,31,148,31,206,31,216,31,131,31,164,31,242,31,3,31,249,31,163,31,32,31,73,31,73,30,161,31,71,31,93,31,93,30,213,31,34,31,34,30,15,31,238,31,229,31,90,31,209,31,10,31,10,30,17,31,130,31,192,31,72,31,72,30,74,31,74,30,70,31,142,31,210,31,34,31,148,31,148,30,37,31,205,31,15,31,164,31,107,31,252,31,146,31,60,31,22,31,191,31,191,30,167,31,167,30,209,31,205,31,205,30,189,31,178,31,24,31,175,31,182,31,135,31,236,31,139,31,139,30,48,31,156,31,235,31,235,30,235,29,206,31,194,31,232,31,224,31,63,31,35,31,194,31,94,31,251,31,228,31,55,31,202,31,148,31,62,31,62,30,78,31,134,31,106,31,95,31,81,31,72,31,17,31,191,31,26,31,100,31,186,31,22,31,22,30,200,31,200,30,20,31,237,31,146,31,68,31,91,31,19,31,202,31,41,31,73,31,161,31,208,31,147,31,147,30,39,31,39,30,166,31,47,31,83,31,214,31,214,30,15,31,15,30,57,31,171,31,171,30,38,31,133,31,133,31,255,31,223,31,223,30,223,29,147,31,175,31,199,31,199,30,13,31,150,31,55,31,55,30,156,31,181,31,18,31,166,31,125,31,229,31,146,31,238,31,195,31,195,30,25,31,25,30,13,31,93,31,160,31,76,31,23,31,198,31,198,30,170,31,170,30,170,29,162,31,137,31,29,31,242,31,242,30,13,31,44,31,100,31,32,31,233,31,82,31,50,31,195,31,195,30,224,31,57,31,135,31,86,31,31,31,31,30,63,31,97,31,248,31,72,31,172,31,175,31,184,31,103,31,69,31,191,31,47,31,47,30,230,31,230,30,133,31,67,31,103,31,115,31,139,31,208,31,65,31,54,31,138,31,205,31,27,31,203,31,69,31,253,31,253,30,53,31,79,31,145,31,63,31,63,30,174,31,150,31,79,31,250,31,31,31,149,31,119,31,228,31,117,31,93,31,126,31,244,31,113,31,190,31,190,30,127,31,156,31,156,30,66,31,195,31,230,31,164,31,164,30,237,31,116,31,155,31,155,30,92,31,220,31,146,31,146,30,115,31,115,30,191,31,191,30,3,31,3,30,108,31,162,31,137,31,62,31,21,31,203,31,107,31,187,31,187,30,137,31,212,31,139,31,197,31,197,30,197,29,213,31,9,31,92,31,182,31,182,30,83,31,57,31,153,31,115,31,175,31,20,31,222,31,222,30,117,31,186,31,81,31,81,30,81,29,81,28,121,31,154,31,137,31,137,30,5,31,145,31,145,30,166,31,52,31,91,31,213,31,106,31,230,31,58,31,101,31,6,31,53,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
