-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 916;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (77,0,0,0,122,0,94,0,0,0,0,0,50,0,167,0,218,0,155,0,226,0,163,0,157,0,52,0,217,0,234,0,184,0,0,0,75,0,50,0,236,0,34,0,239,0,0,0,21,0,126,0,26,0,194,0,61,0,245,0,29,0,200,0,97,0,57,0,0,0,0,0,47,0,218,0,0,0,1,0,40,0,198,0,239,0,0,0,222,0,129,0,250,0,168,0,153,0,251,0,207,0,30,0,103,0,121,0,126,0,59,0,0,0,220,0,0,0,9,0,111,0,0,0,249,0,18,0,252,0,18,0,146,0,110,0,140,0,8,0,207,0,29,0,186,0,0,0,0,0,164,0,0,0,39,0,106,0,67,0,149,0,118,0,0,0,144,0,190,0,132,0,213,0,33,0,153,0,230,0,0,0,196,0,48,0,0,0,118,0,232,0,68,0,89,0,189,0,236,0,0,0,141,0,0,0,130,0,253,0,238,0,0,0,46,0,149,0,171,0,217,0,1,0,68,0,17,0,0,0,205,0,26,0,0,0,243,0,76,0,56,0,121,0,160,0,109,0,65,0,253,0,130,0,79,0,193,0,0,0,175,0,0,0,0,0,0,0,191,0,71,0,0,0,220,0,0,0,0,0,6,0,216,0,65,0,39,0,89,0,0,0,19,0,0,0,124,0,6,0,51,0,51,0,176,0,76,0,210,0,156,0,222,0,185,0,35,0,124,0,0,0,135,0,56,0,188,0,218,0,6,0,161,0,78,0,11,0,135,0,0,0,79,0,63,0,231,0,22,0,0,0,218,0,0,0,25,0,201,0,0,0,64,0,17,0,44,0,43,0,135,0,7,0,101,0,189,0,0,0,60,0,253,0,56,0,34,0,0,0,235,0,0,0,0,0,131,0,196,0,0,0,88,0,13,0,72,0,176,0,10,0,40,0,185,0,29,0,44,0,0,0,25,0,9,0,28,0,139,0,0,0,119,0,167,0,0,0,101,0,240,0,165,0,34,0,98,0,0,0,27,0,138,0,72,0,0,0,131,0,0,0,171,0,0,0,0,0,236,0,17,0,187,0,162,0,161,0,44,0,63,0,152,0,46,0,28,0,68,0,242,0,0,0,0,0,0,0,0,0,101,0,28,0,38,0,0,0,142,0,249,0,0,0,0,0,0,0,216,0,206,0,195,0,156,0,242,0,82,0,124,0,0,0,0,0,0,0,86,0,0,0,228,0,199,0,0,0,234,0,102,0,33,0,0,0,0,0,0,0,0,0,76,0,132,0,123,0,48,0,57,0,0,0,0,0,134,0,85,0,249,0,15,0,1,0,162,0,13,0,3,0,83,0,15,0,127,0,246,0,72,0,0,0,237,0,0,0,34,0,0,0,0,0,150,0,0,0,16,0,18,0,71,0,76,0,56,0,0,0,37,0,248,0,33,0,203,0,222,0,15,0,12,0,76,0,202,0,0,0,211,0,0,0,68,0,68,0,140,0,0,0,22,0,73,0,39,0,237,0,207,0,6,0,193,0,86,0,0,0,0,0,223,0,217,0,238,0,17,0,0,0,117,0,212,0,250,0,227,0,234,0,126,0,253,0,179,0,157,0,105,0,192,0,161,0,0,0,84,0,0,0,240,0,0,0,156,0,59,0,1,0,189,0,0,0,109,0,79,0,132,0,75,0,209,0,0,0,211,0,44,0,189,0,238,0,0,0,0,0,14,0,30,0,176,0,228,0,6,0,0,0,191,0,181,0,82,0,161,0,152,0,137,0,7,0,14,0,202,0,49,0,56,0,136,0,57,0,0,0,209,0,121,0,169,0,106,0,0,0,198,0,4,0,109,0,0,0,134,0,72,0,141,0,210,0,11,0,56,0,0,0,0,0,48,0,90,0,215,0,154,0,144,0,0,0,0,0,54,0,178,0,89,0,23,0,233,0,231,0,35,0,100,0,117,0,243,0,80,0,133,0,128,0,0,0,158,0,95,0,107,0,0,0,52,0,0,0,103,0,244,0,0,0,252,0,119,0,41,0,55,0,0,0,156,0,181,0,163,0,0,0,143,0,224,0,86,0,0,0,247,0,125,0,46,0,31,0,101,0,59,0,81,0,35,0,34,0,138,0,0,0,0,0,17,0,123,0,228,0,9,0,0,0,221,0,214,0,241,0,0,0,204,0,249,0,165,0,0,0,0,0,33,0,10,0,72,0,26,0,127,0,210,0,103,0,0,0,0,0,197,0,67,0,56,0,212,0,5,0,0,0,0,0,145,0,3,0,0,0,0,0,0,0,152,0,45,0,0,0,140,0,171,0,50,0,48,0,0,0,128,0,157,0,163,0,95,0,99,0,0,0,0,0,119,0,225,0,85,0,155,0,84,0,13,0,41,0,170,0,69,0,255,0,134,0,0,0,0,0,0,0,0,0,38,0,184,0,240,0,133,0,84,0,0,0,28,0,0,0,0,0,99,0,158,0,230,0,146,0,164,0,0,0,84,0,81,0,0,0,0,0,202,0,155,0,233,0,204,0,227,0,0,0,82,0,63,0,16,0,17,0,62,0,238,0,254,0,211,0,0,0,167,0,0,0,205,0,226,0,248,0,153,0,0,0,174,0,0,0,40,0,0,0,113,0,235,0,0,0,76,0,37,0,0,0,64,0,169,0,71,0,4,0,59,0,72,0,0,0,85,0,163,0,176,0,165,0,214,0,188,0,0,0,219,0,108,0,16,0,185,0,252,0,0,0,96,0,212,0,143,0,45,0,122,0,225,0,155,0,151,0,189,0,1,0,54,0,250,0,49,0,5,0,50,0,0,0,227,0,45,0,241,0,2,0,0,0,105,0,68,0,253,0,0,0,105,0,0,0,215,0,218,0,34,0,33,0,240,0,0,0,180,0,74,0,134,0,0,0,54,0,195,0,39,0,128,0,187,0,141,0,0,0,128,0,247,0,122,0,81,0,52,0,0,0,44,0,168,0,148,0,230,0,0,0,1,0,43,0,211,0,5,0,178,0,100,0,242,0,226,0,250,0,137,0,235,0,65,0,48,0,247,0,26,0,67,0,113,0,8,0,180,0,59,0,0,0,62,0,57,0,139,0,54,0,149,0,62,0,229,0,30,0,0,0,55,0,0,0,47,0,39,0,185,0,181,0,0,0,41,0,107,0,23,0,24,0,92,0,227,0,146,0,96,0,194,0,88,0,39,0,0,0,147,0,159,0,86,0,0,0,0,0,0,0,252,0,103,0,241,0,0,0,68,0,0,0,121,0,96,0,147,0,206,0,62,0,198,0,95,0,196,0,144,0,172,0,131,0,0,0,119,0,16,0,0,0,0,0,0,0,116,0,0,0,44,0,74,0,103,0,10,0,237,0,124,0,107,0,0,0,44,0,116,0,9,0,152,0,150,0,83,0,44,0,0,0,240,0,200,0,0,0,29,0,47,0,240,0,99,0,0,0,188,0,100,0,41,0,216,0,132,0,128,0,132,0,89,0,242,0,0,0,172,0,134,0,171,0,44,0,169,0,120,0,10,0,207,0,116,0,155,0,122,0,132,0,203,0,0,0,108,0,52,0,126,0,200,0,208,0,88,0,75,0,207,0,69,0,0,0,253,0,16,0,14,0,0,0,109,0,123,0,0,0,69,0,58,0,18,0,37,0,0,0,175,0,74,0,23,0,69,0,45,0,29,0,0,0,0,0,201,0,102,0,135,0,0,0,194,0,251,0,211,0,89,0,29,0,23,0,0,0,56,0,161,0,255,0,231,0,88,0,0,0,205,0,6,0,138,0,86,0,40,0,128,0,161,0,135,0,135,0,191,0,57,0,190,0,211,0,115,0,5,0,201,0,222,0,254,0,0,0,92,0,144,0,0,0,125,0,153,0,126,0,157,0,130,0,255,0,238,0,156,0,118,0,33,0,208,0,92,0,1,0,206,0,91,0,196,0,2,0,241,0,9,0,0,0,140,0,48,0,0,0,154,0,253,0,234,0,29,0,225,0,113,0,61,0,239,0,0,0,103,0,208,0,52,0,204,0,102,0,0,0,0,0,61,0,254,0,70,0,100,0,0,0,83,0,0,0,0,0,24,0,0,0,60,0,132,0,87,0,0,0,197,0,0,0,26,0);
signal scenario_full  : scenario_type := (77,31,77,30,122,31,94,31,94,30,94,29,50,31,167,31,218,31,155,31,226,31,163,31,157,31,52,31,217,31,234,31,184,31,184,30,75,31,50,31,236,31,34,31,239,31,239,30,21,31,126,31,26,31,194,31,61,31,245,31,29,31,200,31,97,31,57,31,57,30,57,29,47,31,218,31,218,30,1,31,40,31,198,31,239,31,239,30,222,31,129,31,250,31,168,31,153,31,251,31,207,31,30,31,103,31,121,31,126,31,59,31,59,30,220,31,220,30,9,31,111,31,111,30,249,31,18,31,252,31,18,31,146,31,110,31,140,31,8,31,207,31,29,31,186,31,186,30,186,29,164,31,164,30,39,31,106,31,67,31,149,31,118,31,118,30,144,31,190,31,132,31,213,31,33,31,153,31,230,31,230,30,196,31,48,31,48,30,118,31,232,31,68,31,89,31,189,31,236,31,236,30,141,31,141,30,130,31,253,31,238,31,238,30,46,31,149,31,171,31,217,31,1,31,68,31,17,31,17,30,205,31,26,31,26,30,243,31,76,31,56,31,121,31,160,31,109,31,65,31,253,31,130,31,79,31,193,31,193,30,175,31,175,30,175,29,175,28,191,31,71,31,71,30,220,31,220,30,220,29,6,31,216,31,65,31,39,31,89,31,89,30,19,31,19,30,124,31,6,31,51,31,51,31,176,31,76,31,210,31,156,31,222,31,185,31,35,31,124,31,124,30,135,31,56,31,188,31,218,31,6,31,161,31,78,31,11,31,135,31,135,30,79,31,63,31,231,31,22,31,22,30,218,31,218,30,25,31,201,31,201,30,64,31,17,31,44,31,43,31,135,31,7,31,101,31,189,31,189,30,60,31,253,31,56,31,34,31,34,30,235,31,235,30,235,29,131,31,196,31,196,30,88,31,13,31,72,31,176,31,10,31,40,31,185,31,29,31,44,31,44,30,25,31,9,31,28,31,139,31,139,30,119,31,167,31,167,30,101,31,240,31,165,31,34,31,98,31,98,30,27,31,138,31,72,31,72,30,131,31,131,30,171,31,171,30,171,29,236,31,17,31,187,31,162,31,161,31,44,31,63,31,152,31,46,31,28,31,68,31,242,31,242,30,242,29,242,28,242,27,101,31,28,31,38,31,38,30,142,31,249,31,249,30,249,29,249,28,216,31,206,31,195,31,156,31,242,31,82,31,124,31,124,30,124,29,124,28,86,31,86,30,228,31,199,31,199,30,234,31,102,31,33,31,33,30,33,29,33,28,33,27,76,31,132,31,123,31,48,31,57,31,57,30,57,29,134,31,85,31,249,31,15,31,1,31,162,31,13,31,3,31,83,31,15,31,127,31,246,31,72,31,72,30,237,31,237,30,34,31,34,30,34,29,150,31,150,30,16,31,18,31,71,31,76,31,56,31,56,30,37,31,248,31,33,31,203,31,222,31,15,31,12,31,76,31,202,31,202,30,211,31,211,30,68,31,68,31,140,31,140,30,22,31,73,31,39,31,237,31,207,31,6,31,193,31,86,31,86,30,86,29,223,31,217,31,238,31,17,31,17,30,117,31,212,31,250,31,227,31,234,31,126,31,253,31,179,31,157,31,105,31,192,31,161,31,161,30,84,31,84,30,240,31,240,30,156,31,59,31,1,31,189,31,189,30,109,31,79,31,132,31,75,31,209,31,209,30,211,31,44,31,189,31,238,31,238,30,238,29,14,31,30,31,176,31,228,31,6,31,6,30,191,31,181,31,82,31,161,31,152,31,137,31,7,31,14,31,202,31,49,31,56,31,136,31,57,31,57,30,209,31,121,31,169,31,106,31,106,30,198,31,4,31,109,31,109,30,134,31,72,31,141,31,210,31,11,31,56,31,56,30,56,29,48,31,90,31,215,31,154,31,144,31,144,30,144,29,54,31,178,31,89,31,23,31,233,31,231,31,35,31,100,31,117,31,243,31,80,31,133,31,128,31,128,30,158,31,95,31,107,31,107,30,52,31,52,30,103,31,244,31,244,30,252,31,119,31,41,31,55,31,55,30,156,31,181,31,163,31,163,30,143,31,224,31,86,31,86,30,247,31,125,31,46,31,31,31,101,31,59,31,81,31,35,31,34,31,138,31,138,30,138,29,17,31,123,31,228,31,9,31,9,30,221,31,214,31,241,31,241,30,204,31,249,31,165,31,165,30,165,29,33,31,10,31,72,31,26,31,127,31,210,31,103,31,103,30,103,29,197,31,67,31,56,31,212,31,5,31,5,30,5,29,145,31,3,31,3,30,3,29,3,28,152,31,45,31,45,30,140,31,171,31,50,31,48,31,48,30,128,31,157,31,163,31,95,31,99,31,99,30,99,29,119,31,225,31,85,31,155,31,84,31,13,31,41,31,170,31,69,31,255,31,134,31,134,30,134,29,134,28,134,27,38,31,184,31,240,31,133,31,84,31,84,30,28,31,28,30,28,29,99,31,158,31,230,31,146,31,164,31,164,30,84,31,81,31,81,30,81,29,202,31,155,31,233,31,204,31,227,31,227,30,82,31,63,31,16,31,17,31,62,31,238,31,254,31,211,31,211,30,167,31,167,30,205,31,226,31,248,31,153,31,153,30,174,31,174,30,40,31,40,30,113,31,235,31,235,30,76,31,37,31,37,30,64,31,169,31,71,31,4,31,59,31,72,31,72,30,85,31,163,31,176,31,165,31,214,31,188,31,188,30,219,31,108,31,16,31,185,31,252,31,252,30,96,31,212,31,143,31,45,31,122,31,225,31,155,31,151,31,189,31,1,31,54,31,250,31,49,31,5,31,50,31,50,30,227,31,45,31,241,31,2,31,2,30,105,31,68,31,253,31,253,30,105,31,105,30,215,31,218,31,34,31,33,31,240,31,240,30,180,31,74,31,134,31,134,30,54,31,195,31,39,31,128,31,187,31,141,31,141,30,128,31,247,31,122,31,81,31,52,31,52,30,44,31,168,31,148,31,230,31,230,30,1,31,43,31,211,31,5,31,178,31,100,31,242,31,226,31,250,31,137,31,235,31,65,31,48,31,247,31,26,31,67,31,113,31,8,31,180,31,59,31,59,30,62,31,57,31,139,31,54,31,149,31,62,31,229,31,30,31,30,30,55,31,55,30,47,31,39,31,185,31,181,31,181,30,41,31,107,31,23,31,24,31,92,31,227,31,146,31,96,31,194,31,88,31,39,31,39,30,147,31,159,31,86,31,86,30,86,29,86,28,252,31,103,31,241,31,241,30,68,31,68,30,121,31,96,31,147,31,206,31,62,31,198,31,95,31,196,31,144,31,172,31,131,31,131,30,119,31,16,31,16,30,16,29,16,28,116,31,116,30,44,31,74,31,103,31,10,31,237,31,124,31,107,31,107,30,44,31,116,31,9,31,152,31,150,31,83,31,44,31,44,30,240,31,200,31,200,30,29,31,47,31,240,31,99,31,99,30,188,31,100,31,41,31,216,31,132,31,128,31,132,31,89,31,242,31,242,30,172,31,134,31,171,31,44,31,169,31,120,31,10,31,207,31,116,31,155,31,122,31,132,31,203,31,203,30,108,31,52,31,126,31,200,31,208,31,88,31,75,31,207,31,69,31,69,30,253,31,16,31,14,31,14,30,109,31,123,31,123,30,69,31,58,31,18,31,37,31,37,30,175,31,74,31,23,31,69,31,45,31,29,31,29,30,29,29,201,31,102,31,135,31,135,30,194,31,251,31,211,31,89,31,29,31,23,31,23,30,56,31,161,31,255,31,231,31,88,31,88,30,205,31,6,31,138,31,86,31,40,31,128,31,161,31,135,31,135,31,191,31,57,31,190,31,211,31,115,31,5,31,201,31,222,31,254,31,254,30,92,31,144,31,144,30,125,31,153,31,126,31,157,31,130,31,255,31,238,31,156,31,118,31,33,31,208,31,92,31,1,31,206,31,91,31,196,31,2,31,241,31,9,31,9,30,140,31,48,31,48,30,154,31,253,31,234,31,29,31,225,31,113,31,61,31,239,31,239,30,103,31,208,31,52,31,204,31,102,31,102,30,102,29,61,31,254,31,70,31,100,31,100,30,83,31,83,30,83,29,24,31,24,30,60,31,132,31,87,31,87,30,197,31,197,30,26,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
