-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_457 is
end project_tb_457;

architecture project_tb_arch_457 of project_tb_457 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 442;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,142,0,175,0,0,0,139,0,55,0,149,0,178,0,74,0,246,0,161,0,202,0,218,0,233,0,176,0,243,0,184,0,0,0,34,0,135,0,52,0,0,0,135,0,89,0,28,0,93,0,197,0,104,0,216,0,105,0,93,0,107,0,170,0,38,0,116,0,240,0,59,0,0,0,120,0,21,0,103,0,229,0,105,0,0,0,130,0,62,0,215,0,250,0,205,0,161,0,96,0,0,0,0,0,35,0,208,0,166,0,0,0,0,0,176,0,0,0,129,0,127,0,0,0,222,0,39,0,0,0,0,0,51,0,179,0,92,0,0,0,0,0,15,0,0,0,66,0,195,0,226,0,238,0,113,0,0,0,0,0,160,0,143,0,156,0,29,0,252,0,206,0,0,0,210,0,71,0,0,0,47,0,169,0,142,0,113,0,81,0,25,0,0,0,169,0,32,0,254,0,14,0,222,0,0,0,84,0,49,0,145,0,168,0,200,0,0,0,86,0,0,0,0,0,188,0,184,0,0,0,76,0,204,0,163,0,130,0,222,0,159,0,95,0,206,0,97,0,217,0,0,0,185,0,210,0,0,0,168,0,136,0,178,0,80,0,13,0,161,0,0,0,0,0,48,0,214,0,104,0,41,0,31,0,47,0,32,0,0,0,24,0,103,0,88,0,20,0,0,0,26,0,254,0,0,0,227,0,153,0,56,0,106,0,24,0,185,0,249,0,8,0,200,0,247,0,249,0,0,0,145,0,131,0,16,0,133,0,83,0,0,0,0,0,0,0,254,0,74,0,195,0,238,0,0,0,255,0,145,0,0,0,110,0,0,0,0,0,18,0,60,0,187,0,124,0,0,0,0,0,48,0,3,0,46,0,116,0,0,0,197,0,196,0,107,0,175,0,14,0,168,0,53,0,38,0,97,0,172,0,245,0,0,0,110,0,136,0,0,0,60,0,88,0,224,0,208,0,40,0,9,0,46,0,125,0,163,0,0,0,21,0,148,0,58,0,0,0,172,0,28,0,63,0,76,0,0,0,0,0,0,0,0,0,55,0,0,0,0,0,0,0,0,0,221,0,200,0,14,0,145,0,0,0,0,0,154,0,136,0,116,0,0,0,162,0,29,0,93,0,142,0,218,0,54,0,0,0,10,0,218,0,0,0,18,0,47,0,136,0,0,0,0,0,0,0,186,0,107,0,47,0,240,0,130,0,40,0,0,0,198,0,192,0,69,0,0,0,55,0,239,0,167,0,0,0,0,0,0,0,0,0,233,0,0,0,228,0,218,0,124,0,0,0,120,0,0,0,10,0,58,0,0,0,251,0,154,0,134,0,0,0,0,0,60,0,98,0,106,0,127,0,208,0,153,0,188,0,0,0,182,0,25,0,193,0,215,0,237,0,200,0,147,0,127,0,135,0,199,0,7,0,31,0,5,0,21,0,246,0,233,0,146,0,112,0,0,0,0,0,230,0,106,0,87,0,229,0,210,0,185,0,0,0,80,0,229,0,32,0,42,0,19,0,80,0,91,0,1,0,0,0,43,0,48,0,53,0,0,0,205,0,187,0,0,0,0,0,68,0,7,0,0,0,101,0,182,0,74,0,145,0,149,0,0,0,0,0,166,0,208,0,255,0,51,0,92,0,0,0,0,0,198,0,0,0,122,0,7,0,136,0,51,0,186,0,230,0,155,0,214,0,73,0,0,0,154,0,0,0,254,0,0,0,64,0,23,0,239,0,32,0,21,0,181,0,0,0,0,0,240,0,202,0,18,0,103,0,221,0,145,0,0,0,89,0,30,0,88,0,186,0,0,0,139,0,0,0,0,0,129,0,65,0,44,0,48,0,47,0,120,0,113,0,245,0,0,0,216,0,110,0,58,0,19,0,93,0,200,0,159,0,130,0,237,0,0,0,0,0,142,0,39,0,21,0,0,0,255,0,192,0,226,0,229,0,7,0,0,0,240,0,0,0,101,0,213,0,0,0);
signal scenario_full  : scenario_type := (0,0,0,0,142,31,175,31,175,30,139,31,55,31,149,31,178,31,74,31,246,31,161,31,202,31,218,31,233,31,176,31,243,31,184,31,184,30,34,31,135,31,52,31,52,30,135,31,89,31,28,31,93,31,197,31,104,31,216,31,105,31,93,31,107,31,170,31,38,31,116,31,240,31,59,31,59,30,120,31,21,31,103,31,229,31,105,31,105,30,130,31,62,31,215,31,250,31,205,31,161,31,96,31,96,30,96,29,35,31,208,31,166,31,166,30,166,29,176,31,176,30,129,31,127,31,127,30,222,31,39,31,39,30,39,29,51,31,179,31,92,31,92,30,92,29,15,31,15,30,66,31,195,31,226,31,238,31,113,31,113,30,113,29,160,31,143,31,156,31,29,31,252,31,206,31,206,30,210,31,71,31,71,30,47,31,169,31,142,31,113,31,81,31,25,31,25,30,169,31,32,31,254,31,14,31,222,31,222,30,84,31,49,31,145,31,168,31,200,31,200,30,86,31,86,30,86,29,188,31,184,31,184,30,76,31,204,31,163,31,130,31,222,31,159,31,95,31,206,31,97,31,217,31,217,30,185,31,210,31,210,30,168,31,136,31,178,31,80,31,13,31,161,31,161,30,161,29,48,31,214,31,104,31,41,31,31,31,47,31,32,31,32,30,24,31,103,31,88,31,20,31,20,30,26,31,254,31,254,30,227,31,153,31,56,31,106,31,24,31,185,31,249,31,8,31,200,31,247,31,249,31,249,30,145,31,131,31,16,31,133,31,83,31,83,30,83,29,83,28,254,31,74,31,195,31,238,31,238,30,255,31,145,31,145,30,110,31,110,30,110,29,18,31,60,31,187,31,124,31,124,30,124,29,48,31,3,31,46,31,116,31,116,30,197,31,196,31,107,31,175,31,14,31,168,31,53,31,38,31,97,31,172,31,245,31,245,30,110,31,136,31,136,30,60,31,88,31,224,31,208,31,40,31,9,31,46,31,125,31,163,31,163,30,21,31,148,31,58,31,58,30,172,31,28,31,63,31,76,31,76,30,76,29,76,28,76,27,55,31,55,30,55,29,55,28,55,27,221,31,200,31,14,31,145,31,145,30,145,29,154,31,136,31,116,31,116,30,162,31,29,31,93,31,142,31,218,31,54,31,54,30,10,31,218,31,218,30,18,31,47,31,136,31,136,30,136,29,136,28,186,31,107,31,47,31,240,31,130,31,40,31,40,30,198,31,192,31,69,31,69,30,55,31,239,31,167,31,167,30,167,29,167,28,167,27,233,31,233,30,228,31,218,31,124,31,124,30,120,31,120,30,10,31,58,31,58,30,251,31,154,31,134,31,134,30,134,29,60,31,98,31,106,31,127,31,208,31,153,31,188,31,188,30,182,31,25,31,193,31,215,31,237,31,200,31,147,31,127,31,135,31,199,31,7,31,31,31,5,31,21,31,246,31,233,31,146,31,112,31,112,30,112,29,230,31,106,31,87,31,229,31,210,31,185,31,185,30,80,31,229,31,32,31,42,31,19,31,80,31,91,31,1,31,1,30,43,31,48,31,53,31,53,30,205,31,187,31,187,30,187,29,68,31,7,31,7,30,101,31,182,31,74,31,145,31,149,31,149,30,149,29,166,31,208,31,255,31,51,31,92,31,92,30,92,29,198,31,198,30,122,31,7,31,136,31,51,31,186,31,230,31,155,31,214,31,73,31,73,30,154,31,154,30,254,31,254,30,64,31,23,31,239,31,32,31,21,31,181,31,181,30,181,29,240,31,202,31,18,31,103,31,221,31,145,31,145,30,89,31,30,31,88,31,186,31,186,30,139,31,139,30,139,29,129,31,65,31,44,31,48,31,47,31,120,31,113,31,245,31,245,30,216,31,110,31,58,31,19,31,93,31,200,31,159,31,130,31,237,31,237,30,237,29,142,31,39,31,21,31,21,30,255,31,192,31,226,31,229,31,7,31,7,30,240,31,240,30,101,31,213,31,213,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
