-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_103 is
end project_tb_103;

architecture project_tb_arch_103 of project_tb_103 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 627;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (33,0,0,0,61,0,244,0,96,0,6,0,230,0,61,0,71,0,0,0,0,0,170,0,221,0,0,0,129,0,155,0,77,0,155,0,86,0,0,0,10,0,200,0,189,0,92,0,213,0,43,0,89,0,0,0,252,0,130,0,0,0,154,0,0,0,35,0,2,0,0,0,31,0,94,0,123,0,38,0,239,0,0,0,55,0,245,0,20,0,0,0,251,0,231,0,0,0,0,0,0,0,147,0,0,0,233,0,89,0,0,0,41,0,48,0,17,0,125,0,28,0,0,0,100,0,51,0,123,0,0,0,239,0,155,0,174,0,137,0,123,0,241,0,58,0,161,0,50,0,87,0,105,0,196,0,13,0,0,0,165,0,232,0,225,0,202,0,153,0,199,0,201,0,182,0,36,0,24,0,138,0,176,0,0,0,194,0,98,0,192,0,0,0,122,0,24,0,0,0,146,0,13,0,76,0,88,0,213,0,63,0,196,0,243,0,169,0,90,0,0,0,197,0,173,0,0,0,117,0,211,0,0,0,206,0,97,0,0,0,0,0,158,0,165,0,161,0,48,0,36,0,177,0,44,0,0,0,147,0,181,0,95,0,129,0,0,0,197,0,20,0,202,0,68,0,0,0,193,0,166,0,16,0,135,0,21,0,178,0,0,0,146,0,116,0,56,0,95,0,0,0,150,0,138,0,200,0,87,0,147,0,222,0,150,0,217,0,0,0,196,0,0,0,114,0,253,0,149,0,203,0,42,0,0,0,233,0,0,0,145,0,112,0,205,0,29,0,0,0,60,0,97,0,0,0,136,0,29,0,224,0,172,0,182,0,129,0,5,0,140,0,51,0,252,0,76,0,236,0,240,0,14,0,0,0,198,0,96,0,16,0,57,0,53,0,242,0,0,0,228,0,186,0,0,0,0,0,178,0,59,0,44,0,168,0,240,0,213,0,25,0,180,0,0,0,132,0,0,0,0,0,248,0,253,0,183,0,0,0,40,0,73,0,91,0,19,0,84,0,222,0,71,0,30,0,66,0,82,0,78,0,211,0,180,0,166,0,230,0,22,0,114,0,70,0,153,0,45,0,81,0,223,0,0,0,15,0,86,0,81,0,209,0,169,0,73,0,172,0,188,0,123,0,0,0,78,0,123,0,0,0,3,0,0,0,0,0,224,0,0,0,148,0,0,0,33,0,81,0,189,0,236,0,177,0,156,0,1,0,0,0,0,0,165,0,212,0,215,0,0,0,221,0,138,0,237,0,0,0,23,0,92,0,169,0,133,0,24,0,160,0,255,0,100,0,0,0,166,0,49,0,154,0,191,0,0,0,68,0,142,0,206,0,151,0,17,0,92,0,0,0,201,0,35,0,153,0,139,0,110,0,199,0,227,0,0,0,87,0,0,0,207,0,231,0,204,0,0,0,54,0,96,0,0,0,0,0,98,0,0,0,197,0,0,0,164,0,50,0,59,0,149,0,57,0,7,0,140,0,204,0,195,0,9,0,187,0,110,0,54,0,209,0,173,0,134,0,163,0,246,0,44,0,165,0,130,0,0,0,228,0,72,0,88,0,20,0,168,0,74,0,80,0,35,0,180,0,248,0,174,0,119,0,187,0,114,0,120,0,218,0,212,0,40,0,73,0,195,0,85,0,214,0,199,0,81,0,147,0,172,0,0,0,27,0,113,0,0,0,0,0,123,0,222,0,0,0,179,0,114,0,234,0,213,0,89,0,143,0,191,0,95,0,0,0,71,0,137,0,0,0,0,0,0,0,119,0,20,0,105,0,78,0,0,0,0,0,181,0,221,0,161,0,245,0,104,0,1,0,91,0,121,0,93,0,193,0,234,0,0,0,249,0,18,0,143,0,10,0,239,0,59,0,60,0,0,0,237,0,41,0,71,0,128,0,0,0,61,0,40,0,127,0,0,0,39,0,139,0,221,0,210,0,112,0,0,0,159,0,253,0,136,0,148,0,125,0,0,0,223,0,0,0,30,0,47,0,231,0,0,0,95,0,0,0,249,0,240,0,176,0,169,0,0,0,0,0,0,0,180,0,176,0,245,0,11,0,245,0,185,0,0,0,164,0,66,0,249,0,213,0,207,0,0,0,0,0,0,0,52,0,127,0,61,0,0,0,0,0,244,0,0,0,192,0,17,0,222,0,230,0,153,0,0,0,115,0,108,0,132,0,175,0,187,0,180,0,0,0,215,0,44,0,100,0,17,0,181,0,5,0,89,0,0,0,82,0,182,0,80,0,198,0,242,0,0,0,0,0,27,0,210,0,68,0,159,0,156,0,120,0,0,0,229,0,217,0,226,0,56,0,231,0,180,0,252,0,29,0,235,0,190,0,0,0,197,0,252,0,0,0,234,0,0,0,19,0,0,0,70,0,183,0,14,0,254,0,74,0,206,0,232,0,233,0,0,0,153,0,214,0,197,0,249,0,142,0,236,0,0,0,63,0,235,0,27,0,0,0,172,0,225,0,240,0,238,0,126,0,0,0,0,0,205,0,66,0,33,0,144,0,0,0,238,0,233,0,0,0,106,0,52,0,48,0,51,0,160,0,121,0,44,0,131,0,201,0,151,0,85,0,232,0,82,0,105,0,0,0,248,0,205,0,10,0,244,0,246,0,37,0,0,0,0,0,230,0,38,0,0,0,245,0,0,0,201,0,182,0,23,0,0,0,0,0,38,0,234,0,237,0,46,0,152,0,209,0,46,0,212,0,0,0,200,0,73,0,0,0,30,0,243,0,66,0,0,0,169,0,140,0,217,0,33,0,118,0,220,0,230,0,251,0,0,0,119,0,207,0,197,0,119,0);
signal scenario_full  : scenario_type := (33,31,33,30,61,31,244,31,96,31,6,31,230,31,61,31,71,31,71,30,71,29,170,31,221,31,221,30,129,31,155,31,77,31,155,31,86,31,86,30,10,31,200,31,189,31,92,31,213,31,43,31,89,31,89,30,252,31,130,31,130,30,154,31,154,30,35,31,2,31,2,30,31,31,94,31,123,31,38,31,239,31,239,30,55,31,245,31,20,31,20,30,251,31,231,31,231,30,231,29,231,28,147,31,147,30,233,31,89,31,89,30,41,31,48,31,17,31,125,31,28,31,28,30,100,31,51,31,123,31,123,30,239,31,155,31,174,31,137,31,123,31,241,31,58,31,161,31,50,31,87,31,105,31,196,31,13,31,13,30,165,31,232,31,225,31,202,31,153,31,199,31,201,31,182,31,36,31,24,31,138,31,176,31,176,30,194,31,98,31,192,31,192,30,122,31,24,31,24,30,146,31,13,31,76,31,88,31,213,31,63,31,196,31,243,31,169,31,90,31,90,30,197,31,173,31,173,30,117,31,211,31,211,30,206,31,97,31,97,30,97,29,158,31,165,31,161,31,48,31,36,31,177,31,44,31,44,30,147,31,181,31,95,31,129,31,129,30,197,31,20,31,202,31,68,31,68,30,193,31,166,31,16,31,135,31,21,31,178,31,178,30,146,31,116,31,56,31,95,31,95,30,150,31,138,31,200,31,87,31,147,31,222,31,150,31,217,31,217,30,196,31,196,30,114,31,253,31,149,31,203,31,42,31,42,30,233,31,233,30,145,31,112,31,205,31,29,31,29,30,60,31,97,31,97,30,136,31,29,31,224,31,172,31,182,31,129,31,5,31,140,31,51,31,252,31,76,31,236,31,240,31,14,31,14,30,198,31,96,31,16,31,57,31,53,31,242,31,242,30,228,31,186,31,186,30,186,29,178,31,59,31,44,31,168,31,240,31,213,31,25,31,180,31,180,30,132,31,132,30,132,29,248,31,253,31,183,31,183,30,40,31,73,31,91,31,19,31,84,31,222,31,71,31,30,31,66,31,82,31,78,31,211,31,180,31,166,31,230,31,22,31,114,31,70,31,153,31,45,31,81,31,223,31,223,30,15,31,86,31,81,31,209,31,169,31,73,31,172,31,188,31,123,31,123,30,78,31,123,31,123,30,3,31,3,30,3,29,224,31,224,30,148,31,148,30,33,31,81,31,189,31,236,31,177,31,156,31,1,31,1,30,1,29,165,31,212,31,215,31,215,30,221,31,138,31,237,31,237,30,23,31,92,31,169,31,133,31,24,31,160,31,255,31,100,31,100,30,166,31,49,31,154,31,191,31,191,30,68,31,142,31,206,31,151,31,17,31,92,31,92,30,201,31,35,31,153,31,139,31,110,31,199,31,227,31,227,30,87,31,87,30,207,31,231,31,204,31,204,30,54,31,96,31,96,30,96,29,98,31,98,30,197,31,197,30,164,31,50,31,59,31,149,31,57,31,7,31,140,31,204,31,195,31,9,31,187,31,110,31,54,31,209,31,173,31,134,31,163,31,246,31,44,31,165,31,130,31,130,30,228,31,72,31,88,31,20,31,168,31,74,31,80,31,35,31,180,31,248,31,174,31,119,31,187,31,114,31,120,31,218,31,212,31,40,31,73,31,195,31,85,31,214,31,199,31,81,31,147,31,172,31,172,30,27,31,113,31,113,30,113,29,123,31,222,31,222,30,179,31,114,31,234,31,213,31,89,31,143,31,191,31,95,31,95,30,71,31,137,31,137,30,137,29,137,28,119,31,20,31,105,31,78,31,78,30,78,29,181,31,221,31,161,31,245,31,104,31,1,31,91,31,121,31,93,31,193,31,234,31,234,30,249,31,18,31,143,31,10,31,239,31,59,31,60,31,60,30,237,31,41,31,71,31,128,31,128,30,61,31,40,31,127,31,127,30,39,31,139,31,221,31,210,31,112,31,112,30,159,31,253,31,136,31,148,31,125,31,125,30,223,31,223,30,30,31,47,31,231,31,231,30,95,31,95,30,249,31,240,31,176,31,169,31,169,30,169,29,169,28,180,31,176,31,245,31,11,31,245,31,185,31,185,30,164,31,66,31,249,31,213,31,207,31,207,30,207,29,207,28,52,31,127,31,61,31,61,30,61,29,244,31,244,30,192,31,17,31,222,31,230,31,153,31,153,30,115,31,108,31,132,31,175,31,187,31,180,31,180,30,215,31,44,31,100,31,17,31,181,31,5,31,89,31,89,30,82,31,182,31,80,31,198,31,242,31,242,30,242,29,27,31,210,31,68,31,159,31,156,31,120,31,120,30,229,31,217,31,226,31,56,31,231,31,180,31,252,31,29,31,235,31,190,31,190,30,197,31,252,31,252,30,234,31,234,30,19,31,19,30,70,31,183,31,14,31,254,31,74,31,206,31,232,31,233,31,233,30,153,31,214,31,197,31,249,31,142,31,236,31,236,30,63,31,235,31,27,31,27,30,172,31,225,31,240,31,238,31,126,31,126,30,126,29,205,31,66,31,33,31,144,31,144,30,238,31,233,31,233,30,106,31,52,31,48,31,51,31,160,31,121,31,44,31,131,31,201,31,151,31,85,31,232,31,82,31,105,31,105,30,248,31,205,31,10,31,244,31,246,31,37,31,37,30,37,29,230,31,38,31,38,30,245,31,245,30,201,31,182,31,23,31,23,30,23,29,38,31,234,31,237,31,46,31,152,31,209,31,46,31,212,31,212,30,200,31,73,31,73,30,30,31,243,31,66,31,66,30,169,31,140,31,217,31,33,31,118,31,220,31,230,31,251,31,251,30,119,31,207,31,197,31,119,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
