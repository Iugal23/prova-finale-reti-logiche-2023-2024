-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 625;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (96,0,0,0,247,0,0,0,0,0,0,0,189,0,228,0,122,0,0,0,96,0,199,0,101,0,124,0,90,0,185,0,0,0,9,0,188,0,0,0,124,0,110,0,44,0,23,0,209,0,64,0,183,0,112,0,244,0,0,0,0,0,79,0,112,0,188,0,106,0,131,0,62,0,0,0,112,0,0,0,184,0,179,0,62,0,199,0,151,0,122,0,102,0,63,0,28,0,210,0,241,0,198,0,240,0,188,0,158,0,143,0,0,0,244,0,55,0,226,0,0,0,132,0,131,0,0,0,173,0,240,0,60,0,141,0,218,0,0,0,140,0,80,0,179,0,72,0,48,0,62,0,22,0,178,0,204,0,73,0,121,0,0,0,0,0,26,0,255,0,118,0,0,0,0,0,17,0,0,0,6,0,82,0,21,0,186,0,0,0,21,0,1,0,233,0,0,0,0,0,64,0,237,0,183,0,163,0,93,0,55,0,194,0,27,0,0,0,124,0,0,0,0,0,0,0,2,0,19,0,252,0,0,0,50,0,106,0,178,0,228,0,81,0,98,0,124,0,2,0,127,0,246,0,223,0,253,0,242,0,133,0,0,0,98,0,32,0,75,0,86,0,0,0,0,0,197,0,0,0,236,0,101,0,27,0,78,0,196,0,149,0,49,0,248,0,229,0,155,0,210,0,171,0,221,0,147,0,11,0,124,0,225,0,186,0,0,0,61,0,49,0,0,0,116,0,169,0,170,0,195,0,93,0,119,0,237,0,0,0,163,0,102,0,170,0,226,0,73,0,0,0,28,0,76,0,0,0,4,0,77,0,0,0,208,0,193,0,59,0,192,0,23,0,178,0,77,0,246,0,97,0,0,0,239,0,27,0,180,0,238,0,122,0,227,0,236,0,171,0,1,0,243,0,0,0,130,0,0,0,147,0,24,0,26,0,19,0,133,0,45,0,133,0,2,0,160,0,0,0,188,0,222,0,83,0,0,0,0,0,181,0,152,0,107,0,66,0,129,0,34,0,202,0,61,0,166,0,195,0,43,0,98,0,53,0,86,0,49,0,238,0,103,0,164,0,32,0,185,0,81,0,243,0,0,0,95,0,55,0,59,0,0,0,20,0,176,0,109,0,250,0,128,0,179,0,168,0,199,0,224,0,203,0,244,0,190,0,88,0,0,0,54,0,3,0,41,0,30,0,220,0,197,0,73,0,246,0,0,0,239,0,35,0,93,0,202,0,0,0,17,0,219,0,109,0,226,0,0,0,193,0,61,0,193,0,5,0,200,0,116,0,176,0,146,0,36,0,0,0,127,0,0,0,57,0,0,0,48,0,82,0,0,0,136,0,193,0,13,0,252,0,76,0,0,0,3,0,48,0,236,0,201,0,129,0,125,0,39,0,84,0,180,0,0,0,171,0,137,0,40,0,198,0,41,0,143,0,77,0,88,0,184,0,243,0,0,0,252,0,236,0,0,0,0,0,202,0,48,0,161,0,0,0,142,0,57,0,221,0,190,0,89,0,191,0,214,0,0,0,211,0,35,0,197,0,254,0,0,0,14,0,85,0,197,0,91,0,181,0,236,0,114,0,78,0,147,0,136,0,225,0,0,0,0,0,23,0,67,0,17,0,138,0,0,0,2,0,65,0,222,0,44,0,0,0,67,0,209,0,26,0,157,0,194,0,187,0,230,0,169,0,0,0,11,0,165,0,0,0,216,0,148,0,29,0,19,0,102,0,32,0,55,0,38,0,34,0,194,0,228,0,49,0,149,0,206,0,70,0,8,0,97,0,246,0,91,0,50,0,0,0,38,0,1,0,158,0,90,0,6,0,0,0,39,0,254,0,108,0,0,0,54,0,250,0,231,0,156,0,201,0,27,0,15,0,0,0,53,0,133,0,217,0,46,0,0,0,0,0,0,0,140,0,187,0,53,0,102,0,0,0,214,0,99,0,225,0,39,0,65,0,79,0,63,0,72,0,100,0,18,0,200,0,0,0,248,0,143,0,53,0,247,0,248,0,57,0,73,0,57,0,188,0,0,0,248,0,172,0,0,0,7,0,89,0,241,0,0,0,104,0,60,0,12,0,92,0,0,0,191,0,126,0,143,0,0,0,205,0,92,0,0,0,0,0,218,0,192,0,149,0,83,0,0,0,215,0,0,0,154,0,0,0,141,0,0,0,0,0,44,0,2,0,114,0,213,0,79,0,68,0,102,0,154,0,171,0,160,0,71,0,29,0,44,0,129,0,41,0,187,0,151,0,0,0,105,0,104,0,175,0,14,0,0,0,0,0,0,0,207,0,0,0,0,0,189,0,92,0,245,0,246,0,35,0,197,0,118,0,177,0,120,0,249,0,0,0,151,0,149,0,28,0,74,0,81,0,105,0,33,0,167,0,0,0,12,0,198,0,38,0,132,0,204,0,53,0,138,0,170,0,0,0,0,0,0,0,0,0,130,0,109,0,0,0,169,0,187,0,0,0,19,0,102,0,40,0,0,0,162,0,167,0,205,0,114,0,43,0,55,0,239,0,0,0,11,0,86,0,0,0,168,0,2,0,184,0,115,0,238,0,0,0,69,0,74,0,46,0,0,0,68,0,46,0,0,0,143,0,150,0,69,0,82,0,0,0,0,0,62,0,26,0,147,0,62,0,0,0,87,0,78,0,141,0,0,0,50,0,22,0,35,0,42,0,213,0,123,0,81,0,176,0,48,0,195,0,67,0,177,0,75,0,128,0,81,0,241,0,0,0,202,0,185,0,253,0,212,0,239,0,0,0,175,0,67,0,186,0,25,0,219,0,240,0,129,0,0,0);
signal scenario_full  : scenario_type := (96,31,96,30,247,31,247,30,247,29,247,28,189,31,228,31,122,31,122,30,96,31,199,31,101,31,124,31,90,31,185,31,185,30,9,31,188,31,188,30,124,31,110,31,44,31,23,31,209,31,64,31,183,31,112,31,244,31,244,30,244,29,79,31,112,31,188,31,106,31,131,31,62,31,62,30,112,31,112,30,184,31,179,31,62,31,199,31,151,31,122,31,102,31,63,31,28,31,210,31,241,31,198,31,240,31,188,31,158,31,143,31,143,30,244,31,55,31,226,31,226,30,132,31,131,31,131,30,173,31,240,31,60,31,141,31,218,31,218,30,140,31,80,31,179,31,72,31,48,31,62,31,22,31,178,31,204,31,73,31,121,31,121,30,121,29,26,31,255,31,118,31,118,30,118,29,17,31,17,30,6,31,82,31,21,31,186,31,186,30,21,31,1,31,233,31,233,30,233,29,64,31,237,31,183,31,163,31,93,31,55,31,194,31,27,31,27,30,124,31,124,30,124,29,124,28,2,31,19,31,252,31,252,30,50,31,106,31,178,31,228,31,81,31,98,31,124,31,2,31,127,31,246,31,223,31,253,31,242,31,133,31,133,30,98,31,32,31,75,31,86,31,86,30,86,29,197,31,197,30,236,31,101,31,27,31,78,31,196,31,149,31,49,31,248,31,229,31,155,31,210,31,171,31,221,31,147,31,11,31,124,31,225,31,186,31,186,30,61,31,49,31,49,30,116,31,169,31,170,31,195,31,93,31,119,31,237,31,237,30,163,31,102,31,170,31,226,31,73,31,73,30,28,31,76,31,76,30,4,31,77,31,77,30,208,31,193,31,59,31,192,31,23,31,178,31,77,31,246,31,97,31,97,30,239,31,27,31,180,31,238,31,122,31,227,31,236,31,171,31,1,31,243,31,243,30,130,31,130,30,147,31,24,31,26,31,19,31,133,31,45,31,133,31,2,31,160,31,160,30,188,31,222,31,83,31,83,30,83,29,181,31,152,31,107,31,66,31,129,31,34,31,202,31,61,31,166,31,195,31,43,31,98,31,53,31,86,31,49,31,238,31,103,31,164,31,32,31,185,31,81,31,243,31,243,30,95,31,55,31,59,31,59,30,20,31,176,31,109,31,250,31,128,31,179,31,168,31,199,31,224,31,203,31,244,31,190,31,88,31,88,30,54,31,3,31,41,31,30,31,220,31,197,31,73,31,246,31,246,30,239,31,35,31,93,31,202,31,202,30,17,31,219,31,109,31,226,31,226,30,193,31,61,31,193,31,5,31,200,31,116,31,176,31,146,31,36,31,36,30,127,31,127,30,57,31,57,30,48,31,82,31,82,30,136,31,193,31,13,31,252,31,76,31,76,30,3,31,48,31,236,31,201,31,129,31,125,31,39,31,84,31,180,31,180,30,171,31,137,31,40,31,198,31,41,31,143,31,77,31,88,31,184,31,243,31,243,30,252,31,236,31,236,30,236,29,202,31,48,31,161,31,161,30,142,31,57,31,221,31,190,31,89,31,191,31,214,31,214,30,211,31,35,31,197,31,254,31,254,30,14,31,85,31,197,31,91,31,181,31,236,31,114,31,78,31,147,31,136,31,225,31,225,30,225,29,23,31,67,31,17,31,138,31,138,30,2,31,65,31,222,31,44,31,44,30,67,31,209,31,26,31,157,31,194,31,187,31,230,31,169,31,169,30,11,31,165,31,165,30,216,31,148,31,29,31,19,31,102,31,32,31,55,31,38,31,34,31,194,31,228,31,49,31,149,31,206,31,70,31,8,31,97,31,246,31,91,31,50,31,50,30,38,31,1,31,158,31,90,31,6,31,6,30,39,31,254,31,108,31,108,30,54,31,250,31,231,31,156,31,201,31,27,31,15,31,15,30,53,31,133,31,217,31,46,31,46,30,46,29,46,28,140,31,187,31,53,31,102,31,102,30,214,31,99,31,225,31,39,31,65,31,79,31,63,31,72,31,100,31,18,31,200,31,200,30,248,31,143,31,53,31,247,31,248,31,57,31,73,31,57,31,188,31,188,30,248,31,172,31,172,30,7,31,89,31,241,31,241,30,104,31,60,31,12,31,92,31,92,30,191,31,126,31,143,31,143,30,205,31,92,31,92,30,92,29,218,31,192,31,149,31,83,31,83,30,215,31,215,30,154,31,154,30,141,31,141,30,141,29,44,31,2,31,114,31,213,31,79,31,68,31,102,31,154,31,171,31,160,31,71,31,29,31,44,31,129,31,41,31,187,31,151,31,151,30,105,31,104,31,175,31,14,31,14,30,14,29,14,28,207,31,207,30,207,29,189,31,92,31,245,31,246,31,35,31,197,31,118,31,177,31,120,31,249,31,249,30,151,31,149,31,28,31,74,31,81,31,105,31,33,31,167,31,167,30,12,31,198,31,38,31,132,31,204,31,53,31,138,31,170,31,170,30,170,29,170,28,170,27,130,31,109,31,109,30,169,31,187,31,187,30,19,31,102,31,40,31,40,30,162,31,167,31,205,31,114,31,43,31,55,31,239,31,239,30,11,31,86,31,86,30,168,31,2,31,184,31,115,31,238,31,238,30,69,31,74,31,46,31,46,30,68,31,46,31,46,30,143,31,150,31,69,31,82,31,82,30,82,29,62,31,26,31,147,31,62,31,62,30,87,31,78,31,141,31,141,30,50,31,22,31,35,31,42,31,213,31,123,31,81,31,176,31,48,31,195,31,67,31,177,31,75,31,128,31,81,31,241,31,241,30,202,31,185,31,253,31,212,31,239,31,239,30,175,31,67,31,186,31,25,31,219,31,240,31,129,31,129,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
