-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 356;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (64,0,116,0,232,0,0,0,0,0,73,0,74,0,189,0,99,0,113,0,0,0,16,0,80,0,113,0,84,0,0,0,109,0,145,0,167,0,54,0,227,0,19,0,165,0,0,0,169,0,108,0,176,0,135,0,189,0,0,0,0,0,1,0,24,0,154,0,0,0,77,0,150,0,0,0,233,0,90,0,80,0,0,0,57,0,244,0,0,0,17,0,155,0,186,0,245,0,102,0,51,0,215,0,58,0,235,0,169,0,107,0,226,0,218,0,224,0,230,0,0,0,37,0,240,0,39,0,103,0,171,0,87,0,3,0,55,0,241,0,239,0,157,0,36,0,45,0,242,0,119,0,75,0,24,0,111,0,86,0,0,0,35,0,102,0,103,0,0,0,61,0,83,0,120,0,243,0,54,0,15,0,0,0,132,0,82,0,0,0,143,0,210,0,161,0,125,0,228,0,0,0,63,0,213,0,215,0,64,0,138,0,238,0,185,0,0,0,142,0,122,0,0,0,72,0,97,0,183,0,134,0,144,0,64,0,94,0,245,0,0,0,207,0,0,0,100,0,31,0,189,0,80,0,0,0,120,0,37,0,17,0,27,0,11,0,61,0,11,0,0,0,194,0,78,0,96,0,0,0,148,0,0,0,143,0,87,0,179,0,79,0,244,0,50,0,127,0,0,0,29,0,89,0,175,0,94,0,194,0,84,0,245,0,82,0,243,0,0,0,211,0,141,0,0,0,210,0,102,0,101,0,34,0,165,0,55,0,134,0,0,0,111,0,0,0,91,0,106,0,126,0,0,0,157,0,124,0,224,0,0,0,12,0,217,0,0,0,46,0,0,0,88,0,30,0,0,0,0,0,128,0,0,0,175,0,67,0,0,0,190,0,98,0,205,0,34,0,0,0,79,0,21,0,0,0,249,0,225,0,90,0,107,0,13,0,214,0,163,0,0,0,25,0,22,0,97,0,215,0,0,0,10,0,140,0,130,0,0,0,239,0,23,0,94,0,148,0,91,0,44,0,163,0,6,0,60,0,209,0,0,0,34,0,131,0,86,0,58,0,37,0,244,0,53,0,227,0,107,0,110,0,151,0,43,0,177,0,201,0,172,0,224,0,0,0,26,0,16,0,138,0,101,0,48,0,11,0,158,0,0,0,209,0,0,0,164,0,163,0,91,0,200,0,207,0,16,0,226,0,2,0,93,0,170,0,0,0,251,0,196,0,60,0,132,0,22,0,0,0,0,0,244,0,238,0,87,0,0,0,116,0,198,0,249,0,36,0,83,0,222,0,27,0,110,0,207,0,40,0,139,0,0,0,12,0,83,0,194,0,160,0,255,0,0,0,183,0,235,0,139,0,155,0,160,0,46,0,0,0,24,0,43,0,111,0,15,0,76,0,64,0,183,0,221,0,78,0,35,0,96,0,38,0,181,0,184,0,223,0,0,0,237,0,7,0,4,0,123,0,80,0,64,0,0,0,104,0,231,0,0,0,0,0,0,0,202,0,161,0,249,0,146,0,57,0,121,0,244,0,122,0,144,0,131,0,252,0,0,0,121,0,46,0,183,0,0,0,177,0,0,0,77,0,168,0,240,0,230,0,213,0);
signal scenario_full  : scenario_type := (64,31,116,31,232,31,232,30,232,29,73,31,74,31,189,31,99,31,113,31,113,30,16,31,80,31,113,31,84,31,84,30,109,31,145,31,167,31,54,31,227,31,19,31,165,31,165,30,169,31,108,31,176,31,135,31,189,31,189,30,189,29,1,31,24,31,154,31,154,30,77,31,150,31,150,30,233,31,90,31,80,31,80,30,57,31,244,31,244,30,17,31,155,31,186,31,245,31,102,31,51,31,215,31,58,31,235,31,169,31,107,31,226,31,218,31,224,31,230,31,230,30,37,31,240,31,39,31,103,31,171,31,87,31,3,31,55,31,241,31,239,31,157,31,36,31,45,31,242,31,119,31,75,31,24,31,111,31,86,31,86,30,35,31,102,31,103,31,103,30,61,31,83,31,120,31,243,31,54,31,15,31,15,30,132,31,82,31,82,30,143,31,210,31,161,31,125,31,228,31,228,30,63,31,213,31,215,31,64,31,138,31,238,31,185,31,185,30,142,31,122,31,122,30,72,31,97,31,183,31,134,31,144,31,64,31,94,31,245,31,245,30,207,31,207,30,100,31,31,31,189,31,80,31,80,30,120,31,37,31,17,31,27,31,11,31,61,31,11,31,11,30,194,31,78,31,96,31,96,30,148,31,148,30,143,31,87,31,179,31,79,31,244,31,50,31,127,31,127,30,29,31,89,31,175,31,94,31,194,31,84,31,245,31,82,31,243,31,243,30,211,31,141,31,141,30,210,31,102,31,101,31,34,31,165,31,55,31,134,31,134,30,111,31,111,30,91,31,106,31,126,31,126,30,157,31,124,31,224,31,224,30,12,31,217,31,217,30,46,31,46,30,88,31,30,31,30,30,30,29,128,31,128,30,175,31,67,31,67,30,190,31,98,31,205,31,34,31,34,30,79,31,21,31,21,30,249,31,225,31,90,31,107,31,13,31,214,31,163,31,163,30,25,31,22,31,97,31,215,31,215,30,10,31,140,31,130,31,130,30,239,31,23,31,94,31,148,31,91,31,44,31,163,31,6,31,60,31,209,31,209,30,34,31,131,31,86,31,58,31,37,31,244,31,53,31,227,31,107,31,110,31,151,31,43,31,177,31,201,31,172,31,224,31,224,30,26,31,16,31,138,31,101,31,48,31,11,31,158,31,158,30,209,31,209,30,164,31,163,31,91,31,200,31,207,31,16,31,226,31,2,31,93,31,170,31,170,30,251,31,196,31,60,31,132,31,22,31,22,30,22,29,244,31,238,31,87,31,87,30,116,31,198,31,249,31,36,31,83,31,222,31,27,31,110,31,207,31,40,31,139,31,139,30,12,31,83,31,194,31,160,31,255,31,255,30,183,31,235,31,139,31,155,31,160,31,46,31,46,30,24,31,43,31,111,31,15,31,76,31,64,31,183,31,221,31,78,31,35,31,96,31,38,31,181,31,184,31,223,31,223,30,237,31,7,31,4,31,123,31,80,31,64,31,64,30,104,31,231,31,231,30,231,29,231,28,202,31,161,31,249,31,146,31,57,31,121,31,244,31,122,31,144,31,131,31,252,31,252,30,121,31,46,31,183,31,183,30,177,31,177,30,77,31,168,31,240,31,230,31,213,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
