-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 688;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,123,0,60,0,185,0,12,0,29,0,244,0,53,0,95,0,77,0,163,0,244,0,48,0,0,0,237,0,167,0,224,0,65,0,164,0,38,0,110,0,45,0,0,0,142,0,163,0,20,0,79,0,173,0,91,0,55,0,34,0,218,0,122,0,127,0,65,0,127,0,102,0,209,0,50,0,38,0,1,0,0,0,205,0,116,0,172,0,114,0,140,0,200,0,74,0,192,0,228,0,0,0,210,0,4,0,123,0,78,0,0,0,206,0,0,0,116,0,25,0,96,0,110,0,202,0,199,0,0,0,59,0,114,0,160,0,29,0,211,0,180,0,64,0,76,0,236,0,199,0,0,0,3,0,64,0,53,0,109,0,141,0,238,0,0,0,0,0,9,0,41,0,196,0,208,0,17,0,69,0,0,0,0,0,227,0,0,0,0,0,183,0,30,0,134,0,92,0,131,0,2,0,132,0,147,0,151,0,209,0,124,0,0,0,0,0,0,0,81,0,222,0,44,0,157,0,189,0,0,0,213,0,0,0,63,0,192,0,238,0,204,0,108,0,111,0,0,0,233,0,191,0,0,0,159,0,21,0,33,0,121,0,222,0,17,0,242,0,179,0,44,0,0,0,124,0,29,0,101,0,0,0,234,0,54,0,148,0,62,0,49,0,201,0,90,0,114,0,135,0,53,0,177,0,50,0,170,0,204,0,144,0,198,0,20,0,108,0,5,0,222,0,108,0,175,0,240,0,229,0,144,0,100,0,0,0,107,0,0,0,125,0,91,0,48,0,122,0,105,0,237,0,207,0,116,0,210,0,59,0,117,0,0,0,62,0,0,0,84,0,191,0,47,0,86,0,218,0,181,0,125,0,0,0,192,0,14,0,157,0,116,0,59,0,36,0,131,0,68,0,249,0,0,0,0,0,20,0,0,0,77,0,170,0,126,0,157,0,0,0,134,0,210,0,133,0,0,0,224,0,78,0,252,0,0,0,13,0,140,0,0,0,113,0,208,0,6,0,98,0,0,0,0,0,162,0,7,0,118,0,0,0,245,0,0,0,154,0,0,0,0,0,32,0,18,0,22,0,230,0,129,0,106,0,65,0,0,0,15,0,0,0,207,0,159,0,34,0,0,0,72,0,60,0,0,0,125,0,189,0,100,0,27,0,114,0,80,0,206,0,55,0,212,0,245,0,150,0,0,0,187,0,39,0,85,0,59,0,210,0,170,0,12,0,200,0,79,0,139,0,206,0,34,0,81,0,57,0,220,0,0,0,78,0,209,0,38,0,97,0,97,0,0,0,0,0,44,0,0,0,185,0,0,0,197,0,139,0,242,0,102,0,23,0,150,0,0,0,74,0,47,0,241,0,57,0,43,0,5,0,111,0,56,0,174,0,59,0,251,0,196,0,193,0,41,0,95,0,17,0,151,0,81,0,44,0,0,0,23,0,234,0,99,0,233,0,111,0,0,0,84,0,93,0,104,0,0,0,0,0,0,0,148,0,55,0,13,0,148,0,236,0,167,0,72,0,37,0,40,0,22,0,159,0,224,0,0,0,63,0,36,0,200,0,121,0,162,0,120,0,131,0,5,0,0,0,186,0,165,0,0,0,148,0,0,0,9,0,0,0,174,0,150,0,76,0,50,0,15,0,218,0,0,0,226,0,250,0,59,0,205,0,192,0,63,0,200,0,15,0,133,0,33,0,218,0,71,0,12,0,131,0,240,0,167,0,59,0,3,0,86,0,0,0,0,0,162,0,0,0,209,0,241,0,100,0,50,0,251,0,17,0,23,0,168,0,235,0,78,0,67,0,157,0,0,0,1,0,93,0,110,0,0,0,129,0,137,0,236,0,168,0,0,0,218,0,101,0,0,0,51,0,253,0,125,0,161,0,222,0,0,0,147,0,131,0,39,0,29,0,163,0,0,0,207,0,159,0,243,0,138,0,188,0,178,0,222,0,0,0,58,0,29,0,104,0,171,0,118,0,144,0,233,0,138,0,151,0,127,0,0,0,0,0,0,0,12,0,209,0,26,0,175,0,60,0,213,0,1,0,90,0,210,0,77,0,0,0,0,0,6,0,240,0,252,0,235,0,0,0,130,0,100,0,111,0,1,0,217,0,249,0,224,0,0,0,235,0,93,0,61,0,42,0,0,0,0,0,6,0,0,0,125,0,0,0,150,0,0,0,180,0,0,0,194,0,161,0,233,0,237,0,0,0,112,0,18,0,0,0,154,0,145,0,72,0,0,0,0,0,83,0,121,0,248,0,212,0,0,0,79,0,249,0,72,0,131,0,107,0,17,0,218,0,112,0,183,0,0,0,0,0,0,0,46,0,166,0,148,0,169,0,213,0,250,0,121,0,19,0,247,0,71,0,0,0,224,0,0,0,214,0,239,0,50,0,233,0,169,0,201,0,0,0,53,0,170,0,204,0,0,0,0,0,197,0,146,0,136,0,227,0,98,0,168,0,96,0,16,0,112,0,203,0,4,0,137,0,42,0,167,0,246,0,77,0,0,0,46,0,249,0,50,0,119,0,0,0,0,0,206,0,19,0,212,0,204,0,150,0,211,0,238,0,0,0,252,0,166,0,252,0,12,0,151,0,23,0,249,0,227,0,210,0,219,0,39,0,42,0,0,0,14,0,0,0,11,0,15,0,6,0,189,0,194,0,0,0,57,0,0,0,0,0,48,0,95,0,169,0,243,0,71,0,45,0,95,0,0,0,0,0,165,0,12,0,209,0,229,0,128,0,12,0,76,0,180,0,180,0,0,0,45,0,0,0,118,0,162,0,140,0,109,0,161,0,131,0,20,0,37,0,89,0,194,0,9,0,0,0,0,0,153,0,237,0,0,0,0,0,155,0,0,0,203,0,167,0,192,0,234,0,216,0,122,0,55,0,0,0,0,0,7,0,0,0,122,0,46,0,0,0,39,0,137,0,41,0,214,0,248,0,220,0,0,0,52,0,89,0,15,0,0,0,188,0,198,0,44,0,0,0,182,0,147,0,73,0,246,0,94,0,0,0,150,0,82,0,242,0,115,0,22,0,53,0,81,0,142,0,113,0,200,0,44,0,194,0,174,0,0,0,0,0);
signal scenario_full  : scenario_type := (0,0,123,31,60,31,185,31,12,31,29,31,244,31,53,31,95,31,77,31,163,31,244,31,48,31,48,30,237,31,167,31,224,31,65,31,164,31,38,31,110,31,45,31,45,30,142,31,163,31,20,31,79,31,173,31,91,31,55,31,34,31,218,31,122,31,127,31,65,31,127,31,102,31,209,31,50,31,38,31,1,31,1,30,205,31,116,31,172,31,114,31,140,31,200,31,74,31,192,31,228,31,228,30,210,31,4,31,123,31,78,31,78,30,206,31,206,30,116,31,25,31,96,31,110,31,202,31,199,31,199,30,59,31,114,31,160,31,29,31,211,31,180,31,64,31,76,31,236,31,199,31,199,30,3,31,64,31,53,31,109,31,141,31,238,31,238,30,238,29,9,31,41,31,196,31,208,31,17,31,69,31,69,30,69,29,227,31,227,30,227,29,183,31,30,31,134,31,92,31,131,31,2,31,132,31,147,31,151,31,209,31,124,31,124,30,124,29,124,28,81,31,222,31,44,31,157,31,189,31,189,30,213,31,213,30,63,31,192,31,238,31,204,31,108,31,111,31,111,30,233,31,191,31,191,30,159,31,21,31,33,31,121,31,222,31,17,31,242,31,179,31,44,31,44,30,124,31,29,31,101,31,101,30,234,31,54,31,148,31,62,31,49,31,201,31,90,31,114,31,135,31,53,31,177,31,50,31,170,31,204,31,144,31,198,31,20,31,108,31,5,31,222,31,108,31,175,31,240,31,229,31,144,31,100,31,100,30,107,31,107,30,125,31,91,31,48,31,122,31,105,31,237,31,207,31,116,31,210,31,59,31,117,31,117,30,62,31,62,30,84,31,191,31,47,31,86,31,218,31,181,31,125,31,125,30,192,31,14,31,157,31,116,31,59,31,36,31,131,31,68,31,249,31,249,30,249,29,20,31,20,30,77,31,170,31,126,31,157,31,157,30,134,31,210,31,133,31,133,30,224,31,78,31,252,31,252,30,13,31,140,31,140,30,113,31,208,31,6,31,98,31,98,30,98,29,162,31,7,31,118,31,118,30,245,31,245,30,154,31,154,30,154,29,32,31,18,31,22,31,230,31,129,31,106,31,65,31,65,30,15,31,15,30,207,31,159,31,34,31,34,30,72,31,60,31,60,30,125,31,189,31,100,31,27,31,114,31,80,31,206,31,55,31,212,31,245,31,150,31,150,30,187,31,39,31,85,31,59,31,210,31,170,31,12,31,200,31,79,31,139,31,206,31,34,31,81,31,57,31,220,31,220,30,78,31,209,31,38,31,97,31,97,31,97,30,97,29,44,31,44,30,185,31,185,30,197,31,139,31,242,31,102,31,23,31,150,31,150,30,74,31,47,31,241,31,57,31,43,31,5,31,111,31,56,31,174,31,59,31,251,31,196,31,193,31,41,31,95,31,17,31,151,31,81,31,44,31,44,30,23,31,234,31,99,31,233,31,111,31,111,30,84,31,93,31,104,31,104,30,104,29,104,28,148,31,55,31,13,31,148,31,236,31,167,31,72,31,37,31,40,31,22,31,159,31,224,31,224,30,63,31,36,31,200,31,121,31,162,31,120,31,131,31,5,31,5,30,186,31,165,31,165,30,148,31,148,30,9,31,9,30,174,31,150,31,76,31,50,31,15,31,218,31,218,30,226,31,250,31,59,31,205,31,192,31,63,31,200,31,15,31,133,31,33,31,218,31,71,31,12,31,131,31,240,31,167,31,59,31,3,31,86,31,86,30,86,29,162,31,162,30,209,31,241,31,100,31,50,31,251,31,17,31,23,31,168,31,235,31,78,31,67,31,157,31,157,30,1,31,93,31,110,31,110,30,129,31,137,31,236,31,168,31,168,30,218,31,101,31,101,30,51,31,253,31,125,31,161,31,222,31,222,30,147,31,131,31,39,31,29,31,163,31,163,30,207,31,159,31,243,31,138,31,188,31,178,31,222,31,222,30,58,31,29,31,104,31,171,31,118,31,144,31,233,31,138,31,151,31,127,31,127,30,127,29,127,28,12,31,209,31,26,31,175,31,60,31,213,31,1,31,90,31,210,31,77,31,77,30,77,29,6,31,240,31,252,31,235,31,235,30,130,31,100,31,111,31,1,31,217,31,249,31,224,31,224,30,235,31,93,31,61,31,42,31,42,30,42,29,6,31,6,30,125,31,125,30,150,31,150,30,180,31,180,30,194,31,161,31,233,31,237,31,237,30,112,31,18,31,18,30,154,31,145,31,72,31,72,30,72,29,83,31,121,31,248,31,212,31,212,30,79,31,249,31,72,31,131,31,107,31,17,31,218,31,112,31,183,31,183,30,183,29,183,28,46,31,166,31,148,31,169,31,213,31,250,31,121,31,19,31,247,31,71,31,71,30,224,31,224,30,214,31,239,31,50,31,233,31,169,31,201,31,201,30,53,31,170,31,204,31,204,30,204,29,197,31,146,31,136,31,227,31,98,31,168,31,96,31,16,31,112,31,203,31,4,31,137,31,42,31,167,31,246,31,77,31,77,30,46,31,249,31,50,31,119,31,119,30,119,29,206,31,19,31,212,31,204,31,150,31,211,31,238,31,238,30,252,31,166,31,252,31,12,31,151,31,23,31,249,31,227,31,210,31,219,31,39,31,42,31,42,30,14,31,14,30,11,31,15,31,6,31,189,31,194,31,194,30,57,31,57,30,57,29,48,31,95,31,169,31,243,31,71,31,45,31,95,31,95,30,95,29,165,31,12,31,209,31,229,31,128,31,12,31,76,31,180,31,180,31,180,30,45,31,45,30,118,31,162,31,140,31,109,31,161,31,131,31,20,31,37,31,89,31,194,31,9,31,9,30,9,29,153,31,237,31,237,30,237,29,155,31,155,30,203,31,167,31,192,31,234,31,216,31,122,31,55,31,55,30,55,29,7,31,7,30,122,31,46,31,46,30,39,31,137,31,41,31,214,31,248,31,220,31,220,30,52,31,89,31,15,31,15,30,188,31,198,31,44,31,44,30,182,31,147,31,73,31,246,31,94,31,94,30,150,31,82,31,242,31,115,31,22,31,53,31,81,31,142,31,113,31,200,31,44,31,194,31,174,31,174,30,174,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
