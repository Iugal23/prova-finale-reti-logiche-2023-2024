-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 942;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,123,0,24,0,193,0,57,0,106,0,182,0,66,0,0,0,0,0,21,0,0,0,227,0,0,0,221,0,47,0,211,0,0,0,198,0,6,0,191,0,67,0,168,0,106,0,63,0,185,0,118,0,0,0,81,0,0,0,179,0,131,0,169,0,120,0,0,0,191,0,58,0,248,0,249,0,78,0,0,0,0,0,112,0,0,0,182,0,8,0,160,0,200,0,30,0,216,0,249,0,230,0,242,0,183,0,0,0,118,0,166,0,0,0,180,0,101,0,39,0,229,0,0,0,143,0,38,0,200,0,119,0,59,0,248,0,214,0,31,0,241,0,154,0,165,0,72,0,92,0,233,0,158,0,28,0,11,0,46,0,87,0,177,0,242,0,237,0,197,0,138,0,0,0,25,0,228,0,0,0,223,0,168,0,0,0,61,0,11,0,0,0,126,0,3,0,201,0,130,0,66,0,60,0,118,0,33,0,0,0,199,0,58,0,14,0,12,0,124,0,111,0,24,0,196,0,108,0,55,0,101,0,12,0,0,0,13,0,186,0,116,0,0,0,211,0,254,0,252,0,122,0,62,0,237,0,120,0,145,0,59,0,253,0,0,0,3,0,18,0,42,0,9,0,0,0,87,0,105,0,150,0,0,0,45,0,199,0,36,0,135,0,73,0,0,0,58,0,126,0,23,0,165,0,104,0,106,0,23,0,62,0,0,0,174,0,139,0,4,0,210,0,0,0,175,0,207,0,0,0,0,0,0,0,22,0,193,0,40,0,0,0,10,0,214,0,76,0,127,0,213,0,62,0,221,0,208,0,224,0,99,0,189,0,56,0,162,0,168,0,57,0,69,0,112,0,255,0,0,0,241,0,197,0,130,0,247,0,0,0,4,0,172,0,245,0,216,0,0,0,23,0,157,0,224,0,172,0,89,0,159,0,63,0,149,0,147,0,0,0,0,0,37,0,112,0,71,0,0,0,238,0,229,0,33,0,35,0,74,0,69,0,209,0,181,0,54,0,98,0,0,0,0,0,45,0,29,0,122,0,145,0,165,0,27,0,226,0,40,0,153,0,0,0,136,0,0,0,132,0,235,0,1,0,199,0,80,0,186,0,107,0,105,0,152,0,147,0,254,0,0,0,0,0,0,0,147,0,73,0,181,0,196,0,49,0,56,0,222,0,174,0,54,0,0,0,155,0,36,0,248,0,136,0,142,0,51,0,253,0,97,0,167,0,114,0,31,0,153,0,56,0,16,0,160,0,78,0,189,0,40,0,67,0,160,0,109,0,156,0,171,0,233,0,204,0,135,0,0,0,248,0,216,0,247,0,43,0,0,0,0,0,106,0,19,0,201,0,0,0,78,0,53,0,0,0,78,0,172,0,233,0,111,0,50,0,216,0,97,0,60,0,87,0,23,0,7,0,0,0,198,0,0,0,155,0,119,0,0,0,239,0,0,0,78,0,0,0,23,0,172,0,183,0,151,0,172,0,0,0,13,0,197,0,92,0,236,0,17,0,79,0,63,0,165,0,0,0,0,0,181,0,241,0,240,0,12,0,0,0,0,0,105,0,0,0,192,0,0,0,116,0,0,0,85,0,0,0,0,0,76,0,0,0,205,0,0,0,0,0,211,0,0,0,96,0,153,0,38,0,0,0,96,0,94,0,102,0,0,0,234,0,67,0,167,0,0,0,0,0,0,0,249,0,16,0,0,0,232,0,45,0,0,0,22,0,162,0,94,0,199,0,116,0,210,0,93,0,72,0,0,0,0,0,42,0,31,0,0,0,82,0,136,0,232,0,0,0,43,0,0,0,233,0,136,0,0,0,59,0,0,0,0,0,191,0,115,0,0,0,0,0,193,0,162,0,64,0,67,0,0,0,0,0,111,0,86,0,241,0,210,0,8,0,181,0,52,0,62,0,21,0,115,0,238,0,0,0,0,0,199,0,0,0,182,0,228,0,53,0,137,0,18,0,209,0,39,0,29,0,0,0,121,0,216,0,93,0,251,0,78,0,218,0,238,0,12,0,178,0,13,0,6,0,226,0,90,0,0,0,112,0,101,0,0,0,0,0,64,0,126,0,228,0,198,0,0,0,43,0,238,0,125,0,0,0,0,0,13,0,217,0,247,0,0,0,119,0,0,0,0,0,0,0,131,0,34,0,118,0,212,0,59,0,91,0,135,0,32,0,0,0,163,0,0,0,233,0,210,0,40,0,6,0,0,0,255,0,33,0,90,0,0,0,3,0,251,0,0,0,122,0,107,0,118,0,26,0,52,0,209,0,176,0,13,0,0,0,145,0,0,0,63,0,0,0,235,0,13,0,86,0,174,0,11,0,0,0,0,0,211,0,0,0,215,0,14,0,6,0,109,0,0,0,46,0,0,0,200,0,17,0,96,0,99,0,148,0,78,0,31,0,190,0,119,0,126,0,0,0,0,0,48,0,0,0,0,0,192,0,130,0,0,0,133,0,0,0,242,0,206,0,159,0,98,0,0,0,43,0,140,0,0,0,254,0,0,0,0,0,4,0,210,0,12,0,164,0,232,0,183,0,135,0,87,0,151,0,96,0,46,0,78,0,0,0,153,0,153,0,8,0,23,0,85,0,161,0,214,0,154,0,32,0,213,0,112,0,0,0,252,0,24,0,0,0,82,0,199,0,50,0,241,0,0,0,0,0,114,0,202,0,114,0,154,0,250,0,225,0,109,0,104,0,68,0,180,0,212,0,10,0,224,0,16,0,60,0,199,0,193,0,215,0,0,0,131,0,119,0,145,0,208,0,0,0,0,0,206,0,87,0,59,0,30,0,67,0,8,0,54,0,0,0,165,0,153,0,158,0,207,0,216,0,252,0,138,0,0,0,74,0,65,0,243,0,125,0,151,0,151,0,56,0,176,0,26,0,0,0,40,0,41,0,35,0,0,0,200,0,57,0,116,0,83,0,51,0,230,0,121,0,214,0,198,0,211,0,103,0,99,0,0,0,90,0,220,0,221,0,222,0,59,0,12,0,0,0,174,0,0,0,0,0,203,0,0,0,5,0,11,0,105,0,0,0,39,0,154,0,220,0,213,0,28,0,214,0,187,0,147,0,230,0,133,0,175,0,74,0,192,0,29,0,128,0,60,0,245,0,0,0,81,0,0,0,0,0,36,0,0,0,0,0,0,0,31,0,0,0,0,0,80,0,146,0,27,0,220,0,89,0,0,0,244,0,161,0,217,0,62,0,5,0,166,0,200,0,150,0,42,0,218,0,215,0,167,0,187,0,43,0,82,0,215,0,38,0,18,0,210,0,86,0,126,0,208,0,91,0,86,0,204,0,72,0,124,0,201,0,68,0,205,0,109,0,222,0,155,0,3,0,108,0,0,0,116,0,231,0,0,0,23,0,50,0,246,0,53,0,108,0,106,0,121,0,238,0,2,0,163,0,94,0,110,0,86,0,143,0,0,0,12,0,0,0,228,0,67,0,169,0,97,0,203,0,69,0,15,0,0,0,25,0,146,0,47,0,254,0,0,0,6,0,24,0,172,0,121,0,153,0,103,0,0,0,227,0,154,0,204,0,102,0,0,0,61,0,191,0,218,0,0,0,0,0,0,0,181,0,223,0,204,0,72,0,151,0,0,0,251,0,51,0,122,0,51,0,161,0,0,0,108,0,0,0,0,0,0,0,212,0,0,0,136,0,2,0,219,0,192,0,0,0,44,0,201,0,82,0,24,0,0,0,22,0,62,0,128,0,250,0,136,0,210,0,37,0,13,0,142,0,222,0,181,0,171,0,145,0,254,0,0,0,95,0,61,0,109,0,209,0,84,0,86,0,164,0,164,0,165,0,219,0,0,0,0,0,28,0,233,0,235,0,49,0,48,0,118,0,150,0,69,0,93,0,0,0,112,0,74,0,127,0,99,0,239,0,0,0,127,0,0,0,94,0,0,0,9,0,129,0,25,0,125,0,167,0,115,0,190,0,0,0,0,0,93,0,0,0,43,0,0,0,1,0,54,0,153,0,41,0,0,0,215,0,0,0,242,0,246,0,75,0,52,0,0,0,22,0,83,0,67,0,97,0,175,0,0,0,132,0,20,0,96,0,152,0,89,0,235,0,175,0,181,0,104,0,207,0,93,0,212,0,154,0,242,0,72,0,10,0,0,0,0,0,222,0,87,0,140,0,153,0,0,0,126,0,47,0,127,0,0,0,1,0,0,0,16,0,0,0,46,0,216,0,0,0,50,0,0,0);
signal scenario_full  : scenario_type := (0,0,123,31,24,31,193,31,57,31,106,31,182,31,66,31,66,30,66,29,21,31,21,30,227,31,227,30,221,31,47,31,211,31,211,30,198,31,6,31,191,31,67,31,168,31,106,31,63,31,185,31,118,31,118,30,81,31,81,30,179,31,131,31,169,31,120,31,120,30,191,31,58,31,248,31,249,31,78,31,78,30,78,29,112,31,112,30,182,31,8,31,160,31,200,31,30,31,216,31,249,31,230,31,242,31,183,31,183,30,118,31,166,31,166,30,180,31,101,31,39,31,229,31,229,30,143,31,38,31,200,31,119,31,59,31,248,31,214,31,31,31,241,31,154,31,165,31,72,31,92,31,233,31,158,31,28,31,11,31,46,31,87,31,177,31,242,31,237,31,197,31,138,31,138,30,25,31,228,31,228,30,223,31,168,31,168,30,61,31,11,31,11,30,126,31,3,31,201,31,130,31,66,31,60,31,118,31,33,31,33,30,199,31,58,31,14,31,12,31,124,31,111,31,24,31,196,31,108,31,55,31,101,31,12,31,12,30,13,31,186,31,116,31,116,30,211,31,254,31,252,31,122,31,62,31,237,31,120,31,145,31,59,31,253,31,253,30,3,31,18,31,42,31,9,31,9,30,87,31,105,31,150,31,150,30,45,31,199,31,36,31,135,31,73,31,73,30,58,31,126,31,23,31,165,31,104,31,106,31,23,31,62,31,62,30,174,31,139,31,4,31,210,31,210,30,175,31,207,31,207,30,207,29,207,28,22,31,193,31,40,31,40,30,10,31,214,31,76,31,127,31,213,31,62,31,221,31,208,31,224,31,99,31,189,31,56,31,162,31,168,31,57,31,69,31,112,31,255,31,255,30,241,31,197,31,130,31,247,31,247,30,4,31,172,31,245,31,216,31,216,30,23,31,157,31,224,31,172,31,89,31,159,31,63,31,149,31,147,31,147,30,147,29,37,31,112,31,71,31,71,30,238,31,229,31,33,31,35,31,74,31,69,31,209,31,181,31,54,31,98,31,98,30,98,29,45,31,29,31,122,31,145,31,165,31,27,31,226,31,40,31,153,31,153,30,136,31,136,30,132,31,235,31,1,31,199,31,80,31,186,31,107,31,105,31,152,31,147,31,254,31,254,30,254,29,254,28,147,31,73,31,181,31,196,31,49,31,56,31,222,31,174,31,54,31,54,30,155,31,36,31,248,31,136,31,142,31,51,31,253,31,97,31,167,31,114,31,31,31,153,31,56,31,16,31,160,31,78,31,189,31,40,31,67,31,160,31,109,31,156,31,171,31,233,31,204,31,135,31,135,30,248,31,216,31,247,31,43,31,43,30,43,29,106,31,19,31,201,31,201,30,78,31,53,31,53,30,78,31,172,31,233,31,111,31,50,31,216,31,97,31,60,31,87,31,23,31,7,31,7,30,198,31,198,30,155,31,119,31,119,30,239,31,239,30,78,31,78,30,23,31,172,31,183,31,151,31,172,31,172,30,13,31,197,31,92,31,236,31,17,31,79,31,63,31,165,31,165,30,165,29,181,31,241,31,240,31,12,31,12,30,12,29,105,31,105,30,192,31,192,30,116,31,116,30,85,31,85,30,85,29,76,31,76,30,205,31,205,30,205,29,211,31,211,30,96,31,153,31,38,31,38,30,96,31,94,31,102,31,102,30,234,31,67,31,167,31,167,30,167,29,167,28,249,31,16,31,16,30,232,31,45,31,45,30,22,31,162,31,94,31,199,31,116,31,210,31,93,31,72,31,72,30,72,29,42,31,31,31,31,30,82,31,136,31,232,31,232,30,43,31,43,30,233,31,136,31,136,30,59,31,59,30,59,29,191,31,115,31,115,30,115,29,193,31,162,31,64,31,67,31,67,30,67,29,111,31,86,31,241,31,210,31,8,31,181,31,52,31,62,31,21,31,115,31,238,31,238,30,238,29,199,31,199,30,182,31,228,31,53,31,137,31,18,31,209,31,39,31,29,31,29,30,121,31,216,31,93,31,251,31,78,31,218,31,238,31,12,31,178,31,13,31,6,31,226,31,90,31,90,30,112,31,101,31,101,30,101,29,64,31,126,31,228,31,198,31,198,30,43,31,238,31,125,31,125,30,125,29,13,31,217,31,247,31,247,30,119,31,119,30,119,29,119,28,131,31,34,31,118,31,212,31,59,31,91,31,135,31,32,31,32,30,163,31,163,30,233,31,210,31,40,31,6,31,6,30,255,31,33,31,90,31,90,30,3,31,251,31,251,30,122,31,107,31,118,31,26,31,52,31,209,31,176,31,13,31,13,30,145,31,145,30,63,31,63,30,235,31,13,31,86,31,174,31,11,31,11,30,11,29,211,31,211,30,215,31,14,31,6,31,109,31,109,30,46,31,46,30,200,31,17,31,96,31,99,31,148,31,78,31,31,31,190,31,119,31,126,31,126,30,126,29,48,31,48,30,48,29,192,31,130,31,130,30,133,31,133,30,242,31,206,31,159,31,98,31,98,30,43,31,140,31,140,30,254,31,254,30,254,29,4,31,210,31,12,31,164,31,232,31,183,31,135,31,87,31,151,31,96,31,46,31,78,31,78,30,153,31,153,31,8,31,23,31,85,31,161,31,214,31,154,31,32,31,213,31,112,31,112,30,252,31,24,31,24,30,82,31,199,31,50,31,241,31,241,30,241,29,114,31,202,31,114,31,154,31,250,31,225,31,109,31,104,31,68,31,180,31,212,31,10,31,224,31,16,31,60,31,199,31,193,31,215,31,215,30,131,31,119,31,145,31,208,31,208,30,208,29,206,31,87,31,59,31,30,31,67,31,8,31,54,31,54,30,165,31,153,31,158,31,207,31,216,31,252,31,138,31,138,30,74,31,65,31,243,31,125,31,151,31,151,31,56,31,176,31,26,31,26,30,40,31,41,31,35,31,35,30,200,31,57,31,116,31,83,31,51,31,230,31,121,31,214,31,198,31,211,31,103,31,99,31,99,30,90,31,220,31,221,31,222,31,59,31,12,31,12,30,174,31,174,30,174,29,203,31,203,30,5,31,11,31,105,31,105,30,39,31,154,31,220,31,213,31,28,31,214,31,187,31,147,31,230,31,133,31,175,31,74,31,192,31,29,31,128,31,60,31,245,31,245,30,81,31,81,30,81,29,36,31,36,30,36,29,36,28,31,31,31,30,31,29,80,31,146,31,27,31,220,31,89,31,89,30,244,31,161,31,217,31,62,31,5,31,166,31,200,31,150,31,42,31,218,31,215,31,167,31,187,31,43,31,82,31,215,31,38,31,18,31,210,31,86,31,126,31,208,31,91,31,86,31,204,31,72,31,124,31,201,31,68,31,205,31,109,31,222,31,155,31,3,31,108,31,108,30,116,31,231,31,231,30,23,31,50,31,246,31,53,31,108,31,106,31,121,31,238,31,2,31,163,31,94,31,110,31,86,31,143,31,143,30,12,31,12,30,228,31,67,31,169,31,97,31,203,31,69,31,15,31,15,30,25,31,146,31,47,31,254,31,254,30,6,31,24,31,172,31,121,31,153,31,103,31,103,30,227,31,154,31,204,31,102,31,102,30,61,31,191,31,218,31,218,30,218,29,218,28,181,31,223,31,204,31,72,31,151,31,151,30,251,31,51,31,122,31,51,31,161,31,161,30,108,31,108,30,108,29,108,28,212,31,212,30,136,31,2,31,219,31,192,31,192,30,44,31,201,31,82,31,24,31,24,30,22,31,62,31,128,31,250,31,136,31,210,31,37,31,13,31,142,31,222,31,181,31,171,31,145,31,254,31,254,30,95,31,61,31,109,31,209,31,84,31,86,31,164,31,164,31,165,31,219,31,219,30,219,29,28,31,233,31,235,31,49,31,48,31,118,31,150,31,69,31,93,31,93,30,112,31,74,31,127,31,99,31,239,31,239,30,127,31,127,30,94,31,94,30,9,31,129,31,25,31,125,31,167,31,115,31,190,31,190,30,190,29,93,31,93,30,43,31,43,30,1,31,54,31,153,31,41,31,41,30,215,31,215,30,242,31,246,31,75,31,52,31,52,30,22,31,83,31,67,31,97,31,175,31,175,30,132,31,20,31,96,31,152,31,89,31,235,31,175,31,181,31,104,31,207,31,93,31,212,31,154,31,242,31,72,31,10,31,10,30,10,29,222,31,87,31,140,31,153,31,153,30,126,31,47,31,127,31,127,30,1,31,1,30,16,31,16,30,46,31,216,31,216,30,50,31,50,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
