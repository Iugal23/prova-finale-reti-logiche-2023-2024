-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 903;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (81,0,216,0,23,0,140,0,0,0,247,0,75,0,238,0,201,0,197,0,0,0,221,0,0,0,209,0,0,0,183,0,6,0,164,0,228,0,200,0,159,0,43,0,0,0,90,0,0,0,163,0,179,0,186,0,156,0,141,0,137,0,130,0,0,0,135,0,97,0,21,0,178,0,241,0,0,0,31,0,122,0,75,0,157,0,0,0,146,0,3,0,162,0,173,0,0,0,94,0,224,0,0,0,4,0,0,0,64,0,5,0,6,0,63,0,78,0,34,0,228,0,34,0,0,0,56,0,0,0,255,0,214,0,0,0,162,0,119,0,0,0,128,0,49,0,196,0,96,0,0,0,196,0,65,0,0,0,248,0,186,0,168,0,202,0,0,0,190,0,154,0,133,0,52,0,157,0,0,0,32,0,0,0,211,0,105,0,144,0,191,0,0,0,103,0,183,0,176,0,93,0,134,0,191,0,0,0,67,0,186,0,153,0,224,0,241,0,216,0,104,0,215,0,6,0,176,0,0,0,80,0,200,0,29,0,128,0,19,0,146,0,121,0,233,0,252,0,0,0,0,0,84,0,209,0,0,0,54,0,186,0,0,0,0,0,43,0,188,0,192,0,10,0,155,0,0,0,106,0,62,0,58,0,238,0,253,0,0,0,165,0,28,0,182,0,115,0,87,0,0,0,22,0,176,0,70,0,89,0,214,0,116,0,237,0,52,0,31,0,202,0,22,0,92,0,216,0,9,0,150,0,215,0,0,0,123,0,231,0,65,0,0,0,41,0,90,0,202,0,245,0,55,0,26,0,197,0,41,0,0,0,132,0,21,0,28,0,202,0,118,0,0,0,0,0,64,0,155,0,0,0,87,0,37,0,0,0,194,0,105,0,251,0,138,0,118,0,164,0,225,0,140,0,84,0,2,0,0,0,176,0,132,0,240,0,197,0,179,0,0,0,119,0,156,0,133,0,254,0,75,0,154,0,232,0,58,0,136,0,0,0,17,0,31,0,228,0,172,0,206,0,246,0,69,0,152,0,142,0,117,0,130,0,13,0,242,0,42,0,96,0,210,0,25,0,88,0,0,0,72,0,6,0,0,0,26,0,234,0,0,0,181,0,0,0,26,0,158,0,207,0,139,0,0,0,0,0,212,0,18,0,64,0,169,0,136,0,205,0,216,0,149,0,0,0,192,0,0,0,240,0,239,0,239,0,0,0,143,0,29,0,159,0,75,0,205,0,240,0,0,0,0,0,78,0,193,0,134,0,0,0,124,0,69,0,155,0,62,0,0,0,244,0,0,0,227,0,85,0,9,0,0,0,184,0,0,0,2,0,58,0,74,0,10,0,226,0,243,0,15,0,170,0,0,0,157,0,23,0,247,0,54,0,85,0,168,0,13,0,73,0,229,0,0,0,146,0,151,0,255,0,66,0,0,0,154,0,195,0,4,0,202,0,251,0,40,0,181,0,175,0,0,0,142,0,0,0,195,0,0,0,201,0,244,0,71,0,0,0,253,0,221,0,179,0,59,0,135,0,143,0,0,0,149,0,149,0,0,0,77,0,0,0,218,0,134,0,169,0,165,0,62,0,105,0,213,0,195,0,218,0,0,0,231,0,200,0,69,0,76,0,0,0,50,0,186,0,48,0,53,0,2,0,239,0,139,0,0,0,0,0,50,0,220,0,81,0,35,0,31,0,216,0,158,0,88,0,145,0,121,0,64,0,199,0,196,0,44,0,94,0,0,0,0,0,180,0,0,0,147,0,92,0,185,0,51,0,0,0,137,0,16,0,27,0,15,0,224,0,0,0,17,0,151,0,41,0,38,0,19,0,166,0,0,0,156,0,204,0,120,0,230,0,74,0,204,0,28,0,204,0,0,0,0,0,0,0,135,0,0,0,102,0,231,0,0,0,0,0,0,0,173,0,5,0,244,0,187,0,0,0,60,0,0,0,22,0,136,0,43,0,33,0,193,0,0,0,0,0,0,0,22,0,0,0,111,0,246,0,156,0,131,0,255,0,110,0,242,0,0,0,174,0,200,0,36,0,207,0,193,0,149,0,0,0,254,0,216,0,174,0,113,0,180,0,240,0,19,0,149,0,0,0,175,0,87,0,219,0,68,0,164,0,0,0,197,0,107,0,5,0,197,0,0,0,12,0,153,0,156,0,0,0,0,0,164,0,194,0,168,0,0,0,0,0,154,0,240,0,0,0,217,0,0,0,232,0,149,0,131,0,128,0,93,0,0,0,82,0,193,0,92,0,53,0,157,0,214,0,139,0,8,0,50,0,0,0,103,0,69,0,0,0,28,0,123,0,216,0,0,0,167,0,55,0,188,0,0,0,203,0,0,0,0,0,231,0,100,0,36,0,0,0,203,0,145,0,0,0,196,0,64,0,158,0,0,0,136,0,202,0,64,0,134,0,41,0,62,0,120,0,47,0,23,0,0,0,69,0,29,0,220,0,0,0,201,0,106,0,4,0,131,0,151,0,228,0,50,0,128,0,16,0,76,0,0,0,197,0,170,0,0,0,0,0,49,0,3,0,221,0,181,0,3,0,122,0,20,0,0,0,183,0,247,0,112,0,232,0,37,0,188,0,14,0,0,0,136,0,130,0,139,0,154,0,0,0,226,0,65,0,37,0,203,0,55,0,45,0,0,0,174,0,122,0,205,0,93,0,129,0,98,0,34,0,4,0,141,0,19,0,100,0,110,0,48,0,83,0,248,0,253,0,104,0,121,0,75,0,0,0,38,0,144,0,35,0,227,0,132,0,158,0,147,0,162,0,0,0,48,0,228,0,56,0,127,0,133,0,45,0,0,0,110,0,226,0,0,0,160,0,199,0,0,0,75,0,182,0,246,0,64,0,143,0,246,0,72,0,0,0,67,0,59,0,38,0,91,0,216,0,91,0,248,0,0,0,117,0,63,0,181,0,0,0,225,0,205,0,109,0,44,0,191,0,224,0,18,0,119,0,131,0,49,0,96,0,240,0,185,0,124,0,75,0,181,0,188,0,211,0,0,0,217,0,160,0,41,0,37,0,27,0,255,0,35,0,0,0,11,0,143,0,194,0,0,0,15,0,230,0,34,0,0,0,102,0,210,0,56,0,41,0,136,0,152,0,95,0,128,0,97,0,103,0,0,0,37,0,151,0,207,0,69,0,0,0,197,0,130,0,73,0,65,0,83,0,0,0,134,0,243,0,147,0,0,0,182,0,0,0,117,0,0,0,0,0,0,0,130,0,129,0,128,0,81,0,44,0,51,0,93,0,137,0,93,0,138,0,84,0,250,0,78,0,228,0,42,0,181,0,0,0,0,0,130,0,87,0,97,0,197,0,215,0,0,0,158,0,218,0,120,0,22,0,107,0,5,0,159,0,75,0,46,0,129,0,32,0,143,0,239,0,0,0,251,0,194,0,0,0,115,0,147,0,227,0,122,0,69,0,67,0,71,0,0,0,44,0,202,0,0,0,0,0,98,0,202,0,32,0,3,0,132,0,93,0,178,0,0,0,146,0,118,0,104,0,129,0,0,0,234,0,168,0,50,0,117,0,246,0,108,0,91,0,232,0,64,0,0,0,52,0,0,0,120,0,133,0,182,0,12,0,224,0,170,0,204,0,225,0,174,0,0,0,0,0,0,0,0,0,196,0,201,0,147,0,66,0,0,0,35,0,27,0,34,0,136,0,0,0,148,0,44,0,16,0,137,0,5,0,7,0,0,0,199,0,183,0,186,0,88,0,0,0,119,0,0,0,218,0,58,0,65,0,208,0,0,0,0,0,149,0,63,0,152,0,60,0,0,0,0,0,0,0,237,0,41,0,54,0,44,0,238,0,199,0,245,0,77,0,196,0,236,0,43,0,134,0,0,0,17,0,238,0,216,0,39,0,40,0,58,0,23,0,19,0,27,0,47,0,152,0,0,0,146,0,0,0,94,0,78,0,212,0,0,0,113,0,249,0,95,0,13,0,0,0,176,0,0,0,0,0,30,0,96,0,208,0,200,0,237,0,0,0,0,0,83,0,18,0,238,0,234,0,55,0,0,0,88,0,160,0,145,0);
signal scenario_full  : scenario_type := (81,31,216,31,23,31,140,31,140,30,247,31,75,31,238,31,201,31,197,31,197,30,221,31,221,30,209,31,209,30,183,31,6,31,164,31,228,31,200,31,159,31,43,31,43,30,90,31,90,30,163,31,179,31,186,31,156,31,141,31,137,31,130,31,130,30,135,31,97,31,21,31,178,31,241,31,241,30,31,31,122,31,75,31,157,31,157,30,146,31,3,31,162,31,173,31,173,30,94,31,224,31,224,30,4,31,4,30,64,31,5,31,6,31,63,31,78,31,34,31,228,31,34,31,34,30,56,31,56,30,255,31,214,31,214,30,162,31,119,31,119,30,128,31,49,31,196,31,96,31,96,30,196,31,65,31,65,30,248,31,186,31,168,31,202,31,202,30,190,31,154,31,133,31,52,31,157,31,157,30,32,31,32,30,211,31,105,31,144,31,191,31,191,30,103,31,183,31,176,31,93,31,134,31,191,31,191,30,67,31,186,31,153,31,224,31,241,31,216,31,104,31,215,31,6,31,176,31,176,30,80,31,200,31,29,31,128,31,19,31,146,31,121,31,233,31,252,31,252,30,252,29,84,31,209,31,209,30,54,31,186,31,186,30,186,29,43,31,188,31,192,31,10,31,155,31,155,30,106,31,62,31,58,31,238,31,253,31,253,30,165,31,28,31,182,31,115,31,87,31,87,30,22,31,176,31,70,31,89,31,214,31,116,31,237,31,52,31,31,31,202,31,22,31,92,31,216,31,9,31,150,31,215,31,215,30,123,31,231,31,65,31,65,30,41,31,90,31,202,31,245,31,55,31,26,31,197,31,41,31,41,30,132,31,21,31,28,31,202,31,118,31,118,30,118,29,64,31,155,31,155,30,87,31,37,31,37,30,194,31,105,31,251,31,138,31,118,31,164,31,225,31,140,31,84,31,2,31,2,30,176,31,132,31,240,31,197,31,179,31,179,30,119,31,156,31,133,31,254,31,75,31,154,31,232,31,58,31,136,31,136,30,17,31,31,31,228,31,172,31,206,31,246,31,69,31,152,31,142,31,117,31,130,31,13,31,242,31,42,31,96,31,210,31,25,31,88,31,88,30,72,31,6,31,6,30,26,31,234,31,234,30,181,31,181,30,26,31,158,31,207,31,139,31,139,30,139,29,212,31,18,31,64,31,169,31,136,31,205,31,216,31,149,31,149,30,192,31,192,30,240,31,239,31,239,31,239,30,143,31,29,31,159,31,75,31,205,31,240,31,240,30,240,29,78,31,193,31,134,31,134,30,124,31,69,31,155,31,62,31,62,30,244,31,244,30,227,31,85,31,9,31,9,30,184,31,184,30,2,31,58,31,74,31,10,31,226,31,243,31,15,31,170,31,170,30,157,31,23,31,247,31,54,31,85,31,168,31,13,31,73,31,229,31,229,30,146,31,151,31,255,31,66,31,66,30,154,31,195,31,4,31,202,31,251,31,40,31,181,31,175,31,175,30,142,31,142,30,195,31,195,30,201,31,244,31,71,31,71,30,253,31,221,31,179,31,59,31,135,31,143,31,143,30,149,31,149,31,149,30,77,31,77,30,218,31,134,31,169,31,165,31,62,31,105,31,213,31,195,31,218,31,218,30,231,31,200,31,69,31,76,31,76,30,50,31,186,31,48,31,53,31,2,31,239,31,139,31,139,30,139,29,50,31,220,31,81,31,35,31,31,31,216,31,158,31,88,31,145,31,121,31,64,31,199,31,196,31,44,31,94,31,94,30,94,29,180,31,180,30,147,31,92,31,185,31,51,31,51,30,137,31,16,31,27,31,15,31,224,31,224,30,17,31,151,31,41,31,38,31,19,31,166,31,166,30,156,31,204,31,120,31,230,31,74,31,204,31,28,31,204,31,204,30,204,29,204,28,135,31,135,30,102,31,231,31,231,30,231,29,231,28,173,31,5,31,244,31,187,31,187,30,60,31,60,30,22,31,136,31,43,31,33,31,193,31,193,30,193,29,193,28,22,31,22,30,111,31,246,31,156,31,131,31,255,31,110,31,242,31,242,30,174,31,200,31,36,31,207,31,193,31,149,31,149,30,254,31,216,31,174,31,113,31,180,31,240,31,19,31,149,31,149,30,175,31,87,31,219,31,68,31,164,31,164,30,197,31,107,31,5,31,197,31,197,30,12,31,153,31,156,31,156,30,156,29,164,31,194,31,168,31,168,30,168,29,154,31,240,31,240,30,217,31,217,30,232,31,149,31,131,31,128,31,93,31,93,30,82,31,193,31,92,31,53,31,157,31,214,31,139,31,8,31,50,31,50,30,103,31,69,31,69,30,28,31,123,31,216,31,216,30,167,31,55,31,188,31,188,30,203,31,203,30,203,29,231,31,100,31,36,31,36,30,203,31,145,31,145,30,196,31,64,31,158,31,158,30,136,31,202,31,64,31,134,31,41,31,62,31,120,31,47,31,23,31,23,30,69,31,29,31,220,31,220,30,201,31,106,31,4,31,131,31,151,31,228,31,50,31,128,31,16,31,76,31,76,30,197,31,170,31,170,30,170,29,49,31,3,31,221,31,181,31,3,31,122,31,20,31,20,30,183,31,247,31,112,31,232,31,37,31,188,31,14,31,14,30,136,31,130,31,139,31,154,31,154,30,226,31,65,31,37,31,203,31,55,31,45,31,45,30,174,31,122,31,205,31,93,31,129,31,98,31,34,31,4,31,141,31,19,31,100,31,110,31,48,31,83,31,248,31,253,31,104,31,121,31,75,31,75,30,38,31,144,31,35,31,227,31,132,31,158,31,147,31,162,31,162,30,48,31,228,31,56,31,127,31,133,31,45,31,45,30,110,31,226,31,226,30,160,31,199,31,199,30,75,31,182,31,246,31,64,31,143,31,246,31,72,31,72,30,67,31,59,31,38,31,91,31,216,31,91,31,248,31,248,30,117,31,63,31,181,31,181,30,225,31,205,31,109,31,44,31,191,31,224,31,18,31,119,31,131,31,49,31,96,31,240,31,185,31,124,31,75,31,181,31,188,31,211,31,211,30,217,31,160,31,41,31,37,31,27,31,255,31,35,31,35,30,11,31,143,31,194,31,194,30,15,31,230,31,34,31,34,30,102,31,210,31,56,31,41,31,136,31,152,31,95,31,128,31,97,31,103,31,103,30,37,31,151,31,207,31,69,31,69,30,197,31,130,31,73,31,65,31,83,31,83,30,134,31,243,31,147,31,147,30,182,31,182,30,117,31,117,30,117,29,117,28,130,31,129,31,128,31,81,31,44,31,51,31,93,31,137,31,93,31,138,31,84,31,250,31,78,31,228,31,42,31,181,31,181,30,181,29,130,31,87,31,97,31,197,31,215,31,215,30,158,31,218,31,120,31,22,31,107,31,5,31,159,31,75,31,46,31,129,31,32,31,143,31,239,31,239,30,251,31,194,31,194,30,115,31,147,31,227,31,122,31,69,31,67,31,71,31,71,30,44,31,202,31,202,30,202,29,98,31,202,31,32,31,3,31,132,31,93,31,178,31,178,30,146,31,118,31,104,31,129,31,129,30,234,31,168,31,50,31,117,31,246,31,108,31,91,31,232,31,64,31,64,30,52,31,52,30,120,31,133,31,182,31,12,31,224,31,170,31,204,31,225,31,174,31,174,30,174,29,174,28,174,27,196,31,201,31,147,31,66,31,66,30,35,31,27,31,34,31,136,31,136,30,148,31,44,31,16,31,137,31,5,31,7,31,7,30,199,31,183,31,186,31,88,31,88,30,119,31,119,30,218,31,58,31,65,31,208,31,208,30,208,29,149,31,63,31,152,31,60,31,60,30,60,29,60,28,237,31,41,31,54,31,44,31,238,31,199,31,245,31,77,31,196,31,236,31,43,31,134,31,134,30,17,31,238,31,216,31,39,31,40,31,58,31,23,31,19,31,27,31,47,31,152,31,152,30,146,31,146,30,94,31,78,31,212,31,212,30,113,31,249,31,95,31,13,31,13,30,176,31,176,30,176,29,30,31,96,31,208,31,200,31,237,31,237,30,237,29,83,31,18,31,238,31,234,31,55,31,55,30,88,31,160,31,145,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
