-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 750;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,139,0,105,0,0,0,174,0,36,0,240,0,227,0,21,0,127,0,67,0,168,0,146,0,172,0,0,0,0,0,194,0,158,0,0,0,187,0,75,0,44,0,118,0,121,0,140,0,79,0,10,0,0,0,39,0,155,0,204,0,173,0,235,0,0,0,131,0,194,0,30,0,0,0,41,0,101,0,213,0,71,0,91,0,181,0,0,0,0,0,178,0,85,0,236,0,62,0,152,0,94,0,80,0,0,0,0,0,155,0,218,0,238,0,178,0,184,0,0,0,55,0,18,0,0,0,46,0,255,0,120,0,0,0,0,0,141,0,201,0,66,0,57,0,14,0,221,0,182,0,0,0,58,0,14,0,0,0,235,0,83,0,0,0,122,0,0,0,15,0,24,0,25,0,202,0,9,0,0,0,0,0,59,0,96,0,149,0,22,0,0,0,184,0,135,0,136,0,0,0,0,0,235,0,39,0,220,0,46,0,149,0,0,0,243,0,188,0,129,0,0,0,0,0,8,0,34,0,213,0,60,0,112,0,146,0,0,0,0,0,199,0,27,0,0,0,89,0,181,0,109,0,99,0,164,0,253,0,229,0,176,0,69,0,135,0,224,0,69,0,0,0,241,0,0,0,151,0,0,0,0,0,0,0,4,0,13,0,238,0,161,0,70,0,229,0,98,0,0,0,202,0,242,0,207,0,79,0,53,0,0,0,11,0,251,0,0,0,145,0,36,0,198,0,250,0,169,0,112,0,0,0,12,0,244,0,110,0,56,0,217,0,155,0,81,0,118,0,115,0,0,0,135,0,57,0,0,0,157,0,0,0,150,0,235,0,137,0,219,0,0,0,80,0,227,0,0,0,229,0,142,0,213,0,72,0,36,0,0,0,38,0,56,0,229,0,0,0,92,0,196,0,51,0,59,0,170,0,220,0,228,0,184,0,14,0,122,0,23,0,97,0,188,0,254,0,168,0,22,0,197,0,170,0,144,0,0,0,19,0,232,0,0,0,19,0,0,0,0,0,148,0,52,0,162,0,123,0,0,0,0,0,0,0,119,0,170,0,0,0,240,0,0,0,75,0,246,0,114,0,25,0,63,0,75,0,52,0,0,0,0,0,0,0,43,0,44,0,53,0,195,0,111,0,78,0,57,0,186,0,255,0,44,0,0,0,206,0,206,0,80,0,121,0,160,0,113,0,1,0,0,0,10,0,0,0,34,0,173,0,157,0,167,0,119,0,174,0,121,0,135,0,42,0,29,0,0,0,213,0,251,0,0,0,0,0,191,0,33,0,0,0,219,0,66,0,65,0,60,0,123,0,197,0,176,0,0,0,109,0,184,0,108,0,149,0,142,0,143,0,33,0,50,0,142,0,238,0,115,0,152,0,233,0,177,0,22,0,240,0,0,0,163,0,217,0,88,0,166,0,240,0,247,0,184,0,138,0,216,0,134,0,0,0,0,0,0,0,200,0,0,0,147,0,5,0,0,0,43,0,0,0,176,0,198,0,57,0,148,0,0,0,70,0,95,0,171,0,70,0,39,0,0,0,11,0,0,0,8,0,162,0,33,0,8,0,109,0,214,0,0,0,19,0,239,0,96,0,0,0,162,0,25,0,0,0,75,0,148,0,0,0,66,0,242,0,145,0,0,0,196,0,25,0,62,0,112,0,6,0,66,0,32,0,0,0,50,0,160,0,0,0,42,0,185,0,171,0,95,0,225,0,53,0,0,0,239,0,0,0,148,0,233,0,0,0,167,0,0,0,249,0,0,0,212,0,172,0,237,0,0,0,0,0,113,0,0,0,227,0,127,0,46,0,246,0,97,0,202,0,0,0,0,0,203,0,183,0,7,0,241,0,111,0,0,0,17,0,209,0,42,0,125,0,68,0,253,0,238,0,57,0,142,0,0,0,204,0,236,0,127,0,219,0,154,0,0,0,37,0,190,0,0,0,151,0,225,0,99,0,162,0,55,0,0,0,227,0,129,0,142,0,210,0,213,0,243,0,175,0,2,0,162,0,30,0,131,0,242,0,0,0,0,0,26,0,153,0,49,0,0,0,0,0,0,0,67,0,242,0,0,0,160,0,53,0,121,0,219,0,125,0,160,0,96,0,30,0,91,0,233,0,0,0,185,0,130,0,0,0,0,0,0,0,0,0,216,0,0,0,64,0,113,0,144,0,47,0,124,0,0,0,164,0,0,0,17,0,225,0,0,0,101,0,5,0,96,0,153,0,153,0,0,0,190,0,221,0,66,0,4,0,17,0,0,0,0,0,122,0,255,0,14,0,84,0,94,0,22,0,103,0,41,0,1,0,70,0,0,0,48,0,138,0,230,0,0,0,80,0,167,0,106,0,27,0,0,0,18,0,90,0,147,0,119,0,104,0,240,0,0,0,234,0,127,0,60,0,25,0,242,0,88,0,7,0,4,0,88,0,241,0,39,0,204,0,185,0,0,0,76,0,142,0,193,0,25,0,224,0,156,0,248,0,0,0,0,0,178,0,47,0,42,0,0,0,54,0,78,0,114,0,0,0,119,0,181,0,44,0,0,0,82,0,146,0,168,0,228,0,122,0,151,0,0,0,46,0,42,0,82,0,189,0,147,0,115,0,168,0,43,0,196,0,211,0,127,0,79,0,49,0,225,0,0,0,56,0,9,0,0,0,5,0,194,0,50,0,168,0,54,0,83,0,50,0,151,0,0,0,12,0,78,0,32,0,233,0,211,0,0,0,0,0,0,0,107,0,4,0,87,0,129,0,43,0,21,0,221,0,26,0,5,0,0,0,144,0,29,0,6,0,0,0,0,0,24,0,9,0,150,0,0,0,115,0,206,0,106,0,0,0,77,0,0,0,196,0,136,0,0,0,237,0,98,0,50,0,164,0,206,0,149,0,0,0,0,0,22,0,226,0,9,0,129,0,0,0,53,0,79,0,53,0,71,0,202,0,181,0,80,0,0,0,0,0,0,0,192,0,177,0,21,0,0,0,217,0,122,0,144,0,0,0,0,0,0,0,143,0,0,0,198,0,87,0,152,0,246,0,0,0,20,0,171,0,165,0,166,0,0,0,30,0,76,0,114,0,240,0,203,0,251,0,50,0,216,0,0,0,150,0,0,0,28,0,217,0,231,0,220,0,0,0,3,0,255,0,47,0,154,0,82,0,229,0,0,0,104,0,196,0,0,0,226,0,173,0,0,0,89,0,188,0,58,0,194,0,226,0,25,0,69,0,74,0,240,0,109,0,154,0,191,0,252,0,157,0,4,0,0,0,200,0,87,0,88,0,26,0,49,0,49,0,33,0,14,0,0,0,42,0,235,0,81,0,145,0,0,0,152,0,0,0,131,0,0,0,67,0,0,0,38,0,234,0,94,0);
signal scenario_full  : scenario_type := (0,0,139,31,105,31,105,30,174,31,36,31,240,31,227,31,21,31,127,31,67,31,168,31,146,31,172,31,172,30,172,29,194,31,158,31,158,30,187,31,75,31,44,31,118,31,121,31,140,31,79,31,10,31,10,30,39,31,155,31,204,31,173,31,235,31,235,30,131,31,194,31,30,31,30,30,41,31,101,31,213,31,71,31,91,31,181,31,181,30,181,29,178,31,85,31,236,31,62,31,152,31,94,31,80,31,80,30,80,29,155,31,218,31,238,31,178,31,184,31,184,30,55,31,18,31,18,30,46,31,255,31,120,31,120,30,120,29,141,31,201,31,66,31,57,31,14,31,221,31,182,31,182,30,58,31,14,31,14,30,235,31,83,31,83,30,122,31,122,30,15,31,24,31,25,31,202,31,9,31,9,30,9,29,59,31,96,31,149,31,22,31,22,30,184,31,135,31,136,31,136,30,136,29,235,31,39,31,220,31,46,31,149,31,149,30,243,31,188,31,129,31,129,30,129,29,8,31,34,31,213,31,60,31,112,31,146,31,146,30,146,29,199,31,27,31,27,30,89,31,181,31,109,31,99,31,164,31,253,31,229,31,176,31,69,31,135,31,224,31,69,31,69,30,241,31,241,30,151,31,151,30,151,29,151,28,4,31,13,31,238,31,161,31,70,31,229,31,98,31,98,30,202,31,242,31,207,31,79,31,53,31,53,30,11,31,251,31,251,30,145,31,36,31,198,31,250,31,169,31,112,31,112,30,12,31,244,31,110,31,56,31,217,31,155,31,81,31,118,31,115,31,115,30,135,31,57,31,57,30,157,31,157,30,150,31,235,31,137,31,219,31,219,30,80,31,227,31,227,30,229,31,142,31,213,31,72,31,36,31,36,30,38,31,56,31,229,31,229,30,92,31,196,31,51,31,59,31,170,31,220,31,228,31,184,31,14,31,122,31,23,31,97,31,188,31,254,31,168,31,22,31,197,31,170,31,144,31,144,30,19,31,232,31,232,30,19,31,19,30,19,29,148,31,52,31,162,31,123,31,123,30,123,29,123,28,119,31,170,31,170,30,240,31,240,30,75,31,246,31,114,31,25,31,63,31,75,31,52,31,52,30,52,29,52,28,43,31,44,31,53,31,195,31,111,31,78,31,57,31,186,31,255,31,44,31,44,30,206,31,206,31,80,31,121,31,160,31,113,31,1,31,1,30,10,31,10,30,34,31,173,31,157,31,167,31,119,31,174,31,121,31,135,31,42,31,29,31,29,30,213,31,251,31,251,30,251,29,191,31,33,31,33,30,219,31,66,31,65,31,60,31,123,31,197,31,176,31,176,30,109,31,184,31,108,31,149,31,142,31,143,31,33,31,50,31,142,31,238,31,115,31,152,31,233,31,177,31,22,31,240,31,240,30,163,31,217,31,88,31,166,31,240,31,247,31,184,31,138,31,216,31,134,31,134,30,134,29,134,28,200,31,200,30,147,31,5,31,5,30,43,31,43,30,176,31,198,31,57,31,148,31,148,30,70,31,95,31,171,31,70,31,39,31,39,30,11,31,11,30,8,31,162,31,33,31,8,31,109,31,214,31,214,30,19,31,239,31,96,31,96,30,162,31,25,31,25,30,75,31,148,31,148,30,66,31,242,31,145,31,145,30,196,31,25,31,62,31,112,31,6,31,66,31,32,31,32,30,50,31,160,31,160,30,42,31,185,31,171,31,95,31,225,31,53,31,53,30,239,31,239,30,148,31,233,31,233,30,167,31,167,30,249,31,249,30,212,31,172,31,237,31,237,30,237,29,113,31,113,30,227,31,127,31,46,31,246,31,97,31,202,31,202,30,202,29,203,31,183,31,7,31,241,31,111,31,111,30,17,31,209,31,42,31,125,31,68,31,253,31,238,31,57,31,142,31,142,30,204,31,236,31,127,31,219,31,154,31,154,30,37,31,190,31,190,30,151,31,225,31,99,31,162,31,55,31,55,30,227,31,129,31,142,31,210,31,213,31,243,31,175,31,2,31,162,31,30,31,131,31,242,31,242,30,242,29,26,31,153,31,49,31,49,30,49,29,49,28,67,31,242,31,242,30,160,31,53,31,121,31,219,31,125,31,160,31,96,31,30,31,91,31,233,31,233,30,185,31,130,31,130,30,130,29,130,28,130,27,216,31,216,30,64,31,113,31,144,31,47,31,124,31,124,30,164,31,164,30,17,31,225,31,225,30,101,31,5,31,96,31,153,31,153,31,153,30,190,31,221,31,66,31,4,31,17,31,17,30,17,29,122,31,255,31,14,31,84,31,94,31,22,31,103,31,41,31,1,31,70,31,70,30,48,31,138,31,230,31,230,30,80,31,167,31,106,31,27,31,27,30,18,31,90,31,147,31,119,31,104,31,240,31,240,30,234,31,127,31,60,31,25,31,242,31,88,31,7,31,4,31,88,31,241,31,39,31,204,31,185,31,185,30,76,31,142,31,193,31,25,31,224,31,156,31,248,31,248,30,248,29,178,31,47,31,42,31,42,30,54,31,78,31,114,31,114,30,119,31,181,31,44,31,44,30,82,31,146,31,168,31,228,31,122,31,151,31,151,30,46,31,42,31,82,31,189,31,147,31,115,31,168,31,43,31,196,31,211,31,127,31,79,31,49,31,225,31,225,30,56,31,9,31,9,30,5,31,194,31,50,31,168,31,54,31,83,31,50,31,151,31,151,30,12,31,78,31,32,31,233,31,211,31,211,30,211,29,211,28,107,31,4,31,87,31,129,31,43,31,21,31,221,31,26,31,5,31,5,30,144,31,29,31,6,31,6,30,6,29,24,31,9,31,150,31,150,30,115,31,206,31,106,31,106,30,77,31,77,30,196,31,136,31,136,30,237,31,98,31,50,31,164,31,206,31,149,31,149,30,149,29,22,31,226,31,9,31,129,31,129,30,53,31,79,31,53,31,71,31,202,31,181,31,80,31,80,30,80,29,80,28,192,31,177,31,21,31,21,30,217,31,122,31,144,31,144,30,144,29,144,28,143,31,143,30,198,31,87,31,152,31,246,31,246,30,20,31,171,31,165,31,166,31,166,30,30,31,76,31,114,31,240,31,203,31,251,31,50,31,216,31,216,30,150,31,150,30,28,31,217,31,231,31,220,31,220,30,3,31,255,31,47,31,154,31,82,31,229,31,229,30,104,31,196,31,196,30,226,31,173,31,173,30,89,31,188,31,58,31,194,31,226,31,25,31,69,31,74,31,240,31,109,31,154,31,191,31,252,31,157,31,4,31,4,30,200,31,87,31,88,31,26,31,49,31,49,31,33,31,14,31,14,30,42,31,235,31,81,31,145,31,145,30,152,31,152,30,131,31,131,30,67,31,67,30,38,31,234,31,94,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
