-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_328 is
end project_tb_328;

architecture project_tb_arch_328 of project_tb_328 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 817;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (188,0,116,0,36,0,116,0,81,0,0,0,137,0,0,0,0,0,168,0,16,0,241,0,55,0,110,0,45,0,180,0,61,0,48,0,25,0,0,0,194,0,5,0,69,0,0,0,56,0,252,0,232,0,240,0,250,0,105,0,233,0,26,0,170,0,188,0,0,0,174,0,0,0,128,0,94,0,0,0,0,0,126,0,32,0,44,0,0,0,212,0,103,0,223,0,0,0,208,0,211,0,8,0,129,0,25,0,53,0,0,0,254,0,168,0,0,0,184,0,0,0,206,0,188,0,254,0,185,0,237,0,102,0,163,0,0,0,193,0,171,0,208,0,78,0,98,0,244,0,122,0,240,0,233,0,189,0,60,0,0,0,60,0,23,0,224,0,209,0,130,0,0,0,238,0,0,0,10,0,133,0,58,0,177,0,165,0,0,0,0,0,174,0,56,0,43,0,220,0,0,0,206,0,176,0,167,0,0,0,52,0,120,0,0,0,0,0,89,0,120,0,102,0,255,0,131,0,228,0,67,0,23,0,132,0,15,0,14,0,237,0,131,0,192,0,56,0,16,0,190,0,0,0,10,0,150,0,199,0,227,0,0,0,41,0,240,0,201,0,22,0,79,0,0,0,0,0,7,0,35,0,69,0,208,0,58,0,0,0,0,0,130,0,51,0,157,0,107,0,133,0,180,0,68,0,164,0,0,0,164,0,0,0,209,0,70,0,0,0,26,0,146,0,218,0,148,0,0,0,0,0,74,0,181,0,124,0,114,0,214,0,0,0,30,0,54,0,34,0,123,0,79,0,103,0,0,0,183,0,29,0,208,0,235,0,0,0,115,0,162,0,0,0,9,0,201,0,0,0,17,0,181,0,65,0,0,0,0,0,57,0,217,0,156,0,105,0,243,0,226,0,0,0,197,0,0,0,240,0,122,0,188,0,106,0,61,0,132,0,124,0,81,0,208,0,156,0,212,0,0,0,70,0,87,0,0,0,0,0,14,0,79,0,240,0,27,0,219,0,17,0,200,0,0,0,0,0,8,0,250,0,13,0,0,0,0,0,171,0,93,0,42,0,88,0,73,0,187,0,47,0,196,0,153,0,192,0,86,0,0,0,187,0,121,0,0,0,23,0,93,0,0,0,134,0,23,0,105,0,27,0,43,0,0,0,13,0,98,0,0,0,44,0,147,0,219,0,12,0,0,0,8,0,0,0,113,0,176,0,193,0,75,0,128,0,133,0,0,0,243,0,146,0,0,0,172,0,163,0,93,0,36,0,195,0,170,0,60,0,208,0,151,0,135,0,14,0,180,0,104,0,0,0,144,0,148,0,111,0,97,0,189,0,24,0,119,0,0,0,152,0,51,0,98,0,0,0,0,0,113,0,80,0,192,0,75,0,184,0,22,0,199,0,74,0,233,0,141,0,141,0,204,0,80,0,4,0,179,0,255,0,219,0,167,0,0,0,100,0,157,0,0,0,0,0,193,0,178,0,201,0,154,0,0,0,136,0,167,0,0,0,144,0,23,0,0,0,208,0,35,0,198,0,241,0,53,0,25,0,41,0,12,0,177,0,96,0,80,0,0,0,53,0,50,0,164,0,196,0,51,0,86,0,95,0,32,0,1,0,94,0,0,0,65,0,0,0,0,0,126,0,0,0,236,0,174,0,237,0,237,0,247,0,224,0,91,0,102,0,50,0,197,0,23,0,224,0,0,0,114,0,115,0,154,0,191,0,105,0,180,0,0,0,151,0,102,0,94,0,113,0,144,0,152,0,62,0,182,0,48,0,183,0,227,0,212,0,41,0,235,0,39,0,75,0,0,0,223,0,49,0,104,0,116,0,234,0,243,0,0,0,15,0,167,0,98,0,27,0,166,0,0,0,0,0,6,0,75,0,0,0,170,0,94,0,22,0,48,0,51,0,0,0,0,0,107,0,72,0,160,0,87,0,179,0,68,0,0,0,99,0,0,0,176,0,19,0,217,0,203,0,126,0,168,0,0,0,132,0,128,0,142,0,4,0,75,0,0,0,0,0,174,0,226,0,61,0,15,0,238,0,194,0,173,0,136,0,94,0,241,0,72,0,70,0,215,0,192,0,29,0,96,0,151,0,216,0,84,0,132,0,224,0,12,0,197,0,0,0,105,0,255,0,229,0,28,0,23,0,252,0,32,0,0,0,62,0,100,0,174,0,112,0,0,0,0,0,137,0,159,0,108,0,152,0,182,0,0,0,98,0,178,0,115,0,33,0,160,0,0,0,37,0,200,0,131,0,40,0,133,0,57,0,0,0,179,0,38,0,70,0,24,0,198,0,26,0,40,0,127,0,117,0,204,0,242,0,187,0,233,0,138,0,44,0,112,0,112,0,142,0,155,0,0,0,140,0,56,0,87,0,30,0,0,0,0,0,175,0,174,0,0,0,61,0,9,0,65,0,32,0,0,0,49,0,116,0,55,0,210,0,167,0,0,0,212,0,137,0,76,0,152,0,189,0,211,0,99,0,17,0,4,0,120,0,27,0,0,0,70,0,33,0,174,0,151,0,246,0,96,0,123,0,192,0,95,0,0,0,0,0,84,0,168,0,0,0,0,0,112,0,62,0,0,0,17,0,0,0,114,0,30,0,18,0,0,0,0,0,231,0,184,0,106,0,110,0,53,0,141,0,114,0,0,0,59,0,19,0,43,0,66,0,207,0,253,0,6,0,137,0,0,0,42,0,158,0,0,0,42,0,111,0,97,0,248,0,232,0,187,0,0,0,0,0,149,0,44,0,201,0,161,0,208,0,0,0,153,0,178,0,243,0,0,0,96,0,24,0,42,0,164,0,254,0,119,0,254,0,55,0,78,0,147,0,251,0,20,0,196,0,151,0,236,0,251,0,252,0,0,0,113,0,219,0,110,0,117,0,211,0,65,0,132,0,253,0,191,0,0,0,186,0,0,0,70,0,0,0,190,0,0,0,199,0,76,0,157,0,44,0,0,0,115,0,189,0,239,0,124,0,58,0,176,0,0,0,191,0,226,0,0,0,108,0,52,0,21,0,0,0,34,0,184,0,77,0,79,0,170,0,55,0,123,0,54,0,149,0,174,0,0,0,0,0,32,0,16,0,0,0,0,0,72,0,12,0,106,0,64,0,60,0,219,0,0,0,0,0,131,0,150,0,116,0,130,0,117,0,237,0,74,0,0,0,20,0,19,0,209,0,203,0,63,0,231,0,219,0,89,0,48,0,0,0,143,0,175,0,157,0,57,0,163,0,203,0,74,0,177,0,233,0,181,0,0,0,145,0,234,0,0,0,72,0,144,0,255,0,16,0,168,0,7,0,128,0,159,0,232,0,134,0,220,0,0,0,74,0,58,0,125,0,232,0,163,0,184,0,200,0,30,0,0,0,0,0,13,0,178,0,241,0,112,0,115,0,61,0,0,0,0,0,155,0,219,0,69,0,70,0,59,0,126,0,0,0,0,0,20,0,204,0,183,0,0,0,135,0,111,0,74,0,42,0,78,0,248,0,216,0,120,0,29,0,101,0,17,0,90,0,62,0,0,0,0,0,160,0,124,0,0,0,235,0,248,0,165,0,0,0,230,0,159,0,215,0,156,0,82,0,180,0,222,0,68,0,0,0,0,0,139,0,29,0,65,0,235,0,11,0,0,0,85,0,62,0,0,0,158,0,45,0);
signal scenario_full  : scenario_type := (188,31,116,31,36,31,116,31,81,31,81,30,137,31,137,30,137,29,168,31,16,31,241,31,55,31,110,31,45,31,180,31,61,31,48,31,25,31,25,30,194,31,5,31,69,31,69,30,56,31,252,31,232,31,240,31,250,31,105,31,233,31,26,31,170,31,188,31,188,30,174,31,174,30,128,31,94,31,94,30,94,29,126,31,32,31,44,31,44,30,212,31,103,31,223,31,223,30,208,31,211,31,8,31,129,31,25,31,53,31,53,30,254,31,168,31,168,30,184,31,184,30,206,31,188,31,254,31,185,31,237,31,102,31,163,31,163,30,193,31,171,31,208,31,78,31,98,31,244,31,122,31,240,31,233,31,189,31,60,31,60,30,60,31,23,31,224,31,209,31,130,31,130,30,238,31,238,30,10,31,133,31,58,31,177,31,165,31,165,30,165,29,174,31,56,31,43,31,220,31,220,30,206,31,176,31,167,31,167,30,52,31,120,31,120,30,120,29,89,31,120,31,102,31,255,31,131,31,228,31,67,31,23,31,132,31,15,31,14,31,237,31,131,31,192,31,56,31,16,31,190,31,190,30,10,31,150,31,199,31,227,31,227,30,41,31,240,31,201,31,22,31,79,31,79,30,79,29,7,31,35,31,69,31,208,31,58,31,58,30,58,29,130,31,51,31,157,31,107,31,133,31,180,31,68,31,164,31,164,30,164,31,164,30,209,31,70,31,70,30,26,31,146,31,218,31,148,31,148,30,148,29,74,31,181,31,124,31,114,31,214,31,214,30,30,31,54,31,34,31,123,31,79,31,103,31,103,30,183,31,29,31,208,31,235,31,235,30,115,31,162,31,162,30,9,31,201,31,201,30,17,31,181,31,65,31,65,30,65,29,57,31,217,31,156,31,105,31,243,31,226,31,226,30,197,31,197,30,240,31,122,31,188,31,106,31,61,31,132,31,124,31,81,31,208,31,156,31,212,31,212,30,70,31,87,31,87,30,87,29,14,31,79,31,240,31,27,31,219,31,17,31,200,31,200,30,200,29,8,31,250,31,13,31,13,30,13,29,171,31,93,31,42,31,88,31,73,31,187,31,47,31,196,31,153,31,192,31,86,31,86,30,187,31,121,31,121,30,23,31,93,31,93,30,134,31,23,31,105,31,27,31,43,31,43,30,13,31,98,31,98,30,44,31,147,31,219,31,12,31,12,30,8,31,8,30,113,31,176,31,193,31,75,31,128,31,133,31,133,30,243,31,146,31,146,30,172,31,163,31,93,31,36,31,195,31,170,31,60,31,208,31,151,31,135,31,14,31,180,31,104,31,104,30,144,31,148,31,111,31,97,31,189,31,24,31,119,31,119,30,152,31,51,31,98,31,98,30,98,29,113,31,80,31,192,31,75,31,184,31,22,31,199,31,74,31,233,31,141,31,141,31,204,31,80,31,4,31,179,31,255,31,219,31,167,31,167,30,100,31,157,31,157,30,157,29,193,31,178,31,201,31,154,31,154,30,136,31,167,31,167,30,144,31,23,31,23,30,208,31,35,31,198,31,241,31,53,31,25,31,41,31,12,31,177,31,96,31,80,31,80,30,53,31,50,31,164,31,196,31,51,31,86,31,95,31,32,31,1,31,94,31,94,30,65,31,65,30,65,29,126,31,126,30,236,31,174,31,237,31,237,31,247,31,224,31,91,31,102,31,50,31,197,31,23,31,224,31,224,30,114,31,115,31,154,31,191,31,105,31,180,31,180,30,151,31,102,31,94,31,113,31,144,31,152,31,62,31,182,31,48,31,183,31,227,31,212,31,41,31,235,31,39,31,75,31,75,30,223,31,49,31,104,31,116,31,234,31,243,31,243,30,15,31,167,31,98,31,27,31,166,31,166,30,166,29,6,31,75,31,75,30,170,31,94,31,22,31,48,31,51,31,51,30,51,29,107,31,72,31,160,31,87,31,179,31,68,31,68,30,99,31,99,30,176,31,19,31,217,31,203,31,126,31,168,31,168,30,132,31,128,31,142,31,4,31,75,31,75,30,75,29,174,31,226,31,61,31,15,31,238,31,194,31,173,31,136,31,94,31,241,31,72,31,70,31,215,31,192,31,29,31,96,31,151,31,216,31,84,31,132,31,224,31,12,31,197,31,197,30,105,31,255,31,229,31,28,31,23,31,252,31,32,31,32,30,62,31,100,31,174,31,112,31,112,30,112,29,137,31,159,31,108,31,152,31,182,31,182,30,98,31,178,31,115,31,33,31,160,31,160,30,37,31,200,31,131,31,40,31,133,31,57,31,57,30,179,31,38,31,70,31,24,31,198,31,26,31,40,31,127,31,117,31,204,31,242,31,187,31,233,31,138,31,44,31,112,31,112,31,142,31,155,31,155,30,140,31,56,31,87,31,30,31,30,30,30,29,175,31,174,31,174,30,61,31,9,31,65,31,32,31,32,30,49,31,116,31,55,31,210,31,167,31,167,30,212,31,137,31,76,31,152,31,189,31,211,31,99,31,17,31,4,31,120,31,27,31,27,30,70,31,33,31,174,31,151,31,246,31,96,31,123,31,192,31,95,31,95,30,95,29,84,31,168,31,168,30,168,29,112,31,62,31,62,30,17,31,17,30,114,31,30,31,18,31,18,30,18,29,231,31,184,31,106,31,110,31,53,31,141,31,114,31,114,30,59,31,19,31,43,31,66,31,207,31,253,31,6,31,137,31,137,30,42,31,158,31,158,30,42,31,111,31,97,31,248,31,232,31,187,31,187,30,187,29,149,31,44,31,201,31,161,31,208,31,208,30,153,31,178,31,243,31,243,30,96,31,24,31,42,31,164,31,254,31,119,31,254,31,55,31,78,31,147,31,251,31,20,31,196,31,151,31,236,31,251,31,252,31,252,30,113,31,219,31,110,31,117,31,211,31,65,31,132,31,253,31,191,31,191,30,186,31,186,30,70,31,70,30,190,31,190,30,199,31,76,31,157,31,44,31,44,30,115,31,189,31,239,31,124,31,58,31,176,31,176,30,191,31,226,31,226,30,108,31,52,31,21,31,21,30,34,31,184,31,77,31,79,31,170,31,55,31,123,31,54,31,149,31,174,31,174,30,174,29,32,31,16,31,16,30,16,29,72,31,12,31,106,31,64,31,60,31,219,31,219,30,219,29,131,31,150,31,116,31,130,31,117,31,237,31,74,31,74,30,20,31,19,31,209,31,203,31,63,31,231,31,219,31,89,31,48,31,48,30,143,31,175,31,157,31,57,31,163,31,203,31,74,31,177,31,233,31,181,31,181,30,145,31,234,31,234,30,72,31,144,31,255,31,16,31,168,31,7,31,128,31,159,31,232,31,134,31,220,31,220,30,74,31,58,31,125,31,232,31,163,31,184,31,200,31,30,31,30,30,30,29,13,31,178,31,241,31,112,31,115,31,61,31,61,30,61,29,155,31,219,31,69,31,70,31,59,31,126,31,126,30,126,29,20,31,204,31,183,31,183,30,135,31,111,31,74,31,42,31,78,31,248,31,216,31,120,31,29,31,101,31,17,31,90,31,62,31,62,30,62,29,160,31,124,31,124,30,235,31,248,31,165,31,165,30,230,31,159,31,215,31,156,31,82,31,180,31,222,31,68,31,68,30,68,29,139,31,29,31,65,31,235,31,11,31,11,30,85,31,62,31,62,30,158,31,45,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
