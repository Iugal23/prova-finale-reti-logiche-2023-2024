-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 892;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (106,0,210,0,249,0,34,0,79,0,0,0,179,0,0,0,103,0,63,0,62,0,0,0,120,0,57,0,0,0,34,0,0,0,0,0,165,0,29,0,62,0,244,0,5,0,240,0,167,0,0,0,161,0,48,0,92,0,3,0,0,0,184,0,88,0,41,0,0,0,165,0,37,0,79,0,0,0,208,0,136,0,189,0,52,0,0,0,0,0,28,0,62,0,216,0,0,0,229,0,186,0,208,0,16,0,171,0,67,0,64,0,74,0,154,0,110,0,90,0,40,0,115,0,31,0,0,0,177,0,80,0,190,0,181,0,0,0,131,0,172,0,124,0,0,0,72,0,237,0,0,0,70,0,181,0,59,0,14,0,71,0,237,0,202,0,162,0,235,0,87,0,0,0,70,0,40,0,0,0,74,0,0,0,79,0,4,0,98,0,73,0,0,0,0,0,175,0,0,0,114,0,99,0,227,0,0,0,151,0,90,0,165,0,43,0,132,0,0,0,162,0,36,0,19,0,127,0,0,0,137,0,20,0,48,0,98,0,30,0,4,0,214,0,79,0,62,0,0,0,234,0,115,0,5,0,0,0,0,0,0,0,195,0,0,0,0,0,188,0,31,0,16,0,93,0,232,0,244,0,212,0,108,0,137,0,212,0,245,0,165,0,0,0,171,0,224,0,234,0,133,0,52,0,51,0,129,0,165,0,170,0,212,0,0,0,252,0,106,0,40,0,171,0,0,0,178,0,26,0,141,0,117,0,174,0,228,0,246,0,0,0,0,0,113,0,15,0,61,0,0,0,0,0,0,0,76,0,130,0,85,0,192,0,0,0,249,0,191,0,131,0,0,0,37,0,164,0,0,0,94,0,0,0,28,0,198,0,243,0,189,0,0,0,90,0,146,0,0,0,0,0,32,0,117,0,0,0,221,0,252,0,0,0,86,0,0,0,238,0,116,0,61,0,132,0,102,0,188,0,128,0,136,0,63,0,0,0,37,0,113,0,239,0,142,0,235,0,220,0,175,0,217,0,136,0,12,0,46,0,0,0,126,0,12,0,224,0,54,0,95,0,50,0,212,0,182,0,203,0,0,0,54,0,202,0,0,0,0,0,254,0,3,0,8,0,161,0,137,0,0,0,176,0,0,0,113,0,88,0,167,0,0,0,100,0,144,0,107,0,231,0,26,0,208,0,0,0,24,0,13,0,59,0,45,0,226,0,0,0,69,0,186,0,0,0,6,0,60,0,0,0,158,0,123,0,247,0,172,0,196,0,153,0,196,0,232,0,76,0,210,0,234,0,182,0,151,0,87,0,251,0,27,0,181,0,164,0,0,0,194,0,76,0,249,0,0,0,138,0,27,0,0,0,141,0,213,0,1,0,157,0,242,0,189,0,0,0,245,0,179,0,195,0,90,0,0,0,143,0,248,0,252,0,157,0,49,0,26,0,60,0,0,0,79,0,0,0,0,0,236,0,32,0,209,0,120,0,0,0,0,0,123,0,0,0,0,0,0,0,82,0,56,0,0,0,82,0,234,0,207,0,114,0,167,0,150,0,28,0,94,0,32,0,0,0,43,0,123,0,244,0,204,0,239,0,0,0,133,0,0,0,210,0,146,0,171,0,62,0,186,0,4,0,146,0,255,0,68,0,146,0,166,0,0,0,227,0,159,0,43,0,0,0,220,0,8,0,187,0,0,0,106,0,0,0,157,0,101,0,66,0,245,0,0,0,0,0,151,0,136,0,68,0,0,0,0,0,62,0,224,0,253,0,143,0,115,0,100,0,72,0,0,0,36,0,191,0,0,0,45,0,130,0,255,0,61,0,4,0,101,0,225,0,186,0,0,0,180,0,68,0,0,0,207,0,201,0,147,0,10,0,170,0,23,0,39,0,157,0,153,0,111,0,244,0,182,0,129,0,117,0,175,0,161,0,0,0,0,0,153,0,159,0,161,0,0,0,7,0,88,0,19,0,96,0,213,0,50,0,74,0,173,0,158,0,210,0,81,0,202,0,62,0,0,0,94,0,241,0,0,0,134,0,157,0,251,0,249,0,133,0,253,0,69,0,0,0,125,0,146,0,169,0,0,0,66,0,113,0,218,0,83,0,124,0,39,0,0,0,18,0,101,0,61,0,220,0,177,0,90,0,4,0,228,0,172,0,74,0,27,0,0,0,235,0,0,0,49,0,128,0,203,0,97,0,150,0,57,0,0,0,28,0,33,0,237,0,46,0,75,0,138,0,20,0,34,0,44,0,237,0,0,0,66,0,86,0,0,0,128,0,206,0,0,0,16,0,52,0,31,0,62,0,105,0,73,0,55,0,153,0,219,0,160,0,25,0,0,0,240,0,150,0,134,0,11,0,223,0,48,0,0,0,11,0,194,0,14,0,80,0,31,0,66,0,241,0,238,0,252,0,36,0,0,0,78,0,233,0,0,0,5,0,130,0,104,0,0,0,0,0,192,0,46,0,0,0,235,0,0,0,103,0,151,0,117,0,177,0,0,0,210,0,0,0,57,0,65,0,144,0,0,0,220,0,89,0,159,0,0,0,0,0,240,0,0,0,0,0,188,0,0,0,29,0,84,0,35,0,62,0,80,0,45,0,97,0,43,0,246,0,0,0,71,0,113,0,0,0,200,0,252,0,0,0,249,0,0,0,0,0,0,0,124,0,183,0,181,0,146,0,113,0,251,0,49,0,0,0,9,0,10,0,132,0,224,0,100,0,1,0,226,0,116,0,0,0,174,0,104,0,68,0,223,0,182,0,162,0,98,0,167,0,118,0,92,0,251,0,142,0,0,0,0,0,0,0,0,0,233,0,235,0,66,0,42,0,169,0,204,0,0,0,65,0,123,0,27,0,158,0,116,0,0,0,0,0,126,0,0,0,12,0,117,0,121,0,18,0,219,0,164,0,19,0,16,0,110,0,0,0,38,0,30,0,136,0,241,0,119,0,189,0,12,0,56,0,213,0,38,0,0,0,172,0,0,0,184,0,96,0,33,0,195,0,164,0,32,0,212,0,14,0,47,0,0,0,218,0,13,0,36,0,232,0,0,0,131,0,0,0,0,0,37,0,110,0,19,0,182,0,0,0,0,0,209,0,122,0,208,0,47,0,25,0,6,0,196,0,144,0,59,0,0,0,73,0,199,0,126,0,61,0,0,0,0,0,134,0,221,0,0,0,0,0,0,0,0,0,53,0,0,0,219,0,216,0,133,0,119,0,219,0,190,0,57,0,181,0,217,0,216,0,163,0,0,0,28,0,128,0,122,0,0,0,221,0,0,0,155,0,0,0,0,0,0,0,0,0,148,0,95,0,157,0,64,0,123,0,80,0,200,0,192,0,0,0,156,0,216,0,36,0,164,0,55,0,160,0,7,0,43,0,0,0,29,0,136,0,199,0,204,0,167,0,17,0,205,0,0,0,237,0,0,0,146,0,112,0,32,0,216,0,99,0,210,0,0,0,133,0,46,0,231,0,142,0,189,0,0,0,49,0,98,0,237,0,191,0,77,0,16,0,109,0,65,0,10,0,214,0,41,0,23,0,208,0,19,0,144,0,32,0,103,0,253,0,20,0,0,0,246,0,19,0,3,0,186,0,125,0,217,0,104,0,0,0,0,0,109,0,15,0,0,0,190,0,197,0,43,0,217,0,242,0,0,0,184,0,197,0,57,0,224,0,15,0,119,0,0,0,99,0,241,0,26,0,0,0,0,0,125,0,0,0,143,0,186,0,195,0,0,0,235,0,32,0,45,0,67,0,51,0,11,0,120,0,187,0,40,0,153,0,142,0,7,0,0,0,116,0,164,0,110,0,93,0,70,0,99,0,57,0,240,0,6,0,27,0,138,0,3,0,224,0,2,0,0,0,209,0,208,0,99,0,18,0,36,0,1,0,31,0,0,0,60,0,8,0,0,0,35,0,0,0,182,0,0,0,17,0,0,0,57,0,0,0,58,0,214,0,208,0,7,0,26,0,182,0,202,0,0,0,191,0,31,0,22,0,90,0,0,0);
signal scenario_full  : scenario_type := (106,31,210,31,249,31,34,31,79,31,79,30,179,31,179,30,103,31,63,31,62,31,62,30,120,31,57,31,57,30,34,31,34,30,34,29,165,31,29,31,62,31,244,31,5,31,240,31,167,31,167,30,161,31,48,31,92,31,3,31,3,30,184,31,88,31,41,31,41,30,165,31,37,31,79,31,79,30,208,31,136,31,189,31,52,31,52,30,52,29,28,31,62,31,216,31,216,30,229,31,186,31,208,31,16,31,171,31,67,31,64,31,74,31,154,31,110,31,90,31,40,31,115,31,31,31,31,30,177,31,80,31,190,31,181,31,181,30,131,31,172,31,124,31,124,30,72,31,237,31,237,30,70,31,181,31,59,31,14,31,71,31,237,31,202,31,162,31,235,31,87,31,87,30,70,31,40,31,40,30,74,31,74,30,79,31,4,31,98,31,73,31,73,30,73,29,175,31,175,30,114,31,99,31,227,31,227,30,151,31,90,31,165,31,43,31,132,31,132,30,162,31,36,31,19,31,127,31,127,30,137,31,20,31,48,31,98,31,30,31,4,31,214,31,79,31,62,31,62,30,234,31,115,31,5,31,5,30,5,29,5,28,195,31,195,30,195,29,188,31,31,31,16,31,93,31,232,31,244,31,212,31,108,31,137,31,212,31,245,31,165,31,165,30,171,31,224,31,234,31,133,31,52,31,51,31,129,31,165,31,170,31,212,31,212,30,252,31,106,31,40,31,171,31,171,30,178,31,26,31,141,31,117,31,174,31,228,31,246,31,246,30,246,29,113,31,15,31,61,31,61,30,61,29,61,28,76,31,130,31,85,31,192,31,192,30,249,31,191,31,131,31,131,30,37,31,164,31,164,30,94,31,94,30,28,31,198,31,243,31,189,31,189,30,90,31,146,31,146,30,146,29,32,31,117,31,117,30,221,31,252,31,252,30,86,31,86,30,238,31,116,31,61,31,132,31,102,31,188,31,128,31,136,31,63,31,63,30,37,31,113,31,239,31,142,31,235,31,220,31,175,31,217,31,136,31,12,31,46,31,46,30,126,31,12,31,224,31,54,31,95,31,50,31,212,31,182,31,203,31,203,30,54,31,202,31,202,30,202,29,254,31,3,31,8,31,161,31,137,31,137,30,176,31,176,30,113,31,88,31,167,31,167,30,100,31,144,31,107,31,231,31,26,31,208,31,208,30,24,31,13,31,59,31,45,31,226,31,226,30,69,31,186,31,186,30,6,31,60,31,60,30,158,31,123,31,247,31,172,31,196,31,153,31,196,31,232,31,76,31,210,31,234,31,182,31,151,31,87,31,251,31,27,31,181,31,164,31,164,30,194,31,76,31,249,31,249,30,138,31,27,31,27,30,141,31,213,31,1,31,157,31,242,31,189,31,189,30,245,31,179,31,195,31,90,31,90,30,143,31,248,31,252,31,157,31,49,31,26,31,60,31,60,30,79,31,79,30,79,29,236,31,32,31,209,31,120,31,120,30,120,29,123,31,123,30,123,29,123,28,82,31,56,31,56,30,82,31,234,31,207,31,114,31,167,31,150,31,28,31,94,31,32,31,32,30,43,31,123,31,244,31,204,31,239,31,239,30,133,31,133,30,210,31,146,31,171,31,62,31,186,31,4,31,146,31,255,31,68,31,146,31,166,31,166,30,227,31,159,31,43,31,43,30,220,31,8,31,187,31,187,30,106,31,106,30,157,31,101,31,66,31,245,31,245,30,245,29,151,31,136,31,68,31,68,30,68,29,62,31,224,31,253,31,143,31,115,31,100,31,72,31,72,30,36,31,191,31,191,30,45,31,130,31,255,31,61,31,4,31,101,31,225,31,186,31,186,30,180,31,68,31,68,30,207,31,201,31,147,31,10,31,170,31,23,31,39,31,157,31,153,31,111,31,244,31,182,31,129,31,117,31,175,31,161,31,161,30,161,29,153,31,159,31,161,31,161,30,7,31,88,31,19,31,96,31,213,31,50,31,74,31,173,31,158,31,210,31,81,31,202,31,62,31,62,30,94,31,241,31,241,30,134,31,157,31,251,31,249,31,133,31,253,31,69,31,69,30,125,31,146,31,169,31,169,30,66,31,113,31,218,31,83,31,124,31,39,31,39,30,18,31,101,31,61,31,220,31,177,31,90,31,4,31,228,31,172,31,74,31,27,31,27,30,235,31,235,30,49,31,128,31,203,31,97,31,150,31,57,31,57,30,28,31,33,31,237,31,46,31,75,31,138,31,20,31,34,31,44,31,237,31,237,30,66,31,86,31,86,30,128,31,206,31,206,30,16,31,52,31,31,31,62,31,105,31,73,31,55,31,153,31,219,31,160,31,25,31,25,30,240,31,150,31,134,31,11,31,223,31,48,31,48,30,11,31,194,31,14,31,80,31,31,31,66,31,241,31,238,31,252,31,36,31,36,30,78,31,233,31,233,30,5,31,130,31,104,31,104,30,104,29,192,31,46,31,46,30,235,31,235,30,103,31,151,31,117,31,177,31,177,30,210,31,210,30,57,31,65,31,144,31,144,30,220,31,89,31,159,31,159,30,159,29,240,31,240,30,240,29,188,31,188,30,29,31,84,31,35,31,62,31,80,31,45,31,97,31,43,31,246,31,246,30,71,31,113,31,113,30,200,31,252,31,252,30,249,31,249,30,249,29,249,28,124,31,183,31,181,31,146,31,113,31,251,31,49,31,49,30,9,31,10,31,132,31,224,31,100,31,1,31,226,31,116,31,116,30,174,31,104,31,68,31,223,31,182,31,162,31,98,31,167,31,118,31,92,31,251,31,142,31,142,30,142,29,142,28,142,27,233,31,235,31,66,31,42,31,169,31,204,31,204,30,65,31,123,31,27,31,158,31,116,31,116,30,116,29,126,31,126,30,12,31,117,31,121,31,18,31,219,31,164,31,19,31,16,31,110,31,110,30,38,31,30,31,136,31,241,31,119,31,189,31,12,31,56,31,213,31,38,31,38,30,172,31,172,30,184,31,96,31,33,31,195,31,164,31,32,31,212,31,14,31,47,31,47,30,218,31,13,31,36,31,232,31,232,30,131,31,131,30,131,29,37,31,110,31,19,31,182,31,182,30,182,29,209,31,122,31,208,31,47,31,25,31,6,31,196,31,144,31,59,31,59,30,73,31,199,31,126,31,61,31,61,30,61,29,134,31,221,31,221,30,221,29,221,28,221,27,53,31,53,30,219,31,216,31,133,31,119,31,219,31,190,31,57,31,181,31,217,31,216,31,163,31,163,30,28,31,128,31,122,31,122,30,221,31,221,30,155,31,155,30,155,29,155,28,155,27,148,31,95,31,157,31,64,31,123,31,80,31,200,31,192,31,192,30,156,31,216,31,36,31,164,31,55,31,160,31,7,31,43,31,43,30,29,31,136,31,199,31,204,31,167,31,17,31,205,31,205,30,237,31,237,30,146,31,112,31,32,31,216,31,99,31,210,31,210,30,133,31,46,31,231,31,142,31,189,31,189,30,49,31,98,31,237,31,191,31,77,31,16,31,109,31,65,31,10,31,214,31,41,31,23,31,208,31,19,31,144,31,32,31,103,31,253,31,20,31,20,30,246,31,19,31,3,31,186,31,125,31,217,31,104,31,104,30,104,29,109,31,15,31,15,30,190,31,197,31,43,31,217,31,242,31,242,30,184,31,197,31,57,31,224,31,15,31,119,31,119,30,99,31,241,31,26,31,26,30,26,29,125,31,125,30,143,31,186,31,195,31,195,30,235,31,32,31,45,31,67,31,51,31,11,31,120,31,187,31,40,31,153,31,142,31,7,31,7,30,116,31,164,31,110,31,93,31,70,31,99,31,57,31,240,31,6,31,27,31,138,31,3,31,224,31,2,31,2,30,209,31,208,31,99,31,18,31,36,31,1,31,31,31,31,30,60,31,8,31,8,30,35,31,35,30,182,31,182,30,17,31,17,30,57,31,57,30,58,31,214,31,208,31,7,31,26,31,182,31,202,31,202,30,191,31,31,31,22,31,90,31,90,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
