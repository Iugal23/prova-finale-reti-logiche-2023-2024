-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_577 is
end project_tb_577;

architecture project_tb_arch_577 of project_tb_577 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 577;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (222,0,15,0,90,0,201,0,154,0,0,0,200,0,209,0,28,0,153,0,0,0,9,0,68,0,222,0,0,0,216,0,187,0,132,0,0,0,182,0,19,0,36,0,174,0,0,0,160,0,182,0,218,0,62,0,106,0,204,0,45,0,0,0,169,0,41,0,200,0,1,0,196,0,127,0,170,0,128,0,132,0,183,0,36,0,216,0,141,0,0,0,103,0,0,0,68,0,230,0,0,0,0,0,0,0,44,0,197,0,85,0,72,0,176,0,113,0,15,0,0,0,43,0,243,0,0,0,0,0,86,0,201,0,0,0,115,0,0,0,206,0,127,0,90,0,9,0,233,0,220,0,0,0,240,0,178,0,167,0,187,0,3,0,245,0,0,0,54,0,4,0,184,0,0,0,69,0,5,0,61,0,47,0,92,0,0,0,246,0,112,0,150,0,19,0,138,0,138,0,199,0,37,0,116,0,3,0,137,0,124,0,107,0,125,0,132,0,112,0,248,0,100,0,205,0,16,0,10,0,72,0,174,0,133,0,195,0,0,0,0,0,10,0,95,0,147,0,223,0,244,0,255,0,48,0,172,0,177,0,167,0,166,0,144,0,187,0,23,0,140,0,91,0,0,0,115,0,88,0,80,0,109,0,161,0,57,0,186,0,86,0,0,0,176,0,244,0,2,0,0,0,57,0,0,0,112,0,0,0,116,0,225,0,230,0,143,0,69,0,184,0,217,0,210,0,219,0,25,0,230,0,119,0,0,0,3,0,0,0,78,0,229,0,242,0,185,0,132,0,213,0,17,0,154,0,142,0,29,0,234,0,33,0,173,0,5,0,249,0,0,0,218,0,23,0,0,0,104,0,115,0,0,0,141,0,233,0,128,0,0,0,26,0,161,0,82,0,154,0,21,0,149,0,20,0,178,0,84,0,46,0,0,0,0,0,201,0,0,0,167,0,26,0,13,0,137,0,121,0,43,0,25,0,79,0,65,0,19,0,247,0,83,0,148,0,76,0,253,0,0,0,42,0,84,0,0,0,0,0,220,0,0,0,0,0,45,0,0,0,65,0,195,0,210,0,80,0,36,0,107,0,7,0,0,0,18,0,32,0,90,0,160,0,254,0,99,0,44,0,212,0,0,0,98,0,248,0,10,0,13,0,140,0,188,0,231,0,86,0,190,0,121,0,54,0,134,0,255,0,48,0,140,0,6,0,36,0,204,0,49,0,246,0,231,0,127,0,186,0,96,0,7,0,81,0,0,0,246,0,0,0,0,0,85,0,0,0,131,0,0,0,0,0,109,0,166,0,193,0,10,0,64,0,80,0,252,0,71,0,225,0,54,0,165,0,0,0,67,0,153,0,31,0,216,0,106,0,60,0,177,0,77,0,214,0,126,0,111,0,203,0,71,0,73,0,193,0,52,0,218,0,160,0,0,0,228,0,167,0,113,0,158,0,11,0,14,0,0,0,94,0,117,0,127,0,54,0,0,0,38,0,34,0,221,0,20,0,202,0,29,0,10,0,187,0,105,0,51,0,65,0,241,0,91,0,62,0,191,0,240,0,0,0,245,0,238,0,204,0,120,0,0,0,145,0,171,0,209,0,19,0,70,0,87,0,212,0,8,0,0,0,221,0,156,0,69,0,0,0,0,0,33,0,146,0,200,0,39,0,85,0,197,0,172,0,186,0,117,0,186,0,50,0,94,0,0,0,67,0,119,0,5,0,165,0,250,0,0,0,235,0,183,0,25,0,24,0,0,0,118,0,15,0,216,0,0,0,68,0,61,0,231,0,44,0,219,0,60,0,52,0,0,0,190,0,230,0,153,0,0,0,165,0,105,0,28,0,98,0,0,0,196,0,183,0,201,0,167,0,224,0,172,0,0,0,219,0,213,0,158,0,248,0,132,0,0,0,57,0,246,0,71,0,161,0,121,0,0,0,56,0,107,0,0,0,65,0,131,0,79,0,0,0,16,0,100,0,22,0,141,0,101,0,232,0,199,0,156,0,238,0,61,0,235,0,0,0,225,0,0,0,0,0,7,0,15,0,58,0,37,0,97,0,188,0,164,0,244,0,205,0,108,0,35,0,210,0,0,0,0,0,128,0,99,0,0,0,66,0,0,0,207,0,26,0,123,0,175,0,209,0,24,0,175,0,0,0,218,0,0,0,155,0,245,0,216,0,109,0,209,0,97,0,88,0,252,0,0,0,179,0,242,0,10,0,160,0,0,0,38,0,242,0,88,0,223,0,155,0,56,0,112,0,0,0,0,0,129,0,0,0,0,0,141,0,252,0,0,0,109,0,221,0,43,0,148,0,206,0,174,0,71,0,81,0,119,0,0,0,73,0,164,0,216,0,128,0,207,0,228,0,173,0,121,0,108,0,43,0,53,0,251,0,25,0,92,0,207,0,174,0,210,0,28,0,0,0,191,0,0,0,162,0,114,0,106,0,0,0,40,0,109,0,29,0,114,0,0,0,18,0,103,0,228,0,0,0,193,0,0,0,89,0,102,0,118,0,179,0,50,0,254,0,192,0,28,0,206,0,78,0,117,0,192,0,64,0,0,0,0,0,21,0,51,0,0,0,49,0,88,0,199,0);
signal scenario_full  : scenario_type := (222,31,15,31,90,31,201,31,154,31,154,30,200,31,209,31,28,31,153,31,153,30,9,31,68,31,222,31,222,30,216,31,187,31,132,31,132,30,182,31,19,31,36,31,174,31,174,30,160,31,182,31,218,31,62,31,106,31,204,31,45,31,45,30,169,31,41,31,200,31,1,31,196,31,127,31,170,31,128,31,132,31,183,31,36,31,216,31,141,31,141,30,103,31,103,30,68,31,230,31,230,30,230,29,230,28,44,31,197,31,85,31,72,31,176,31,113,31,15,31,15,30,43,31,243,31,243,30,243,29,86,31,201,31,201,30,115,31,115,30,206,31,127,31,90,31,9,31,233,31,220,31,220,30,240,31,178,31,167,31,187,31,3,31,245,31,245,30,54,31,4,31,184,31,184,30,69,31,5,31,61,31,47,31,92,31,92,30,246,31,112,31,150,31,19,31,138,31,138,31,199,31,37,31,116,31,3,31,137,31,124,31,107,31,125,31,132,31,112,31,248,31,100,31,205,31,16,31,10,31,72,31,174,31,133,31,195,31,195,30,195,29,10,31,95,31,147,31,223,31,244,31,255,31,48,31,172,31,177,31,167,31,166,31,144,31,187,31,23,31,140,31,91,31,91,30,115,31,88,31,80,31,109,31,161,31,57,31,186,31,86,31,86,30,176,31,244,31,2,31,2,30,57,31,57,30,112,31,112,30,116,31,225,31,230,31,143,31,69,31,184,31,217,31,210,31,219,31,25,31,230,31,119,31,119,30,3,31,3,30,78,31,229,31,242,31,185,31,132,31,213,31,17,31,154,31,142,31,29,31,234,31,33,31,173,31,5,31,249,31,249,30,218,31,23,31,23,30,104,31,115,31,115,30,141,31,233,31,128,31,128,30,26,31,161,31,82,31,154,31,21,31,149,31,20,31,178,31,84,31,46,31,46,30,46,29,201,31,201,30,167,31,26,31,13,31,137,31,121,31,43,31,25,31,79,31,65,31,19,31,247,31,83,31,148,31,76,31,253,31,253,30,42,31,84,31,84,30,84,29,220,31,220,30,220,29,45,31,45,30,65,31,195,31,210,31,80,31,36,31,107,31,7,31,7,30,18,31,32,31,90,31,160,31,254,31,99,31,44,31,212,31,212,30,98,31,248,31,10,31,13,31,140,31,188,31,231,31,86,31,190,31,121,31,54,31,134,31,255,31,48,31,140,31,6,31,36,31,204,31,49,31,246,31,231,31,127,31,186,31,96,31,7,31,81,31,81,30,246,31,246,30,246,29,85,31,85,30,131,31,131,30,131,29,109,31,166,31,193,31,10,31,64,31,80,31,252,31,71,31,225,31,54,31,165,31,165,30,67,31,153,31,31,31,216,31,106,31,60,31,177,31,77,31,214,31,126,31,111,31,203,31,71,31,73,31,193,31,52,31,218,31,160,31,160,30,228,31,167,31,113,31,158,31,11,31,14,31,14,30,94,31,117,31,127,31,54,31,54,30,38,31,34,31,221,31,20,31,202,31,29,31,10,31,187,31,105,31,51,31,65,31,241,31,91,31,62,31,191,31,240,31,240,30,245,31,238,31,204,31,120,31,120,30,145,31,171,31,209,31,19,31,70,31,87,31,212,31,8,31,8,30,221,31,156,31,69,31,69,30,69,29,33,31,146,31,200,31,39,31,85,31,197,31,172,31,186,31,117,31,186,31,50,31,94,31,94,30,67,31,119,31,5,31,165,31,250,31,250,30,235,31,183,31,25,31,24,31,24,30,118,31,15,31,216,31,216,30,68,31,61,31,231,31,44,31,219,31,60,31,52,31,52,30,190,31,230,31,153,31,153,30,165,31,105,31,28,31,98,31,98,30,196,31,183,31,201,31,167,31,224,31,172,31,172,30,219,31,213,31,158,31,248,31,132,31,132,30,57,31,246,31,71,31,161,31,121,31,121,30,56,31,107,31,107,30,65,31,131,31,79,31,79,30,16,31,100,31,22,31,141,31,101,31,232,31,199,31,156,31,238,31,61,31,235,31,235,30,225,31,225,30,225,29,7,31,15,31,58,31,37,31,97,31,188,31,164,31,244,31,205,31,108,31,35,31,210,31,210,30,210,29,128,31,99,31,99,30,66,31,66,30,207,31,26,31,123,31,175,31,209,31,24,31,175,31,175,30,218,31,218,30,155,31,245,31,216,31,109,31,209,31,97,31,88,31,252,31,252,30,179,31,242,31,10,31,160,31,160,30,38,31,242,31,88,31,223,31,155,31,56,31,112,31,112,30,112,29,129,31,129,30,129,29,141,31,252,31,252,30,109,31,221,31,43,31,148,31,206,31,174,31,71,31,81,31,119,31,119,30,73,31,164,31,216,31,128,31,207,31,228,31,173,31,121,31,108,31,43,31,53,31,251,31,25,31,92,31,207,31,174,31,210,31,28,31,28,30,191,31,191,30,162,31,114,31,106,31,106,30,40,31,109,31,29,31,114,31,114,30,18,31,103,31,228,31,228,30,193,31,193,30,89,31,102,31,118,31,179,31,50,31,254,31,192,31,28,31,206,31,78,31,117,31,192,31,64,31,64,30,64,29,21,31,51,31,51,30,49,31,88,31,199,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
