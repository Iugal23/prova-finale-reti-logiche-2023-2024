-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_98 is
end project_tb_98;

architecture project_tb_arch_98 of project_tb_98 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 243;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (240,0,0,0,144,0,119,0,238,0,180,0,205,0,76,0,226,0,111,0,0,0,0,0,158,0,236,0,73,0,247,0,0,0,196,0,179,0,0,0,100,0,35,0,154,0,0,0,65,0,10,0,107,0,14,0,244,0,32,0,132,0,208,0,192,0,122,0,0,0,149,0,0,0,143,0,232,0,226,0,0,0,43,0,145,0,141,0,23,0,44,0,0,0,58,0,156,0,220,0,0,0,0,0,210,0,0,0,11,0,213,0,106,0,225,0,0,0,18,0,0,0,118,0,0,0,134,0,16,0,0,0,120,0,174,0,166,0,0,0,227,0,129,0,0,0,157,0,62,0,32,0,22,0,0,0,88,0,88,0,118,0,185,0,241,0,0,0,0,0,96,0,0,0,196,0,174,0,31,0,51,0,233,0,119,0,5,0,119,0,114,0,0,0,0,0,191,0,230,0,2,0,0,0,0,0,214,0,49,0,0,0,10,0,127,0,209,0,213,0,191,0,186,0,39,0,233,0,216,0,0,0,85,0,189,0,146,0,184,0,142,0,76,0,58,0,50,0,108,0,98,0,137,0,23,0,193,0,152,0,19,0,35,0,21,0,131,0,47,0,2,0,64,0,175,0,16,0,37,0,224,0,83,0,23,0,0,0,0,0,8,0,189,0,25,0,0,0,158,0,0,0,97,0,239,0,62,0,0,0,43,0,84,0,67,0,193,0,163,0,115,0,0,0,110,0,139,0,43,0,135,0,235,0,227,0,208,0,164,0,89,0,139,0,65,0,0,0,104,0,205,0,0,0,104,0,0,0,122,0,136,0,132,0,225,0,134,0,245,0,16,0,213,0,0,0,108,0,0,0,166,0,117,0,0,0,123,0,0,0,0,0,121,0,0,0,84,0,114,0,0,0,175,0,85,0,0,0,0,0,168,0,226,0,0,0,0,0,0,0,194,0,0,0,228,0,117,0,232,0,168,0,0,0,105,0,249,0,24,0,189,0,255,0,114,0,88,0,47,0,123,0,0,0,44,0,44,0,146,0,19,0,42,0,54,0,119,0,61,0,0,0,123,0,0,0,69,0,202,0,79,0,193,0,152,0);
signal scenario_full  : scenario_type := (240,31,240,30,144,31,119,31,238,31,180,31,205,31,76,31,226,31,111,31,111,30,111,29,158,31,236,31,73,31,247,31,247,30,196,31,179,31,179,30,100,31,35,31,154,31,154,30,65,31,10,31,107,31,14,31,244,31,32,31,132,31,208,31,192,31,122,31,122,30,149,31,149,30,143,31,232,31,226,31,226,30,43,31,145,31,141,31,23,31,44,31,44,30,58,31,156,31,220,31,220,30,220,29,210,31,210,30,11,31,213,31,106,31,225,31,225,30,18,31,18,30,118,31,118,30,134,31,16,31,16,30,120,31,174,31,166,31,166,30,227,31,129,31,129,30,157,31,62,31,32,31,22,31,22,30,88,31,88,31,118,31,185,31,241,31,241,30,241,29,96,31,96,30,196,31,174,31,31,31,51,31,233,31,119,31,5,31,119,31,114,31,114,30,114,29,191,31,230,31,2,31,2,30,2,29,214,31,49,31,49,30,10,31,127,31,209,31,213,31,191,31,186,31,39,31,233,31,216,31,216,30,85,31,189,31,146,31,184,31,142,31,76,31,58,31,50,31,108,31,98,31,137,31,23,31,193,31,152,31,19,31,35,31,21,31,131,31,47,31,2,31,64,31,175,31,16,31,37,31,224,31,83,31,23,31,23,30,23,29,8,31,189,31,25,31,25,30,158,31,158,30,97,31,239,31,62,31,62,30,43,31,84,31,67,31,193,31,163,31,115,31,115,30,110,31,139,31,43,31,135,31,235,31,227,31,208,31,164,31,89,31,139,31,65,31,65,30,104,31,205,31,205,30,104,31,104,30,122,31,136,31,132,31,225,31,134,31,245,31,16,31,213,31,213,30,108,31,108,30,166,31,117,31,117,30,123,31,123,30,123,29,121,31,121,30,84,31,114,31,114,30,175,31,85,31,85,30,85,29,168,31,226,31,226,30,226,29,226,28,194,31,194,30,228,31,117,31,232,31,168,31,168,30,105,31,249,31,24,31,189,31,255,31,114,31,88,31,47,31,123,31,123,30,44,31,44,31,146,31,19,31,42,31,54,31,119,31,61,31,61,30,123,31,123,30,69,31,202,31,79,31,193,31,152,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
