-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_899 is
end project_tb_899;

architecture project_tb_arch_899 of project_tb_899 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 789;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (24,0,127,0,0,0,195,0,27,0,217,0,96,0,64,0,68,0,93,0,120,0,208,0,150,0,142,0,121,0,0,0,0,0,185,0,233,0,252,0,22,0,154,0,23,0,91,0,188,0,0,0,0,0,0,0,194,0,58,0,0,0,56,0,49,0,111,0,65,0,15,0,0,0,0,0,136,0,162,0,97,0,218,0,199,0,184,0,4,0,73,0,73,0,13,0,106,0,75,0,43,0,218,0,0,0,113,0,6,0,231,0,0,0,192,0,81,0,162,0,53,0,195,0,102,0,218,0,0,0,0,0,213,0,0,0,228,0,252,0,217,0,21,0,107,0,25,0,0,0,135,0,110,0,87,0,211,0,0,0,246,0,166,0,50,0,3,0,133,0,34,0,172,0,37,0,155,0,121,0,139,0,78,0,8,0,124,0,128,0,175,0,0,0,0,0,177,0,60,0,202,0,177,0,31,0,219,0,169,0,46,0,109,0,200,0,208,0,0,0,0,0,72,0,7,0,212,0,61,0,139,0,227,0,154,0,99,0,55,0,0,0,77,0,38,0,116,0,164,0,229,0,209,0,169,0,15,0,33,0,198,0,57,0,120,0,140,0,75,0,247,0,242,0,220,0,82,0,134,0,48,0,226,0,176,0,87,0,242,0,189,0,70,0,122,0,0,0,163,0,43,0,0,0,236,0,151,0,48,0,204,0,0,0,228,0,171,0,115,0,12,0,38,0,13,0,92,0,236,0,229,0,154,0,77,0,0,0,199,0,128,0,233,0,142,0,190,0,0,0,65,0,157,0,53,0,0,0,226,0,0,0,234,0,82,0,244,0,201,0,46,0,104,0,232,0,207,0,53,0,209,0,0,0,69,0,189,0,241,0,116,0,222,0,213,0,4,0,185,0,156,0,65,0,183,0,95,0,91,0,117,0,0,0,157,0,0,0,18,0,108,0,34,0,67,0,18,0,159,0,40,0,138,0,76,0,36,0,113,0,0,0,174,0,47,0,0,0,37,0,92,0,124,0,137,0,0,0,0,0,52,0,0,0,65,0,142,0,183,0,69,0,0,0,61,0,203,0,91,0,80,0,0,0,236,0,38,0,85,0,21,0,158,0,0,0,186,0,154,0,0,0,174,0,0,0,83,0,114,0,1,0,166,0,210,0,27,0,144,0,166,0,135,0,0,0,119,0,226,0,0,0,140,0,0,0,61,0,173,0,15,0,17,0,252,0,185,0,245,0,173,0,225,0,54,0,46,0,16,0,25,0,59,0,221,0,86,0,112,0,114,0,91,0,29,0,131,0,133,0,68,0,168,0,102,0,105,0,235,0,243,0,171,0,108,0,0,0,29,0,146,0,0,0,212,0,42,0,148,0,0,0,0,0,234,0,0,0,189,0,49,0,0,0,166,0,15,0,119,0,0,0,187,0,73,0,112,0,122,0,146,0,105,0,92,0,0,0,0,0,0,0,88,0,13,0,246,0,0,0,198,0,210,0,0,0,82,0,207,0,0,0,228,0,223,0,1,0,0,0,192,0,101,0,0,0,50,0,0,0,108,0,0,0,5,0,83,0,0,0,33,0,43,0,144,0,0,0,67,0,61,0,110,0,143,0,0,0,0,0,55,0,165,0,2,0,89,0,118,0,113,0,193,0,0,0,0,0,204,0,175,0,234,0,147,0,121,0,225,0,104,0,216,0,7,0,73,0,79,0,240,0,79,0,48,0,68,0,114,0,252,0,123,0,39,0,116,0,0,0,0,0,174,0,72,0,0,0,147,0,0,0,0,0,98,0,0,0,173,0,202,0,0,0,32,0,56,0,234,0,154,0,16,0,218,0,225,0,0,0,22,0,38,0,116,0,100,0,0,0,244,0,204,0,0,0,0,0,0,0,191,0,117,0,137,0,194,0,86,0,54,0,0,0,148,0,64,0,80,0,252,0,94,0,126,0,18,0,59,0,139,0,0,0,84,0,186,0,0,0,126,0,118,0,0,0,121,0,129,0,118,0,0,0,86,0,43,0,78,0,227,0,55,0,152,0,126,0,176,0,216,0,56,0,0,0,54,0,127,0,179,0,241,0,134,0,70,0,124,0,36,0,160,0,15,0,173,0,112,0,76,0,218,0,0,0,0,0,9,0,252,0,0,0,101,0,33,0,171,0,140,0,230,0,251,0,23,0,0,0,189,0,78,0,225,0,219,0,201,0,119,0,0,0,108,0,48,0,0,0,69,0,0,0,193,0,119,0,0,0,119,0,45,0,235,0,6,0,195,0,32,0,65,0,0,0,0,0,238,0,206,0,0,0,225,0,0,0,106,0,103,0,0,0,0,0,163,0,185,0,0,0,108,0,47,0,118,0,0,0,0,0,72,0,129,0,0,0,195,0,153,0,49,0,0,0,115,0,158,0,154,0,2,0,231,0,25,0,1,0,9,0,0,0,31,0,0,0,247,0,0,0,191,0,23,0,37,0,39,0,132,0,47,0,0,0,48,0,13,0,41,0,155,0,57,0,207,0,125,0,162,0,50,0,0,0,0,0,0,0,244,0,61,0,5,0,0,0,228,0,81,0,0,0,228,0,75,0,94,0,64,0,185,0,249,0,136,0,78,0,72,0,91,0,0,0,90,0,78,0,0,0,23,0,103,0,130,0,125,0,171,0,37,0,39,0,191,0,123,0,81,0,123,0,25,0,238,0,114,0,202,0,217,0,253,0,164,0,120,0,251,0,186,0,115,0,45,0,0,0,0,0,132,0,7,0,4,0,211,0,244,0,206,0,247,0,128,0,80,0,1,0,0,0,187,0,223,0,12,0,141,0,158,0,169,0,186,0,0,0,110,0,134,0,144,0,8,0,0,0,195,0,0,0,0,0,0,0,17,0,0,0,19,0,141,0,87,0,185,0,39,0,29,0,212,0,16,0,163,0,182,0,177,0,116,0,156,0,166,0,144,0,0,0,0,0,192,0,101,0,154,0,0,0,230,0,169,0,46,0,131,0,229,0,0,0,105,0,104,0,0,0,250,0,174,0,30,0,85,0,12,0,0,0,46,0,0,0,26,0,20,0,121,0,166,0,180,0,0,0,88,0,165,0,89,0,74,0,129,0,234,0,31,0,238,0,133,0,196,0,0,0,89,0,0,0,234,0,251,0,145,0,207,0,13,0,0,0,0,0,106,0,165,0,0,0,250,0,224,0,0,0,195,0,120,0,210,0,157,0,125,0,31,0,119,0,135,0,170,0,156,0,56,0,107,0,0,0,61,0,101,0,158,0,71,0,121,0,68,0,182,0,177,0,132,0,222,0,91,0,0,0,7,0,0,0,242,0,64,0,200,0,207,0,241,0,242,0,242,0,21,0,79,0,65,0,150,0,0,0,97,0,0,0,0,0,0,0,120,0,174,0,173,0,50,0,254,0,34,0,79,0,180,0,116,0,24,0,0,0,128,0,0,0,43,0,183,0,132,0,0,0,0,0,9,0,30,0,242,0,72,0,149,0,233,0,3,0,92,0,254,0,162,0,45,0,177,0,14,0,0,0,0,0,177,0,200,0);
signal scenario_full  : scenario_type := (24,31,127,31,127,30,195,31,27,31,217,31,96,31,64,31,68,31,93,31,120,31,208,31,150,31,142,31,121,31,121,30,121,29,185,31,233,31,252,31,22,31,154,31,23,31,91,31,188,31,188,30,188,29,188,28,194,31,58,31,58,30,56,31,49,31,111,31,65,31,15,31,15,30,15,29,136,31,162,31,97,31,218,31,199,31,184,31,4,31,73,31,73,31,13,31,106,31,75,31,43,31,218,31,218,30,113,31,6,31,231,31,231,30,192,31,81,31,162,31,53,31,195,31,102,31,218,31,218,30,218,29,213,31,213,30,228,31,252,31,217,31,21,31,107,31,25,31,25,30,135,31,110,31,87,31,211,31,211,30,246,31,166,31,50,31,3,31,133,31,34,31,172,31,37,31,155,31,121,31,139,31,78,31,8,31,124,31,128,31,175,31,175,30,175,29,177,31,60,31,202,31,177,31,31,31,219,31,169,31,46,31,109,31,200,31,208,31,208,30,208,29,72,31,7,31,212,31,61,31,139,31,227,31,154,31,99,31,55,31,55,30,77,31,38,31,116,31,164,31,229,31,209,31,169,31,15,31,33,31,198,31,57,31,120,31,140,31,75,31,247,31,242,31,220,31,82,31,134,31,48,31,226,31,176,31,87,31,242,31,189,31,70,31,122,31,122,30,163,31,43,31,43,30,236,31,151,31,48,31,204,31,204,30,228,31,171,31,115,31,12,31,38,31,13,31,92,31,236,31,229,31,154,31,77,31,77,30,199,31,128,31,233,31,142,31,190,31,190,30,65,31,157,31,53,31,53,30,226,31,226,30,234,31,82,31,244,31,201,31,46,31,104,31,232,31,207,31,53,31,209,31,209,30,69,31,189,31,241,31,116,31,222,31,213,31,4,31,185,31,156,31,65,31,183,31,95,31,91,31,117,31,117,30,157,31,157,30,18,31,108,31,34,31,67,31,18,31,159,31,40,31,138,31,76,31,36,31,113,31,113,30,174,31,47,31,47,30,37,31,92,31,124,31,137,31,137,30,137,29,52,31,52,30,65,31,142,31,183,31,69,31,69,30,61,31,203,31,91,31,80,31,80,30,236,31,38,31,85,31,21,31,158,31,158,30,186,31,154,31,154,30,174,31,174,30,83,31,114,31,1,31,166,31,210,31,27,31,144,31,166,31,135,31,135,30,119,31,226,31,226,30,140,31,140,30,61,31,173,31,15,31,17,31,252,31,185,31,245,31,173,31,225,31,54,31,46,31,16,31,25,31,59,31,221,31,86,31,112,31,114,31,91,31,29,31,131,31,133,31,68,31,168,31,102,31,105,31,235,31,243,31,171,31,108,31,108,30,29,31,146,31,146,30,212,31,42,31,148,31,148,30,148,29,234,31,234,30,189,31,49,31,49,30,166,31,15,31,119,31,119,30,187,31,73,31,112,31,122,31,146,31,105,31,92,31,92,30,92,29,92,28,88,31,13,31,246,31,246,30,198,31,210,31,210,30,82,31,207,31,207,30,228,31,223,31,1,31,1,30,192,31,101,31,101,30,50,31,50,30,108,31,108,30,5,31,83,31,83,30,33,31,43,31,144,31,144,30,67,31,61,31,110,31,143,31,143,30,143,29,55,31,165,31,2,31,89,31,118,31,113,31,193,31,193,30,193,29,204,31,175,31,234,31,147,31,121,31,225,31,104,31,216,31,7,31,73,31,79,31,240,31,79,31,48,31,68,31,114,31,252,31,123,31,39,31,116,31,116,30,116,29,174,31,72,31,72,30,147,31,147,30,147,29,98,31,98,30,173,31,202,31,202,30,32,31,56,31,234,31,154,31,16,31,218,31,225,31,225,30,22,31,38,31,116,31,100,31,100,30,244,31,204,31,204,30,204,29,204,28,191,31,117,31,137,31,194,31,86,31,54,31,54,30,148,31,64,31,80,31,252,31,94,31,126,31,18,31,59,31,139,31,139,30,84,31,186,31,186,30,126,31,118,31,118,30,121,31,129,31,118,31,118,30,86,31,43,31,78,31,227,31,55,31,152,31,126,31,176,31,216,31,56,31,56,30,54,31,127,31,179,31,241,31,134,31,70,31,124,31,36,31,160,31,15,31,173,31,112,31,76,31,218,31,218,30,218,29,9,31,252,31,252,30,101,31,33,31,171,31,140,31,230,31,251,31,23,31,23,30,189,31,78,31,225,31,219,31,201,31,119,31,119,30,108,31,48,31,48,30,69,31,69,30,193,31,119,31,119,30,119,31,45,31,235,31,6,31,195,31,32,31,65,31,65,30,65,29,238,31,206,31,206,30,225,31,225,30,106,31,103,31,103,30,103,29,163,31,185,31,185,30,108,31,47,31,118,31,118,30,118,29,72,31,129,31,129,30,195,31,153,31,49,31,49,30,115,31,158,31,154,31,2,31,231,31,25,31,1,31,9,31,9,30,31,31,31,30,247,31,247,30,191,31,23,31,37,31,39,31,132,31,47,31,47,30,48,31,13,31,41,31,155,31,57,31,207,31,125,31,162,31,50,31,50,30,50,29,50,28,244,31,61,31,5,31,5,30,228,31,81,31,81,30,228,31,75,31,94,31,64,31,185,31,249,31,136,31,78,31,72,31,91,31,91,30,90,31,78,31,78,30,23,31,103,31,130,31,125,31,171,31,37,31,39,31,191,31,123,31,81,31,123,31,25,31,238,31,114,31,202,31,217,31,253,31,164,31,120,31,251,31,186,31,115,31,45,31,45,30,45,29,132,31,7,31,4,31,211,31,244,31,206,31,247,31,128,31,80,31,1,31,1,30,187,31,223,31,12,31,141,31,158,31,169,31,186,31,186,30,110,31,134,31,144,31,8,31,8,30,195,31,195,30,195,29,195,28,17,31,17,30,19,31,141,31,87,31,185,31,39,31,29,31,212,31,16,31,163,31,182,31,177,31,116,31,156,31,166,31,144,31,144,30,144,29,192,31,101,31,154,31,154,30,230,31,169,31,46,31,131,31,229,31,229,30,105,31,104,31,104,30,250,31,174,31,30,31,85,31,12,31,12,30,46,31,46,30,26,31,20,31,121,31,166,31,180,31,180,30,88,31,165,31,89,31,74,31,129,31,234,31,31,31,238,31,133,31,196,31,196,30,89,31,89,30,234,31,251,31,145,31,207,31,13,31,13,30,13,29,106,31,165,31,165,30,250,31,224,31,224,30,195,31,120,31,210,31,157,31,125,31,31,31,119,31,135,31,170,31,156,31,56,31,107,31,107,30,61,31,101,31,158,31,71,31,121,31,68,31,182,31,177,31,132,31,222,31,91,31,91,30,7,31,7,30,242,31,64,31,200,31,207,31,241,31,242,31,242,31,21,31,79,31,65,31,150,31,150,30,97,31,97,30,97,29,97,28,120,31,174,31,173,31,50,31,254,31,34,31,79,31,180,31,116,31,24,31,24,30,128,31,128,30,43,31,183,31,132,31,132,30,132,29,9,31,30,31,242,31,72,31,149,31,233,31,3,31,92,31,254,31,162,31,45,31,177,31,14,31,14,30,14,29,177,31,200,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
