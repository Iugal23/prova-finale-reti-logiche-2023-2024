-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 289;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (251,0,243,0,154,0,32,0,177,0,0,0,244,0,71,0,193,0,8,0,158,0,184,0,0,0,197,0,150,0,172,0,247,0,102,0,77,0,50,0,229,0,166,0,250,0,35,0,0,0,134,0,109,0,248,0,140,0,57,0,0,0,145,0,127,0,0,0,44,0,233,0,164,0,168,0,158,0,66,0,83,0,0,0,0,0,110,0,28,0,0,0,199,0,134,0,172,0,0,0,222,0,0,0,0,0,7,0,162,0,252,0,204,0,16,0,83,0,233,0,240,0,208,0,20,0,98,0,149,0,132,0,161,0,0,0,254,0,162,0,182,0,63,0,210,0,56,0,0,0,185,0,123,0,8,0,252,0,132,0,0,0,126,0,101,0,251,0,201,0,80,0,65,0,0,0,0,0,51,0,101,0,0,0,185,0,55,0,174,0,132,0,89,0,88,0,122,0,0,0,0,0,211,0,205,0,198,0,147,0,189,0,33,0,98,0,0,0,17,0,234,0,79,0,143,0,76,0,0,0,70,0,195,0,187,0,0,0,113,0,0,0,215,0,74,0,0,0,170,0,31,0,103,0,213,0,225,0,116,0,92,0,143,0,227,0,179,0,99,0,44,0,139,0,158,0,6,0,232,0,203,0,156,0,23,0,0,0,96,0,124,0,222,0,179,0,146,0,0,0,188,0,53,0,141,0,4,0,87,0,243,0,0,0,224,0,54,0,45,0,213,0,248,0,0,0,59,0,212,0,155,0,59,0,0,0,127,0,2,0,0,0,242,0,197,0,238,0,126,0,205,0,0,0,160,0,244,0,129,0,211,0,0,0,150,0,86,0,80,0,98,0,89,0,131,0,17,0,237,0,198,0,170,0,168,0,0,0,156,0,114,0,175,0,0,0,0,0,163,0,117,0,0,0,118,0,153,0,97,0,215,0,56,0,74,0,0,0,148,0,82,0,187,0,39,0,95,0,128,0,0,0,217,0,204,0,132,0,234,0,0,0,129,0,168,0,167,0,20,0,163,0,217,0,0,0,0,0,77,0,0,0,99,0,116,0,255,0,33,0,174,0,0,0,197,0,171,0,58,0,233,0,244,0,0,0,41,0,70,0,39,0,235,0,41,0,116,0,217,0,139,0,0,0,233,0,249,0,0,0,0,0,12,0,159,0,5,0,209,0,135,0,190,0,155,0,215,0,172,0,31,0,2,0,238,0,0,0,233,0,12,0,189,0,92,0,5,0,112,0,203,0,249,0,143,0,174,0,0,0,137,0,0,0,0,0,187,0,242,0,65,0,60,0,0,0,122,0);
signal scenario_full  : scenario_type := (251,31,243,31,154,31,32,31,177,31,177,30,244,31,71,31,193,31,8,31,158,31,184,31,184,30,197,31,150,31,172,31,247,31,102,31,77,31,50,31,229,31,166,31,250,31,35,31,35,30,134,31,109,31,248,31,140,31,57,31,57,30,145,31,127,31,127,30,44,31,233,31,164,31,168,31,158,31,66,31,83,31,83,30,83,29,110,31,28,31,28,30,199,31,134,31,172,31,172,30,222,31,222,30,222,29,7,31,162,31,252,31,204,31,16,31,83,31,233,31,240,31,208,31,20,31,98,31,149,31,132,31,161,31,161,30,254,31,162,31,182,31,63,31,210,31,56,31,56,30,185,31,123,31,8,31,252,31,132,31,132,30,126,31,101,31,251,31,201,31,80,31,65,31,65,30,65,29,51,31,101,31,101,30,185,31,55,31,174,31,132,31,89,31,88,31,122,31,122,30,122,29,211,31,205,31,198,31,147,31,189,31,33,31,98,31,98,30,17,31,234,31,79,31,143,31,76,31,76,30,70,31,195,31,187,31,187,30,113,31,113,30,215,31,74,31,74,30,170,31,31,31,103,31,213,31,225,31,116,31,92,31,143,31,227,31,179,31,99,31,44,31,139,31,158,31,6,31,232,31,203,31,156,31,23,31,23,30,96,31,124,31,222,31,179,31,146,31,146,30,188,31,53,31,141,31,4,31,87,31,243,31,243,30,224,31,54,31,45,31,213,31,248,31,248,30,59,31,212,31,155,31,59,31,59,30,127,31,2,31,2,30,242,31,197,31,238,31,126,31,205,31,205,30,160,31,244,31,129,31,211,31,211,30,150,31,86,31,80,31,98,31,89,31,131,31,17,31,237,31,198,31,170,31,168,31,168,30,156,31,114,31,175,31,175,30,175,29,163,31,117,31,117,30,118,31,153,31,97,31,215,31,56,31,74,31,74,30,148,31,82,31,187,31,39,31,95,31,128,31,128,30,217,31,204,31,132,31,234,31,234,30,129,31,168,31,167,31,20,31,163,31,217,31,217,30,217,29,77,31,77,30,99,31,116,31,255,31,33,31,174,31,174,30,197,31,171,31,58,31,233,31,244,31,244,30,41,31,70,31,39,31,235,31,41,31,116,31,217,31,139,31,139,30,233,31,249,31,249,30,249,29,12,31,159,31,5,31,209,31,135,31,190,31,155,31,215,31,172,31,31,31,2,31,238,31,238,30,233,31,12,31,189,31,92,31,5,31,112,31,203,31,249,31,143,31,174,31,174,30,137,31,137,30,137,29,187,31,242,31,65,31,60,31,60,30,122,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
