-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_447 is
end project_tb_447;

architecture project_tb_arch_447 of project_tb_447 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 500;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (68,0,33,0,255,0,62,0,163,0,0,0,64,0,6,0,245,0,31,0,50,0,84,0,215,0,245,0,78,0,249,0,0,0,2,0,162,0,74,0,122,0,122,0,143,0,94,0,219,0,3,0,29,0,210,0,188,0,0,0,216,0,162,0,184,0,118,0,85,0,199,0,132,0,0,0,120,0,141,0,0,0,6,0,36,0,102,0,127,0,153,0,0,0,11,0,226,0,0,0,0,0,0,0,0,0,193,0,99,0,174,0,244,0,111,0,0,0,197,0,179,0,79,0,0,0,32,0,34,0,0,0,54,0,180,0,112,0,161,0,202,0,0,0,0,0,30,0,46,0,245,0,162,0,29,0,51,0,0,0,201,0,0,0,243,0,116,0,102,0,195,0,16,0,122,0,0,0,25,0,132,0,0,0,57,0,71,0,38,0,76,0,181,0,208,0,184,0,191,0,0,0,0,0,70,0,243,0,23,0,175,0,0,0,2,0,102,0,0,0,238,0,91,0,0,0,0,0,100,0,196,0,161,0,102,0,194,0,172,0,60,0,198,0,122,0,0,0,176,0,0,0,72,0,248,0,219,0,207,0,19,0,31,0,117,0,30,0,196,0,99,0,206,0,116,0,42,0,254,0,9,0,193,0,236,0,210,0,39,0,183,0,193,0,202,0,105,0,241,0,174,0,150,0,161,0,183,0,36,0,143,0,0,0,18,0,0,0,225,0,185,0,37,0,0,0,33,0,111,0,204,0,115,0,249,0,216,0,145,0,94,0,0,0,124,0,63,0,0,0,6,0,29,0,0,0,217,0,180,0,0,0,156,0,164,0,207,0,0,0,135,0,56,0,119,0,68,0,42,0,148,0,0,0,227,0,34,0,190,0,90,0,77,0,110,0,0,0,253,0,85,0,7,0,238,0,170,0,0,0,72,0,145,0,100,0,0,0,93,0,5,0,194,0,162,0,0,0,90,0,177,0,244,0,169,0,169,0,201,0,204,0,0,0,213,0,0,0,235,0,145,0,54,0,0,0,23,0,95,0,0,0,0,0,244,0,174,0,38,0,247,0,0,0,216,0,123,0,196,0,24,0,8,0,25,0,97,0,0,0,131,0,75,0,51,0,0,0,56,0,133,0,0,0,17,0,146,0,215,0,0,0,1,0,127,0,72,0,99,0,238,0,0,0,0,0,232,0,109,0,223,0,100,0,23,0,59,0,169,0,50,0,123,0,166,0,56,0,22,0,255,0,159,0,72,0,0,0,130,0,207,0,93,0,253,0,65,0,211,0,200,0,198,0,0,0,0,0,160,0,0,0,7,0,48,0,0,0,190,0,138,0,184,0,171,0,107,0,231,0,234,0,126,0,189,0,80,0,10,0,215,0,117,0,94,0,181,0,0,0,0,0,15,0,0,0,34,0,0,0,55,0,33,0,0,0,84,0,155,0,91,0,185,0,12,0,0,0,8,0,124,0,83,0,122,0,185,0,80,0,105,0,116,0,68,0,29,0,160,0,130,0,171,0,123,0,0,0,205,0,0,0,152,0,221,0,240,0,75,0,170,0,118,0,0,0,109,0,0,0,62,0,122,0,184,0,253,0,214,0,0,0,84,0,77,0,57,0,86,0,203,0,199,0,0,0,0,0,235,0,213,0,0,0,199,0,71,0,166,0,107,0,122,0,0,0,73,0,160,0,0,0,214,0,100,0,162,0,103,0,3,0,21,0,0,0,86,0,0,0,214,0,206,0,84,0,246,0,105,0,70,0,180,0,0,0,185,0,170,0,156,0,255,0,75,0,243,0,121,0,224,0,51,0,161,0,190,0,250,0,53,0,116,0,162,0,75,0,0,0,25,0,134,0,219,0,255,0,247,0,245,0,40,0,0,0,0,0,195,0,20,0,222,0,32,0,0,0,0,0,103,0,164,0,0,0,40,0,229,0,243,0,0,0,65,0,173,0,81,0,0,0,245,0,89,0,0,0,223,0,132,0,218,0,78,0,148,0,198,0,58,0,50,0,165,0,62,0,59,0,0,0,58,0,234,0,0,0,31,0,188,0,191,0,0,0,0,0,42,0,170,0,60,0,105,0,229,0,0,0,232,0,194,0,207,0,0,0,122,0,6,0,241,0,254,0,0,0,91,0,150,0,75,0,232,0,0,0,37,0,16,0,129,0,0,0,0,0,229,0,0,0,165,0,209,0,84,0,149,0,177,0,240,0,1,0,184,0,0,0,35,0,204,0,244,0,0,0,0,0);
signal scenario_full  : scenario_type := (68,31,33,31,255,31,62,31,163,31,163,30,64,31,6,31,245,31,31,31,50,31,84,31,215,31,245,31,78,31,249,31,249,30,2,31,162,31,74,31,122,31,122,31,143,31,94,31,219,31,3,31,29,31,210,31,188,31,188,30,216,31,162,31,184,31,118,31,85,31,199,31,132,31,132,30,120,31,141,31,141,30,6,31,36,31,102,31,127,31,153,31,153,30,11,31,226,31,226,30,226,29,226,28,226,27,193,31,99,31,174,31,244,31,111,31,111,30,197,31,179,31,79,31,79,30,32,31,34,31,34,30,54,31,180,31,112,31,161,31,202,31,202,30,202,29,30,31,46,31,245,31,162,31,29,31,51,31,51,30,201,31,201,30,243,31,116,31,102,31,195,31,16,31,122,31,122,30,25,31,132,31,132,30,57,31,71,31,38,31,76,31,181,31,208,31,184,31,191,31,191,30,191,29,70,31,243,31,23,31,175,31,175,30,2,31,102,31,102,30,238,31,91,31,91,30,91,29,100,31,196,31,161,31,102,31,194,31,172,31,60,31,198,31,122,31,122,30,176,31,176,30,72,31,248,31,219,31,207,31,19,31,31,31,117,31,30,31,196,31,99,31,206,31,116,31,42,31,254,31,9,31,193,31,236,31,210,31,39,31,183,31,193,31,202,31,105,31,241,31,174,31,150,31,161,31,183,31,36,31,143,31,143,30,18,31,18,30,225,31,185,31,37,31,37,30,33,31,111,31,204,31,115,31,249,31,216,31,145,31,94,31,94,30,124,31,63,31,63,30,6,31,29,31,29,30,217,31,180,31,180,30,156,31,164,31,207,31,207,30,135,31,56,31,119,31,68,31,42,31,148,31,148,30,227,31,34,31,190,31,90,31,77,31,110,31,110,30,253,31,85,31,7,31,238,31,170,31,170,30,72,31,145,31,100,31,100,30,93,31,5,31,194,31,162,31,162,30,90,31,177,31,244,31,169,31,169,31,201,31,204,31,204,30,213,31,213,30,235,31,145,31,54,31,54,30,23,31,95,31,95,30,95,29,244,31,174,31,38,31,247,31,247,30,216,31,123,31,196,31,24,31,8,31,25,31,97,31,97,30,131,31,75,31,51,31,51,30,56,31,133,31,133,30,17,31,146,31,215,31,215,30,1,31,127,31,72,31,99,31,238,31,238,30,238,29,232,31,109,31,223,31,100,31,23,31,59,31,169,31,50,31,123,31,166,31,56,31,22,31,255,31,159,31,72,31,72,30,130,31,207,31,93,31,253,31,65,31,211,31,200,31,198,31,198,30,198,29,160,31,160,30,7,31,48,31,48,30,190,31,138,31,184,31,171,31,107,31,231,31,234,31,126,31,189,31,80,31,10,31,215,31,117,31,94,31,181,31,181,30,181,29,15,31,15,30,34,31,34,30,55,31,33,31,33,30,84,31,155,31,91,31,185,31,12,31,12,30,8,31,124,31,83,31,122,31,185,31,80,31,105,31,116,31,68,31,29,31,160,31,130,31,171,31,123,31,123,30,205,31,205,30,152,31,221,31,240,31,75,31,170,31,118,31,118,30,109,31,109,30,62,31,122,31,184,31,253,31,214,31,214,30,84,31,77,31,57,31,86,31,203,31,199,31,199,30,199,29,235,31,213,31,213,30,199,31,71,31,166,31,107,31,122,31,122,30,73,31,160,31,160,30,214,31,100,31,162,31,103,31,3,31,21,31,21,30,86,31,86,30,214,31,206,31,84,31,246,31,105,31,70,31,180,31,180,30,185,31,170,31,156,31,255,31,75,31,243,31,121,31,224,31,51,31,161,31,190,31,250,31,53,31,116,31,162,31,75,31,75,30,25,31,134,31,219,31,255,31,247,31,245,31,40,31,40,30,40,29,195,31,20,31,222,31,32,31,32,30,32,29,103,31,164,31,164,30,40,31,229,31,243,31,243,30,65,31,173,31,81,31,81,30,245,31,89,31,89,30,223,31,132,31,218,31,78,31,148,31,198,31,58,31,50,31,165,31,62,31,59,31,59,30,58,31,234,31,234,30,31,31,188,31,191,31,191,30,191,29,42,31,170,31,60,31,105,31,229,31,229,30,232,31,194,31,207,31,207,30,122,31,6,31,241,31,254,31,254,30,91,31,150,31,75,31,232,31,232,30,37,31,16,31,129,31,129,30,129,29,229,31,229,30,165,31,209,31,84,31,149,31,177,31,240,31,1,31,184,31,184,30,35,31,204,31,244,31,244,30,244,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
