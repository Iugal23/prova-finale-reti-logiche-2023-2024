-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 175;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (154,0,0,0,123,0,89,0,50,0,255,0,0,0,36,0,243,0,214,0,149,0,110,0,62,0,63,0,184,0,16,0,18,0,93,0,0,0,115,0,148,0,82,0,251,0,224,0,245,0,26,0,28,0,0,0,0,0,252,0,168,0,209,0,225,0,0,0,64,0,22,0,31,0,209,0,192,0,0,0,129,0,121,0,178,0,82,0,0,0,4,0,0,0,191,0,55,0,178,0,0,0,181,0,83,0,59,0,0,0,81,0,255,0,249,0,0,0,0,0,118,0,179,0,100,0,83,0,90,0,186,0,213,0,85,0,33,0,129,0,151,0,22,0,47,0,131,0,232,0,187,0,214,0,0,0,153,0,0,0,0,0,209,0,212,0,54,0,174,0,11,0,185,0,194,0,0,0,79,0,48,0,0,0,1,0,25,0,173,0,59,0,0,0,79,0,84,0,78,0,78,0,195,0,0,0,222,0,8,0,100,0,15,0,0,0,146,0,150,0,97,0,73,0,0,0,8,0,111,0,163,0,77,0,42,0,84,0,173,0,240,0,45,0,136,0,187,0,198,0,202,0,22,0,81,0,157,0,154,0,247,0,206,0,212,0,255,0,24,0,122,0,226,0,53,0,98,0,171,0,154,0,153,0,143,0,6,0,204,0,79,0,4,0,221,0,13,0,145,0,44,0,173,0,40,0,161,0,16,0,172,0,115,0,195,0,29,0,48,0,208,0,53,0,132,0,0,0,0,0,17,0,59,0,0,0,141,0,142,0,0,0,46,0,197,0,43,0,219,0);
signal scenario_full  : scenario_type := (154,31,154,30,123,31,89,31,50,31,255,31,255,30,36,31,243,31,214,31,149,31,110,31,62,31,63,31,184,31,16,31,18,31,93,31,93,30,115,31,148,31,82,31,251,31,224,31,245,31,26,31,28,31,28,30,28,29,252,31,168,31,209,31,225,31,225,30,64,31,22,31,31,31,209,31,192,31,192,30,129,31,121,31,178,31,82,31,82,30,4,31,4,30,191,31,55,31,178,31,178,30,181,31,83,31,59,31,59,30,81,31,255,31,249,31,249,30,249,29,118,31,179,31,100,31,83,31,90,31,186,31,213,31,85,31,33,31,129,31,151,31,22,31,47,31,131,31,232,31,187,31,214,31,214,30,153,31,153,30,153,29,209,31,212,31,54,31,174,31,11,31,185,31,194,31,194,30,79,31,48,31,48,30,1,31,25,31,173,31,59,31,59,30,79,31,84,31,78,31,78,31,195,31,195,30,222,31,8,31,100,31,15,31,15,30,146,31,150,31,97,31,73,31,73,30,8,31,111,31,163,31,77,31,42,31,84,31,173,31,240,31,45,31,136,31,187,31,198,31,202,31,22,31,81,31,157,31,154,31,247,31,206,31,212,31,255,31,24,31,122,31,226,31,53,31,98,31,171,31,154,31,153,31,143,31,6,31,204,31,79,31,4,31,221,31,13,31,145,31,44,31,173,31,40,31,161,31,16,31,172,31,115,31,195,31,29,31,48,31,208,31,53,31,132,31,132,30,132,29,17,31,59,31,59,30,141,31,142,31,142,30,46,31,197,31,43,31,219,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
