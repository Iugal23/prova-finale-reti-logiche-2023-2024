-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 258;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (39,0,98,0,5,0,214,0,189,0,82,0,0,0,2,0,0,0,207,0,90,0,85,0,0,0,138,0,151,0,0,0,76,0,0,0,26,0,32,0,209,0,93,0,37,0,239,0,0,0,17,0,13,0,132,0,20,0,21,0,109,0,0,0,112,0,153,0,188,0,197,0,26,0,37,0,0,0,114,0,147,0,140,0,0,0,164,0,97,0,0,0,62,0,79,0,235,0,52,0,124,0,153,0,0,0,178,0,49,0,77,0,150,0,13,0,0,0,28,0,11,0,130,0,0,0,4,0,232,0,0,0,0,0,35,0,243,0,0,0,134,0,75,0,155,0,176,0,213,0,0,0,0,0,4,0,185,0,180,0,0,0,214,0,205,0,0,0,4,0,178,0,189,0,219,0,236,0,49,0,195,0,48,0,0,0,18,0,160,0,0,0,104,0,10,0,178,0,82,0,86,0,246,0,147,0,4,0,0,0,0,0,239,0,50,0,7,0,42,0,245,0,0,0,106,0,0,0,55,0,78,0,67,0,25,0,112,0,242,0,195,0,27,0,1,0,164,0,0,0,70,0,183,0,167,0,171,0,75,0,207,0,127,0,214,0,51,0,26,0,53,0,26,0,149,0,0,0,127,0,156,0,45,0,2,0,94,0,0,0,0,0,129,0,153,0,0,0,32,0,100,0,174,0,0,0,140,0,113,0,0,0,133,0,131,0,160,0,13,0,232,0,193,0,37,0,0,0,251,0,44,0,24,0,29,0,99,0,93,0,161,0,196,0,0,0,0,0,90,0,66,0,56,0,97,0,45,0,0,0,102,0,171,0,110,0,199,0,200,0,42,0,173,0,0,0,0,0,18,0,170,0,66,0,0,0,0,0,203,0,101,0,0,0,9,0,22,0,64,0,44,0,65,0,104,0,245,0,0,0,0,0,95,0,88,0,0,0,64,0,199,0,223,0,184,0,0,0,103,0,108,0,153,0,86,0,132,0,0,0,40,0,0,0,252,0,21,0,72,0,252,0,246,0,141,0,157,0,36,0,230,0,237,0,127,0,0,0,161,0,161,0,13,0,159,0,200,0,123,0,168,0,193,0,0,0,227,0,233,0,126,0,27,0,22,0,42,0,9,0,54,0,101,0,30,0,211,0,190,0,236,0,121,0,232,0);
signal scenario_full  : scenario_type := (39,31,98,31,5,31,214,31,189,31,82,31,82,30,2,31,2,30,207,31,90,31,85,31,85,30,138,31,151,31,151,30,76,31,76,30,26,31,32,31,209,31,93,31,37,31,239,31,239,30,17,31,13,31,132,31,20,31,21,31,109,31,109,30,112,31,153,31,188,31,197,31,26,31,37,31,37,30,114,31,147,31,140,31,140,30,164,31,97,31,97,30,62,31,79,31,235,31,52,31,124,31,153,31,153,30,178,31,49,31,77,31,150,31,13,31,13,30,28,31,11,31,130,31,130,30,4,31,232,31,232,30,232,29,35,31,243,31,243,30,134,31,75,31,155,31,176,31,213,31,213,30,213,29,4,31,185,31,180,31,180,30,214,31,205,31,205,30,4,31,178,31,189,31,219,31,236,31,49,31,195,31,48,31,48,30,18,31,160,31,160,30,104,31,10,31,178,31,82,31,86,31,246,31,147,31,4,31,4,30,4,29,239,31,50,31,7,31,42,31,245,31,245,30,106,31,106,30,55,31,78,31,67,31,25,31,112,31,242,31,195,31,27,31,1,31,164,31,164,30,70,31,183,31,167,31,171,31,75,31,207,31,127,31,214,31,51,31,26,31,53,31,26,31,149,31,149,30,127,31,156,31,45,31,2,31,94,31,94,30,94,29,129,31,153,31,153,30,32,31,100,31,174,31,174,30,140,31,113,31,113,30,133,31,131,31,160,31,13,31,232,31,193,31,37,31,37,30,251,31,44,31,24,31,29,31,99,31,93,31,161,31,196,31,196,30,196,29,90,31,66,31,56,31,97,31,45,31,45,30,102,31,171,31,110,31,199,31,200,31,42,31,173,31,173,30,173,29,18,31,170,31,66,31,66,30,66,29,203,31,101,31,101,30,9,31,22,31,64,31,44,31,65,31,104,31,245,31,245,30,245,29,95,31,88,31,88,30,64,31,199,31,223,31,184,31,184,30,103,31,108,31,153,31,86,31,132,31,132,30,40,31,40,30,252,31,21,31,72,31,252,31,246,31,141,31,157,31,36,31,230,31,237,31,127,31,127,30,161,31,161,31,13,31,159,31,200,31,123,31,168,31,193,31,193,30,227,31,233,31,126,31,27,31,22,31,42,31,9,31,54,31,101,31,30,31,211,31,190,31,236,31,121,31,232,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
