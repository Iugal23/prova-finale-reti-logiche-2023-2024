-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 243;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (163,0,142,0,90,0,0,0,203,0,77,0,1,0,213,0,103,0,240,0,121,0,68,0,48,0,44,0,75,0,106,0,3,0,0,0,59,0,69,0,61,0,182,0,203,0,0,0,190,0,43,0,0,0,139,0,122,0,0,0,244,0,173,0,184,0,0,0,189,0,0,0,214,0,0,0,0,0,0,0,0,0,0,0,61,0,152,0,0,0,185,0,66,0,184,0,94,0,140,0,0,0,167,0,198,0,0,0,0,0,0,0,21,0,82,0,0,0,59,0,0,0,0,0,0,0,101,0,55,0,182,0,131,0,0,0,89,0,194,0,0,0,156,0,218,0,148,0,83,0,0,0,179,0,0,0,127,0,208,0,105,0,230,0,0,0,62,0,88,0,212,0,0,0,160,0,111,0,18,0,84,0,232,0,149,0,173,0,243,0,223,0,0,0,0,0,176,0,155,0,4,0,0,0,97,0,0,0,136,0,82,0,0,0,191,0,21,0,139,0,195,0,250,0,92,0,197,0,0,0,102,0,0,0,201,0,57,0,232,0,98,0,77,0,121,0,20,0,0,0,0,0,3,0,156,0,0,0,0,0,79,0,0,0,77,0,125,0,114,0,85,0,8,0,168,0,96,0,0,0,0,0,0,0,239,0,138,0,49,0,234,0,143,0,175,0,68,0,132,0,0,0,14,0,216,0,0,0,29,0,52,0,243,0,13,0,146,0,48,0,238,0,200,0,228,0,39,0,163,0,115,0,136,0,212,0,0,0,121,0,183,0,190,0,83,0,28,0,0,0,36,0,153,0,0,0,52,0,147,0,93,0,0,0,16,0,0,0,159,0,206,0,154,0,91,0,207,0,0,0,156,0,251,0,148,0,29,0,87,0,56,0,56,0,38,0,167,0,31,0,137,0,0,0,0,0,141,0,15,0,155,0,210,0,9,0,118,0,104,0,173,0,255,0,0,0,205,0,48,0,199,0,75,0,153,0,0,0,217,0,0,0,195,0,89,0,68,0,205,0,94,0,120,0,243,0,59,0,0,0,24,0,153,0,87,0,207,0,67,0,25,0,194,0,0,0,183,0,78,0,29,0,133,0,187,0);
signal scenario_full  : scenario_type := (163,31,142,31,90,31,90,30,203,31,77,31,1,31,213,31,103,31,240,31,121,31,68,31,48,31,44,31,75,31,106,31,3,31,3,30,59,31,69,31,61,31,182,31,203,31,203,30,190,31,43,31,43,30,139,31,122,31,122,30,244,31,173,31,184,31,184,30,189,31,189,30,214,31,214,30,214,29,214,28,214,27,214,26,61,31,152,31,152,30,185,31,66,31,184,31,94,31,140,31,140,30,167,31,198,31,198,30,198,29,198,28,21,31,82,31,82,30,59,31,59,30,59,29,59,28,101,31,55,31,182,31,131,31,131,30,89,31,194,31,194,30,156,31,218,31,148,31,83,31,83,30,179,31,179,30,127,31,208,31,105,31,230,31,230,30,62,31,88,31,212,31,212,30,160,31,111,31,18,31,84,31,232,31,149,31,173,31,243,31,223,31,223,30,223,29,176,31,155,31,4,31,4,30,97,31,97,30,136,31,82,31,82,30,191,31,21,31,139,31,195,31,250,31,92,31,197,31,197,30,102,31,102,30,201,31,57,31,232,31,98,31,77,31,121,31,20,31,20,30,20,29,3,31,156,31,156,30,156,29,79,31,79,30,77,31,125,31,114,31,85,31,8,31,168,31,96,31,96,30,96,29,96,28,239,31,138,31,49,31,234,31,143,31,175,31,68,31,132,31,132,30,14,31,216,31,216,30,29,31,52,31,243,31,13,31,146,31,48,31,238,31,200,31,228,31,39,31,163,31,115,31,136,31,212,31,212,30,121,31,183,31,190,31,83,31,28,31,28,30,36,31,153,31,153,30,52,31,147,31,93,31,93,30,16,31,16,30,159,31,206,31,154,31,91,31,207,31,207,30,156,31,251,31,148,31,29,31,87,31,56,31,56,31,38,31,167,31,31,31,137,31,137,30,137,29,141,31,15,31,155,31,210,31,9,31,118,31,104,31,173,31,255,31,255,30,205,31,48,31,199,31,75,31,153,31,153,30,217,31,217,30,195,31,89,31,68,31,205,31,94,31,120,31,243,31,59,31,59,30,24,31,153,31,87,31,207,31,67,31,25,31,194,31,194,30,183,31,78,31,29,31,133,31,187,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
