-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 568;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,17,0,182,0,236,0,140,0,0,0,0,0,146,0,63,0,18,0,0,0,215,0,173,0,0,0,43,0,48,0,0,0,36,0,48,0,120,0,0,0,39,0,0,0,164,0,5,0,190,0,242,0,0,0,229,0,46,0,108,0,174,0,64,0,124,0,90,0,0,0,203,0,92,0,0,0,120,0,71,0,0,0,242,0,0,0,115,0,111,0,66,0,219,0,111,0,174,0,0,0,144,0,22,0,245,0,48,0,213,0,8,0,78,0,155,0,106,0,0,0,0,0,248,0,0,0,112,0,149,0,23,0,82,0,50,0,4,0,224,0,59,0,61,0,149,0,16,0,113,0,205,0,158,0,32,0,154,0,0,0,66,0,115,0,24,0,176,0,0,0,36,0,69,0,0,0,205,0,209,0,248,0,51,0,0,0,165,0,249,0,66,0,136,0,133,0,208,0,0,0,255,0,114,0,128,0,221,0,209,0,233,0,0,0,0,0,42,0,126,0,23,0,0,0,190,0,120,0,7,0,35,0,0,0,181,0,0,0,51,0,114,0,235,0,0,0,13,0,109,0,208,0,210,0,0,0,125,0,154,0,206,0,0,0,237,0,0,0,125,0,50,0,206,0,0,0,200,0,48,0,210,0,111,0,0,0,251,0,240,0,0,0,0,0,161,0,147,0,18,0,0,0,254,0,239,0,203,0,80,0,0,0,215,0,129,0,65,0,45,0,80,0,92,0,134,0,153,0,99,0,189,0,102,0,175,0,66,0,184,0,249,0,30,0,26,0,0,0,201,0,150,0,0,0,99,0,152,0,0,0,115,0,129,0,54,0,18,0,125,0,35,0,0,0,0,0,236,0,0,0,25,0,238,0,66,0,0,0,102,0,159,0,0,0,110,0,0,0,118,0,0,0,0,0,165,0,14,0,239,0,198,0,103,0,11,0,0,0,0,0,248,0,0,0,0,0,51,0,0,0,65,0,110,0,213,0,28,0,135,0,100,0,36,0,241,0,0,0,203,0,51,0,135,0,0,0,0,0,198,0,24,0,22,0,30,0,104,0,135,0,0,0,68,0,106,0,9,0,181,0,223,0,192,0,90,0,66,0,253,0,185,0,0,0,0,0,196,0,31,0,74,0,122,0,193,0,110,0,217,0,0,0,6,0,236,0,62,0,0,0,182,0,2,0,0,0,0,0,240,0,53,0,192,0,0,0,118,0,142,0,4,0,0,0,244,0,12,0,68,0,44,0,238,0,21,0,0,0,186,0,106,0,153,0,30,0,57,0,0,0,152,0,245,0,196,0,174,0,112,0,249,0,150,0,0,0,220,0,10,0,4,0,80,0,180,0,128,0,68,0,31,0,232,0,172,0,255,0,10,0,19,0,144,0,102,0,195,0,218,0,194,0,108,0,198,0,43,0,10,0,0,0,195,0,66,0,0,0,207,0,94,0,0,0,0,0,145,0,97,0,154,0,96,0,97,0,241,0,177,0,240,0,0,0,50,0,180,0,92,0,5,0,169,0,18,0,107,0,209,0,247,0,151,0,98,0,190,0,82,0,103,0,0,0,0,0,0,0,0,0,0,0,154,0,71,0,0,0,96,0,11,0,163,0,166,0,0,0,127,0,169,0,0,0,41,0,0,0,0,0,0,0,0,0,41,0,249,0,137,0,121,0,135,0,0,0,246,0,0,0,190,0,0,0,0,0,0,0,182,0,144,0,0,0,129,0,0,0,181,0,40,0,100,0,243,0,0,0,0,0,235,0,116,0,243,0,194,0,114,0,212,0,0,0,119,0,198,0,110,0,66,0,159,0,61,0,225,0,0,0,85,0,0,0,4,0,157,0,78,0,5,0,53,0,0,0,0,0,0,0,224,0,149,0,125,0,46,0,58,0,242,0,0,0,120,0,0,0,93,0,167,0,38,0,51,0,0,0,0,0,0,0,0,0,0,0,44,0,140,0,232,0,115,0,0,0,0,0,0,0,203,0,237,0,0,0,65,0,242,0,126,0,92,0,0,0,27,0,159,0,234,0,53,0,227,0,120,0,166,0,143,0,94,0,204,0,18,0,0,0,82,0,72,0,144,0,174,0,187,0,75,0,246,0,117,0,42,0,93,0,0,0,146,0,74,0,119,0,211,0,75,0,0,0,0,0,0,0,99,0,79,0,56,0,0,0,45,0,71,0,173,0,121,0,208,0,0,0,190,0,33,0,0,0,77,0,193,0,37,0,138,0,203,0,18,0,158,0,0,0,28,0,0,0,81,0,102,0,0,0,132,0,106,0,0,0,4,0,77,0,163,0,205,0,85,0,149,0,188,0,243,0,165,0,0,0,0,0,24,0,16,0,10,0,110,0,94,0,68,0,0,0,0,0,0,0,162,0,240,0,38,0,25,0,156,0,0,0,88,0,67,0,246,0,245,0,0,0,0,0,133,0,251,0,158,0,144,0,64,0,30,0,176,0,207,0,200,0,66,0,201,0,5,0,0,0,61,0,241,0,149,0,209,0,0,0,169,0,211,0,123,0,184,0,46,0,144,0,141,0,132,0,198,0);
signal scenario_full  : scenario_type := (0,0,17,31,182,31,236,31,140,31,140,30,140,29,146,31,63,31,18,31,18,30,215,31,173,31,173,30,43,31,48,31,48,30,36,31,48,31,120,31,120,30,39,31,39,30,164,31,5,31,190,31,242,31,242,30,229,31,46,31,108,31,174,31,64,31,124,31,90,31,90,30,203,31,92,31,92,30,120,31,71,31,71,30,242,31,242,30,115,31,111,31,66,31,219,31,111,31,174,31,174,30,144,31,22,31,245,31,48,31,213,31,8,31,78,31,155,31,106,31,106,30,106,29,248,31,248,30,112,31,149,31,23,31,82,31,50,31,4,31,224,31,59,31,61,31,149,31,16,31,113,31,205,31,158,31,32,31,154,31,154,30,66,31,115,31,24,31,176,31,176,30,36,31,69,31,69,30,205,31,209,31,248,31,51,31,51,30,165,31,249,31,66,31,136,31,133,31,208,31,208,30,255,31,114,31,128,31,221,31,209,31,233,31,233,30,233,29,42,31,126,31,23,31,23,30,190,31,120,31,7,31,35,31,35,30,181,31,181,30,51,31,114,31,235,31,235,30,13,31,109,31,208,31,210,31,210,30,125,31,154,31,206,31,206,30,237,31,237,30,125,31,50,31,206,31,206,30,200,31,48,31,210,31,111,31,111,30,251,31,240,31,240,30,240,29,161,31,147,31,18,31,18,30,254,31,239,31,203,31,80,31,80,30,215,31,129,31,65,31,45,31,80,31,92,31,134,31,153,31,99,31,189,31,102,31,175,31,66,31,184,31,249,31,30,31,26,31,26,30,201,31,150,31,150,30,99,31,152,31,152,30,115,31,129,31,54,31,18,31,125,31,35,31,35,30,35,29,236,31,236,30,25,31,238,31,66,31,66,30,102,31,159,31,159,30,110,31,110,30,118,31,118,30,118,29,165,31,14,31,239,31,198,31,103,31,11,31,11,30,11,29,248,31,248,30,248,29,51,31,51,30,65,31,110,31,213,31,28,31,135,31,100,31,36,31,241,31,241,30,203,31,51,31,135,31,135,30,135,29,198,31,24,31,22,31,30,31,104,31,135,31,135,30,68,31,106,31,9,31,181,31,223,31,192,31,90,31,66,31,253,31,185,31,185,30,185,29,196,31,31,31,74,31,122,31,193,31,110,31,217,31,217,30,6,31,236,31,62,31,62,30,182,31,2,31,2,30,2,29,240,31,53,31,192,31,192,30,118,31,142,31,4,31,4,30,244,31,12,31,68,31,44,31,238,31,21,31,21,30,186,31,106,31,153,31,30,31,57,31,57,30,152,31,245,31,196,31,174,31,112,31,249,31,150,31,150,30,220,31,10,31,4,31,80,31,180,31,128,31,68,31,31,31,232,31,172,31,255,31,10,31,19,31,144,31,102,31,195,31,218,31,194,31,108,31,198,31,43,31,10,31,10,30,195,31,66,31,66,30,207,31,94,31,94,30,94,29,145,31,97,31,154,31,96,31,97,31,241,31,177,31,240,31,240,30,50,31,180,31,92,31,5,31,169,31,18,31,107,31,209,31,247,31,151,31,98,31,190,31,82,31,103,31,103,30,103,29,103,28,103,27,103,26,154,31,71,31,71,30,96,31,11,31,163,31,166,31,166,30,127,31,169,31,169,30,41,31,41,30,41,29,41,28,41,27,41,31,249,31,137,31,121,31,135,31,135,30,246,31,246,30,190,31,190,30,190,29,190,28,182,31,144,31,144,30,129,31,129,30,181,31,40,31,100,31,243,31,243,30,243,29,235,31,116,31,243,31,194,31,114,31,212,31,212,30,119,31,198,31,110,31,66,31,159,31,61,31,225,31,225,30,85,31,85,30,4,31,157,31,78,31,5,31,53,31,53,30,53,29,53,28,224,31,149,31,125,31,46,31,58,31,242,31,242,30,120,31,120,30,93,31,167,31,38,31,51,31,51,30,51,29,51,28,51,27,51,26,44,31,140,31,232,31,115,31,115,30,115,29,115,28,203,31,237,31,237,30,65,31,242,31,126,31,92,31,92,30,27,31,159,31,234,31,53,31,227,31,120,31,166,31,143,31,94,31,204,31,18,31,18,30,82,31,72,31,144,31,174,31,187,31,75,31,246,31,117,31,42,31,93,31,93,30,146,31,74,31,119,31,211,31,75,31,75,30,75,29,75,28,99,31,79,31,56,31,56,30,45,31,71,31,173,31,121,31,208,31,208,30,190,31,33,31,33,30,77,31,193,31,37,31,138,31,203,31,18,31,158,31,158,30,28,31,28,30,81,31,102,31,102,30,132,31,106,31,106,30,4,31,77,31,163,31,205,31,85,31,149,31,188,31,243,31,165,31,165,30,165,29,24,31,16,31,10,31,110,31,94,31,68,31,68,30,68,29,68,28,162,31,240,31,38,31,25,31,156,31,156,30,88,31,67,31,246,31,245,31,245,30,245,29,133,31,251,31,158,31,144,31,64,31,30,31,176,31,207,31,200,31,66,31,201,31,5,31,5,30,61,31,241,31,149,31,209,31,209,30,169,31,211,31,123,31,184,31,46,31,144,31,141,31,132,31,198,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
