-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_211 is
end project_tb_211;

architecture project_tb_arch_211 of project_tb_211 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 504;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (2,0,18,0,57,0,0,0,170,0,32,0,15,0,0,0,184,0,198,0,192,0,215,0,214,0,62,0,29,0,0,0,0,0,0,0,0,0,0,0,97,0,0,0,239,0,178,0,0,0,0,0,226,0,218,0,42,0,21,0,76,0,0,0,161,0,52,0,25,0,43,0,71,0,194,0,196,0,193,0,103,0,0,0,0,0,156,0,145,0,121,0,13,0,47,0,153,0,179,0,230,0,61,0,254,0,68,0,144,0,0,0,88,0,107,0,219,0,71,0,223,0,56,0,86,0,0,0,221,0,64,0,107,0,0,0,237,0,17,0,9,0,91,0,224,0,188,0,0,0,239,0,63,0,96,0,92,0,0,0,250,0,4,0,40,0,223,0,227,0,19,0,107,0,181,0,0,0,161,0,0,0,155,0,242,0,66,0,225,0,133,0,46,0,133,0,217,0,172,0,0,0,19,0,165,0,56,0,159,0,222,0,217,0,31,0,115,0,81,0,0,0,5,0,165,0,0,0,250,0,28,0,29,0,241,0,227,0,0,0,114,0,89,0,238,0,152,0,28,0,53,0,0,0,15,0,0,0,166,0,170,0,129,0,76,0,130,0,36,0,36,0,110,0,67,0,76,0,149,0,219,0,186,0,148,0,235,0,0,0,55,0,151,0,38,0,137,0,0,0,151,0,237,0,65,0,0,0,193,0,226,0,157,0,239,0,179,0,106,0,52,0,160,0,8,0,125,0,46,0,82,0,0,0,219,0,45,0,121,0,0,0,86,0,0,0,241,0,107,0,146,0,0,0,105,0,163,0,137,0,213,0,17,0,123,0,29,0,0,0,0,0,10,0,140,0,0,0,93,0,89,0,187,0,47,0,170,0,59,0,0,0,192,0,0,0,48,0,187,0,162,0,176,0,81,0,215,0,185,0,247,0,57,0,111,0,67,0,102,0,15,0,240,0,76,0,38,0,0,0,116,0,171,0,154,0,133,0,155,0,101,0,251,0,110,0,158,0,112,0,71,0,190,0,194,0,35,0,170,0,0,0,81,0,50,0,0,0,167,0,0,0,0,0,253,0,120,0,152,0,0,0,36,0,178,0,20,0,0,0,0,0,0,0,89,0,0,0,36,0,34,0,104,0,68,0,0,0,86,0,140,0,77,0,132,0,137,0,235,0,49,0,0,0,201,0,107,0,0,0,249,0,127,0,12,0,60,0,0,0,230,0,38,0,0,0,78,0,56,0,66,0,175,0,136,0,0,0,29,0,76,0,22,0,250,0,167,0,205,0,127,0,162,0,144,0,96,0,251,0,142,0,7,0,210,0,85,0,208,0,3,0,12,0,170,0,0,0,92,0,83,0,131,0,87,0,7,0,0,0,110,0,221,0,184,0,219,0,238,0,233,0,0,0,52,0,8,0,121,0,247,0,114,0,4,0,0,0,77,0,147,0,154,0,173,0,16,0,193,0,187,0,220,0,4,0,100,0,228,0,88,0,0,0,53,0,42,0,170,0,0,0,54,0,111,0,40,0,127,0,10,0,97,0,107,0,228,0,0,0,38,0,79,0,70,0,0,0,0,0,0,0,126,0,75,0,141,0,129,0,141,0,77,0,255,0,0,0,0,0,72,0,142,0,232,0,95,0,0,0,81,0,67,0,0,0,98,0,29,0,149,0,216,0,147,0,136,0,103,0,220,0,127,0,73,0,30,0,203,0,37,0,186,0,0,0,12,0,195,0,3,0,73,0,0,0,13,0,104,0,32,0,109,0,148,0,0,0,80,0,178,0,75,0,94,0,75,0,151,0,188,0,0,0,66,0,212,0,177,0,224,0,73,0,0,0,247,0,219,0,3,0,25,0,82,0,156,0,0,0,0,0,90,0,137,0,149,0,0,0,21,0,148,0,253,0,0,0,139,0,27,0,158,0,156,0,174,0,105,0,116,0,28,0,230,0,19,0,2,0,0,0,78,0,246,0,110,0,54,0,0,0,154,0,248,0,25,0,189,0,6,0,135,0,221,0,82,0,29,0,199,0,70,0,0,0,251,0,40,0,22,0,249,0,69,0,230,0,83,0,249,0,70,0,0,0,46,0,253,0,177,0,0,0,118,0,125,0,196,0,255,0,0,0,237,0,0,0,0,0,163,0,152,0,0,0,0,0,50,0,27,0,79,0,0,0,10,0,0,0,8,0,131,0,0,0,227,0,0,0,1,0,0,0,0,0,208,0,20,0,154,0,39,0,34,0,172,0,148,0,205,0,101,0,0,0,28,0);
signal scenario_full  : scenario_type := (2,31,18,31,57,31,57,30,170,31,32,31,15,31,15,30,184,31,198,31,192,31,215,31,214,31,62,31,29,31,29,30,29,29,29,28,29,27,29,26,97,31,97,30,239,31,178,31,178,30,178,29,226,31,218,31,42,31,21,31,76,31,76,30,161,31,52,31,25,31,43,31,71,31,194,31,196,31,193,31,103,31,103,30,103,29,156,31,145,31,121,31,13,31,47,31,153,31,179,31,230,31,61,31,254,31,68,31,144,31,144,30,88,31,107,31,219,31,71,31,223,31,56,31,86,31,86,30,221,31,64,31,107,31,107,30,237,31,17,31,9,31,91,31,224,31,188,31,188,30,239,31,63,31,96,31,92,31,92,30,250,31,4,31,40,31,223,31,227,31,19,31,107,31,181,31,181,30,161,31,161,30,155,31,242,31,66,31,225,31,133,31,46,31,133,31,217,31,172,31,172,30,19,31,165,31,56,31,159,31,222,31,217,31,31,31,115,31,81,31,81,30,5,31,165,31,165,30,250,31,28,31,29,31,241,31,227,31,227,30,114,31,89,31,238,31,152,31,28,31,53,31,53,30,15,31,15,30,166,31,170,31,129,31,76,31,130,31,36,31,36,31,110,31,67,31,76,31,149,31,219,31,186,31,148,31,235,31,235,30,55,31,151,31,38,31,137,31,137,30,151,31,237,31,65,31,65,30,193,31,226,31,157,31,239,31,179,31,106,31,52,31,160,31,8,31,125,31,46,31,82,31,82,30,219,31,45,31,121,31,121,30,86,31,86,30,241,31,107,31,146,31,146,30,105,31,163,31,137,31,213,31,17,31,123,31,29,31,29,30,29,29,10,31,140,31,140,30,93,31,89,31,187,31,47,31,170,31,59,31,59,30,192,31,192,30,48,31,187,31,162,31,176,31,81,31,215,31,185,31,247,31,57,31,111,31,67,31,102,31,15,31,240,31,76,31,38,31,38,30,116,31,171,31,154,31,133,31,155,31,101,31,251,31,110,31,158,31,112,31,71,31,190,31,194,31,35,31,170,31,170,30,81,31,50,31,50,30,167,31,167,30,167,29,253,31,120,31,152,31,152,30,36,31,178,31,20,31,20,30,20,29,20,28,89,31,89,30,36,31,34,31,104,31,68,31,68,30,86,31,140,31,77,31,132,31,137,31,235,31,49,31,49,30,201,31,107,31,107,30,249,31,127,31,12,31,60,31,60,30,230,31,38,31,38,30,78,31,56,31,66,31,175,31,136,31,136,30,29,31,76,31,22,31,250,31,167,31,205,31,127,31,162,31,144,31,96,31,251,31,142,31,7,31,210,31,85,31,208,31,3,31,12,31,170,31,170,30,92,31,83,31,131,31,87,31,7,31,7,30,110,31,221,31,184,31,219,31,238,31,233,31,233,30,52,31,8,31,121,31,247,31,114,31,4,31,4,30,77,31,147,31,154,31,173,31,16,31,193,31,187,31,220,31,4,31,100,31,228,31,88,31,88,30,53,31,42,31,170,31,170,30,54,31,111,31,40,31,127,31,10,31,97,31,107,31,228,31,228,30,38,31,79,31,70,31,70,30,70,29,70,28,126,31,75,31,141,31,129,31,141,31,77,31,255,31,255,30,255,29,72,31,142,31,232,31,95,31,95,30,81,31,67,31,67,30,98,31,29,31,149,31,216,31,147,31,136,31,103,31,220,31,127,31,73,31,30,31,203,31,37,31,186,31,186,30,12,31,195,31,3,31,73,31,73,30,13,31,104,31,32,31,109,31,148,31,148,30,80,31,178,31,75,31,94,31,75,31,151,31,188,31,188,30,66,31,212,31,177,31,224,31,73,31,73,30,247,31,219,31,3,31,25,31,82,31,156,31,156,30,156,29,90,31,137,31,149,31,149,30,21,31,148,31,253,31,253,30,139,31,27,31,158,31,156,31,174,31,105,31,116,31,28,31,230,31,19,31,2,31,2,30,78,31,246,31,110,31,54,31,54,30,154,31,248,31,25,31,189,31,6,31,135,31,221,31,82,31,29,31,199,31,70,31,70,30,251,31,40,31,22,31,249,31,69,31,230,31,83,31,249,31,70,31,70,30,46,31,253,31,177,31,177,30,118,31,125,31,196,31,255,31,255,30,237,31,237,30,237,29,163,31,152,31,152,30,152,29,50,31,27,31,79,31,79,30,10,31,10,30,8,31,131,31,131,30,227,31,227,30,1,31,1,30,1,29,208,31,20,31,154,31,39,31,34,31,172,31,148,31,205,31,101,31,101,30,28,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
