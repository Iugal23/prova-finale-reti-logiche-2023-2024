-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_297 is
end project_tb_297;

architecture project_tb_arch_297 of project_tb_297 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 913;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (201,0,3,0,172,0,71,0,88,0,0,0,82,0,229,0,0,0,30,0,251,0,215,0,142,0,49,0,48,0,180,0,0,0,0,0,80,0,72,0,204,0,145,0,223,0,117,0,23,0,246,0,109,0,179,0,241,0,189,0,54,0,0,0,0,0,152,0,55,0,74,0,16,0,174,0,37,0,227,0,0,0,0,0,184,0,218,0,248,0,42,0,162,0,172,0,145,0,55,0,101,0,110,0,254,0,107,0,45,0,112,0,0,0,194,0,74,0,46,0,228,0,209,0,52,0,155,0,0,0,128,0,252,0,164,0,191,0,0,0,167,0,35,0,162,0,81,0,188,0,0,0,47,0,179,0,0,0,157,0,119,0,86,0,0,0,62,0,131,0,0,0,162,0,154,0,222,0,197,0,169,0,189,0,33,0,175,0,193,0,201,0,113,0,0,0,195,0,64,0,250,0,147,0,227,0,207,0,12,0,205,0,97,0,168,0,171,0,218,0,0,0,59,0,42,0,0,0,114,0,252,0,29,0,109,0,232,0,0,0,0,0,253,0,0,0,255,0,66,0,0,0,202,0,50,0,0,0,56,0,142,0,58,0,178,0,212,0,66,0,131,0,221,0,245,0,31,0,75,0,22,0,0,0,181,0,0,0,142,0,165,0,17,0,231,0,60,0,0,0,0,0,205,0,5,0,0,0,121,0,0,0,15,0,28,0,240,0,208,0,116,0,22,0,227,0,196,0,159,0,116,0,0,0,234,0,139,0,134,0,254,0,0,0,242,0,53,0,10,0,116,0,81,0,214,0,20,0,0,0,103,0,32,0,0,0,13,0,12,0,66,0,0,0,36,0,38,0,34,0,145,0,0,0,208,0,8,0,155,0,133,0,57,0,181,0,231,0,201,0,8,0,0,0,247,0,142,0,0,0,112,0,255,0,37,0,16,0,55,0,217,0,35,0,102,0,35,0,209,0,0,0,0,0,0,0,189,0,65,0,112,0,206,0,0,0,73,0,171,0,8,0,28,0,159,0,23,0,113,0,0,0,0,0,153,0,0,0,70,0,49,0,232,0,64,0,246,0,180,0,224,0,188,0,83,0,229,0,190,0,234,0,226,0,0,0,0,0,184,0,111,0,0,0,75,0,0,0,0,0,0,0,239,0,0,0,143,0,184,0,241,0,0,0,255,0,174,0,143,0,185,0,42,0,7,0,133,0,0,0,65,0,129,0,253,0,71,0,118,0,124,0,35,0,0,0,126,0,0,0,224,0,0,0,186,0,2,0,28,0,226,0,202,0,79,0,0,0,0,0,139,0,116,0,0,0,0,0,205,0,89,0,196,0,160,0,37,0,129,0,140,0,179,0,215,0,83,0,31,0,116,0,136,0,180,0,88,0,0,0,37,0,179,0,150,0,0,0,92,0,217,0,6,0,60,0,96,0,16,0,225,0,232,0,0,0,65,0,9,0,94,0,106,0,140,0,0,0,0,0,242,0,0,0,78,0,0,0,141,0,89,0,0,0,147,0,54,0,191,0,172,0,150,0,80,0,251,0,205,0,19,0,0,0,190,0,136,0,48,0,118,0,154,0,0,0,130,0,229,0,18,0,31,0,101,0,0,0,234,0,245,0,128,0,207,0,24,0,159,0,234,0,150,0,221,0,79,0,0,0,213,0,89,0,194,0,160,0,149,0,0,0,119,0,68,0,238,0,43,0,95,0,191,0,134,0,212,0,72,0,56,0,115,0,230,0,46,0,254,0,9,0,91,0,152,0,11,0,203,0,218,0,148,0,146,0,227,0,235,0,216,0,181,0,29,0,170,0,0,0,0,0,81,0,0,0,106,0,94,0,253,0,29,0,51,0,141,0,181,0,0,0,165,0,160,0,211,0,129,0,22,0,184,0,149,0,121,0,85,0,235,0,190,0,61,0,65,0,0,0,252,0,0,0,112,0,175,0,66,0,23,0,5,0,0,0,194,0,171,0,196,0,0,0,127,0,173,0,133,0,0,0,114,0,216,0,23,0,0,0,219,0,74,0,254,0,238,0,119,0,115,0,121,0,236,0,62,0,0,0,15,0,17,0,83,0,237,0,4,0,16,0,178,0,20,0,33,0,65,0,51,0,0,0,0,0,253,0,225,0,108,0,255,0,250,0,158,0,0,0,88,0,23,0,196,0,174,0,0,0,106,0,144,0,0,0,234,0,134,0,107,0,212,0,52,0,54,0,150,0,152,0,210,0,53,0,228,0,75,0,0,0,232,0,0,0,255,0,127,0,177,0,251,0,154,0,5,0,0,0,132,0,89,0,54,0,239,0,229,0,249,0,0,0,189,0,60,0,218,0,119,0,147,0,240,0,137,0,122,0,104,0,53,0,73,0,107,0,242,0,188,0,0,0,27,0,157,0,156,0,20,0,169,0,206,0,13,0,70,0,0,0,79,0,122,0,0,0,0,0,83,0,175,0,189,0,39,0,254,0,0,0,6,0,45,0,141,0,99,0,62,0,232,0,93,0,54,0,99,0,185,0,218,0,0,0,0,0,235,0,130,0,94,0,32,0,210,0,49,0,39,0,86,0,192,0,210,0,254,0,0,0,93,0,0,0,176,0,0,0,0,0,140,0,141,0,0,0,82,0,98,0,0,0,126,0,210,0,8,0,44,0,0,0,244,0,0,0,0,0,0,0,253,0,0,0,107,0,0,0,0,0,94,0,224,0,199,0,213,0,134,0,215,0,240,0,0,0,0,0,41,0,0,0,0,0,222,0,72,0,154,0,17,0,195,0,217,0,164,0,98,0,160,0,134,0,178,0,152,0,40,0,4,0,155,0,4,0,0,0,104,0,40,0,2,0,240,0,214,0,205,0,202,0,0,0,126,0,62,0,178,0,34,0,188,0,64,0,203,0,50,0,185,0,142,0,38,0,0,0,144,0,49,0,0,0,251,0,24,0,0,0,0,0,5,0,192,0,138,0,0,0,52,0,190,0,255,0,31,0,119,0,185,0,147,0,200,0,55,0,87,0,41,0,125,0,173,0,56,0,240,0,44,0,197,0,84,0,130,0,106,0,248,0,172,0,87,0,36,0,168,0,143,0,0,0,235,0,55,0,49,0,0,0,209,0,87,0,109,0,141,0,213,0,0,0,0,0,235,0,0,0,221,0,59,0,178,0,190,0,0,0,42,0,76,0,1,0,52,0,70,0,99,0,0,0,234,0,0,0,174,0,130,0,224,0,0,0,0,0,237,0,58,0,0,0,22,0,120,0,68,0,0,0,218,0,0,0,84,0,183,0,56,0,93,0,216,0,233,0,91,0,173,0,36,0,103,0,79,0,27,0,126,0,65,0,120,0,244,0,208,0,74,0,0,0,149,0,197,0,138,0,32,0,15,0,74,0,0,0,81,0,92,0,171,0,175,0,152,0,80,0,0,0,85,0,150,0,237,0,116,0,0,0,91,0,130,0,124,0,90,0,0,0,0,0,187,0,165,0,13,0,4,0,162,0,220,0,240,0,0,0,80,0,43,0,13,0,5,0,0,0,0,0,249,0,206,0,27,0,231,0,0,0,0,0,65,0,162,0,0,0,173,0,31,0,86,0,244,0,7,0,91,0,55,0,30,0,165,0,0,0,243,0,136,0,219,0,0,0,15,0,207,0,0,0,0,0,0,0,9,0,189,0,0,0,70,0,92,0,57,0,0,0,0,0,200,0,119,0,235,0,0,0,120,0,207,0,194,0,13,0,140,0,166,0,0,0,177,0,16,0,65,0,14,0,71,0,60,0,207,0,174,0,0,0,249,0,222,0,234,0,119,0,21,0,210,0,48,0,0,0,126,0,28,0,109,0,153,0,135,0,199,0,152,0,163,0,24,0,103,0,0,0,134,0,0,0,219,0,47,0,219,0,0,0,131,0,110,0,58,0,0,0,50,0,201,0,28,0,244,0,0,0,119,0,91,0,105,0,210,0,77,0,0,0,0,0,40,0,183,0,234,0,0,0,26,0,108,0,18,0,42,0,213,0,51,0,0,0,151,0,107,0,192,0,72,0,81,0,0,0,124,0,184,0,120,0,131,0,241,0,255,0,13,0,211,0,142,0,0,0,47,0,0,0);
signal scenario_full  : scenario_type := (201,31,3,31,172,31,71,31,88,31,88,30,82,31,229,31,229,30,30,31,251,31,215,31,142,31,49,31,48,31,180,31,180,30,180,29,80,31,72,31,204,31,145,31,223,31,117,31,23,31,246,31,109,31,179,31,241,31,189,31,54,31,54,30,54,29,152,31,55,31,74,31,16,31,174,31,37,31,227,31,227,30,227,29,184,31,218,31,248,31,42,31,162,31,172,31,145,31,55,31,101,31,110,31,254,31,107,31,45,31,112,31,112,30,194,31,74,31,46,31,228,31,209,31,52,31,155,31,155,30,128,31,252,31,164,31,191,31,191,30,167,31,35,31,162,31,81,31,188,31,188,30,47,31,179,31,179,30,157,31,119,31,86,31,86,30,62,31,131,31,131,30,162,31,154,31,222,31,197,31,169,31,189,31,33,31,175,31,193,31,201,31,113,31,113,30,195,31,64,31,250,31,147,31,227,31,207,31,12,31,205,31,97,31,168,31,171,31,218,31,218,30,59,31,42,31,42,30,114,31,252,31,29,31,109,31,232,31,232,30,232,29,253,31,253,30,255,31,66,31,66,30,202,31,50,31,50,30,56,31,142,31,58,31,178,31,212,31,66,31,131,31,221,31,245,31,31,31,75,31,22,31,22,30,181,31,181,30,142,31,165,31,17,31,231,31,60,31,60,30,60,29,205,31,5,31,5,30,121,31,121,30,15,31,28,31,240,31,208,31,116,31,22,31,227,31,196,31,159,31,116,31,116,30,234,31,139,31,134,31,254,31,254,30,242,31,53,31,10,31,116,31,81,31,214,31,20,31,20,30,103,31,32,31,32,30,13,31,12,31,66,31,66,30,36,31,38,31,34,31,145,31,145,30,208,31,8,31,155,31,133,31,57,31,181,31,231,31,201,31,8,31,8,30,247,31,142,31,142,30,112,31,255,31,37,31,16,31,55,31,217,31,35,31,102,31,35,31,209,31,209,30,209,29,209,28,189,31,65,31,112,31,206,31,206,30,73,31,171,31,8,31,28,31,159,31,23,31,113,31,113,30,113,29,153,31,153,30,70,31,49,31,232,31,64,31,246,31,180,31,224,31,188,31,83,31,229,31,190,31,234,31,226,31,226,30,226,29,184,31,111,31,111,30,75,31,75,30,75,29,75,28,239,31,239,30,143,31,184,31,241,31,241,30,255,31,174,31,143,31,185,31,42,31,7,31,133,31,133,30,65,31,129,31,253,31,71,31,118,31,124,31,35,31,35,30,126,31,126,30,224,31,224,30,186,31,2,31,28,31,226,31,202,31,79,31,79,30,79,29,139,31,116,31,116,30,116,29,205,31,89,31,196,31,160,31,37,31,129,31,140,31,179,31,215,31,83,31,31,31,116,31,136,31,180,31,88,31,88,30,37,31,179,31,150,31,150,30,92,31,217,31,6,31,60,31,96,31,16,31,225,31,232,31,232,30,65,31,9,31,94,31,106,31,140,31,140,30,140,29,242,31,242,30,78,31,78,30,141,31,89,31,89,30,147,31,54,31,191,31,172,31,150,31,80,31,251,31,205,31,19,31,19,30,190,31,136,31,48,31,118,31,154,31,154,30,130,31,229,31,18,31,31,31,101,31,101,30,234,31,245,31,128,31,207,31,24,31,159,31,234,31,150,31,221,31,79,31,79,30,213,31,89,31,194,31,160,31,149,31,149,30,119,31,68,31,238,31,43,31,95,31,191,31,134,31,212,31,72,31,56,31,115,31,230,31,46,31,254,31,9,31,91,31,152,31,11,31,203,31,218,31,148,31,146,31,227,31,235,31,216,31,181,31,29,31,170,31,170,30,170,29,81,31,81,30,106,31,94,31,253,31,29,31,51,31,141,31,181,31,181,30,165,31,160,31,211,31,129,31,22,31,184,31,149,31,121,31,85,31,235,31,190,31,61,31,65,31,65,30,252,31,252,30,112,31,175,31,66,31,23,31,5,31,5,30,194,31,171,31,196,31,196,30,127,31,173,31,133,31,133,30,114,31,216,31,23,31,23,30,219,31,74,31,254,31,238,31,119,31,115,31,121,31,236,31,62,31,62,30,15,31,17,31,83,31,237,31,4,31,16,31,178,31,20,31,33,31,65,31,51,31,51,30,51,29,253,31,225,31,108,31,255,31,250,31,158,31,158,30,88,31,23,31,196,31,174,31,174,30,106,31,144,31,144,30,234,31,134,31,107,31,212,31,52,31,54,31,150,31,152,31,210,31,53,31,228,31,75,31,75,30,232,31,232,30,255,31,127,31,177,31,251,31,154,31,5,31,5,30,132,31,89,31,54,31,239,31,229,31,249,31,249,30,189,31,60,31,218,31,119,31,147,31,240,31,137,31,122,31,104,31,53,31,73,31,107,31,242,31,188,31,188,30,27,31,157,31,156,31,20,31,169,31,206,31,13,31,70,31,70,30,79,31,122,31,122,30,122,29,83,31,175,31,189,31,39,31,254,31,254,30,6,31,45,31,141,31,99,31,62,31,232,31,93,31,54,31,99,31,185,31,218,31,218,30,218,29,235,31,130,31,94,31,32,31,210,31,49,31,39,31,86,31,192,31,210,31,254,31,254,30,93,31,93,30,176,31,176,30,176,29,140,31,141,31,141,30,82,31,98,31,98,30,126,31,210,31,8,31,44,31,44,30,244,31,244,30,244,29,244,28,253,31,253,30,107,31,107,30,107,29,94,31,224,31,199,31,213,31,134,31,215,31,240,31,240,30,240,29,41,31,41,30,41,29,222,31,72,31,154,31,17,31,195,31,217,31,164,31,98,31,160,31,134,31,178,31,152,31,40,31,4,31,155,31,4,31,4,30,104,31,40,31,2,31,240,31,214,31,205,31,202,31,202,30,126,31,62,31,178,31,34,31,188,31,64,31,203,31,50,31,185,31,142,31,38,31,38,30,144,31,49,31,49,30,251,31,24,31,24,30,24,29,5,31,192,31,138,31,138,30,52,31,190,31,255,31,31,31,119,31,185,31,147,31,200,31,55,31,87,31,41,31,125,31,173,31,56,31,240,31,44,31,197,31,84,31,130,31,106,31,248,31,172,31,87,31,36,31,168,31,143,31,143,30,235,31,55,31,49,31,49,30,209,31,87,31,109,31,141,31,213,31,213,30,213,29,235,31,235,30,221,31,59,31,178,31,190,31,190,30,42,31,76,31,1,31,52,31,70,31,99,31,99,30,234,31,234,30,174,31,130,31,224,31,224,30,224,29,237,31,58,31,58,30,22,31,120,31,68,31,68,30,218,31,218,30,84,31,183,31,56,31,93,31,216,31,233,31,91,31,173,31,36,31,103,31,79,31,27,31,126,31,65,31,120,31,244,31,208,31,74,31,74,30,149,31,197,31,138,31,32,31,15,31,74,31,74,30,81,31,92,31,171,31,175,31,152,31,80,31,80,30,85,31,150,31,237,31,116,31,116,30,91,31,130,31,124,31,90,31,90,30,90,29,187,31,165,31,13,31,4,31,162,31,220,31,240,31,240,30,80,31,43,31,13,31,5,31,5,30,5,29,249,31,206,31,27,31,231,31,231,30,231,29,65,31,162,31,162,30,173,31,31,31,86,31,244,31,7,31,91,31,55,31,30,31,165,31,165,30,243,31,136,31,219,31,219,30,15,31,207,31,207,30,207,29,207,28,9,31,189,31,189,30,70,31,92,31,57,31,57,30,57,29,200,31,119,31,235,31,235,30,120,31,207,31,194,31,13,31,140,31,166,31,166,30,177,31,16,31,65,31,14,31,71,31,60,31,207,31,174,31,174,30,249,31,222,31,234,31,119,31,21,31,210,31,48,31,48,30,126,31,28,31,109,31,153,31,135,31,199,31,152,31,163,31,24,31,103,31,103,30,134,31,134,30,219,31,47,31,219,31,219,30,131,31,110,31,58,31,58,30,50,31,201,31,28,31,244,31,244,30,119,31,91,31,105,31,210,31,77,31,77,30,77,29,40,31,183,31,234,31,234,30,26,31,108,31,18,31,42,31,213,31,51,31,51,30,151,31,107,31,192,31,72,31,81,31,81,30,124,31,184,31,120,31,131,31,241,31,255,31,13,31,211,31,142,31,142,30,47,31,47,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
