-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 423;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (13,0,244,0,7,0,146,0,174,0,0,0,0,0,139,0,169,0,50,0,102,0,157,0,0,0,64,0,203,0,7,0,113,0,214,0,238,0,0,0,0,0,223,0,182,0,0,0,34,0,101,0,129,0,216,0,220,0,245,0,0,0,148,0,111,0,111,0,39,0,0,0,148,0,190,0,0,0,251,0,191,0,100,0,109,0,30,0,10,0,0,0,39,0,64,0,236,0,0,0,208,0,92,0,4,0,0,0,0,0,191,0,0,0,117,0,221,0,12,0,0,0,0,0,5,0,217,0,0,0,63,0,27,0,222,0,44,0,0,0,0,0,0,0,8,0,234,0,32,0,244,0,200,0,0,0,171,0,8,0,106,0,233,0,208,0,154,0,3,0,206,0,0,0,57,0,38,0,0,0,220,0,195,0,158,0,32,0,241,0,21,0,140,0,62,0,33,0,65,0,0,0,0,0,0,0,0,0,205,0,252,0,0,0,219,0,52,0,215,0,150,0,80,0,220,0,152,0,56,0,0,0,173,0,79,0,125,0,187,0,153,0,130,0,226,0,0,0,0,0,0,0,213,0,21,0,0,0,0,0,220,0,169,0,179,0,106,0,0,0,0,0,0,0,38,0,62,0,33,0,218,0,228,0,0,0,107,0,0,0,0,0,191,0,25,0,129,0,234,0,0,0,79,0,184,0,68,0,166,0,141,0,219,0,153,0,213,0,217,0,228,0,143,0,74,0,169,0,137,0,45,0,133,0,184,0,40,0,73,0,52,0,0,0,151,0,0,0,11,0,238,0,122,0,68,0,0,0,0,0,108,0,147,0,92,0,156,0,66,0,243,0,15,0,116,0,0,0,161,0,131,0,0,0,220,0,110,0,82,0,0,0,141,0,61,0,34,0,0,0,222,0,176,0,236,0,0,0,206,0,36,0,83,0,169,0,249,0,239,0,0,0,79,0,148,0,160,0,91,0,56,0,136,0,129,0,72,0,134,0,179,0,204,0,48,0,68,0,64,0,225,0,4,0,0,0,46,0,2,0,62,0,234,0,0,0,154,0,28,0,253,0,105,0,251,0,95,0,242,0,165,0,38,0,74,0,145,0,196,0,146,0,152,0,55,0,57,0,187,0,224,0,0,0,88,0,139,0,0,0,168,0,240,0,2,0,212,0,56,0,97,0,157,0,167,0,83,0,12,0,0,0,182,0,10,0,234,0,222,0,154,0,36,0,0,0,0,0,0,0,85,0,0,0,0,0,107,0,7,0,0,0,189,0,61,0,172,0,131,0,145,0,0,0,36,0,113,0,122,0,231,0,75,0,242,0,164,0,23,0,0,0,8,0,243,0,28,0,189,0,0,0,0,0,170,0,43,0,0,0,211,0,161,0,0,0,80,0,0,0,0,0,0,0,64,0,0,0,96,0,0,0,9,0,0,0,0,0,31,0,20,0,20,0,189,0,28,0,148,0,128,0,94,0,252,0,97,0,0,0,208,0,185,0,148,0,4,0,215,0,7,0,231,0,170,0,198,0,0,0,74,0,100,0,0,0,40,0,249,0,176,0,225,0,228,0,0,0,39,0,248,0,0,0,42,0,65,0,49,0,196,0,164,0,25,0,13,0,178,0,67,0,0,0,61,0,235,0,232,0,0,0,36,0,0,0,128,0,210,0,20,0,129,0,234,0,0,0,165,0,0,0,6,0,255,0,51,0,167,0,212,0,121,0,97,0,61,0,124,0,0,0,135,0,211,0,62,0,210,0,208,0,172,0,33,0,26,0,39,0,203,0,221,0,92,0,224,0,0,0,6,0,243,0,92,0,166,0,159,0,153,0,203,0,225,0,0,0,161,0,2,0,21,0,0,0,138,0,42,0,46,0,0,0,132,0,0,0,149,0,149,0,57,0,0,0);
signal scenario_full  : scenario_type := (13,31,244,31,7,31,146,31,174,31,174,30,174,29,139,31,169,31,50,31,102,31,157,31,157,30,64,31,203,31,7,31,113,31,214,31,238,31,238,30,238,29,223,31,182,31,182,30,34,31,101,31,129,31,216,31,220,31,245,31,245,30,148,31,111,31,111,31,39,31,39,30,148,31,190,31,190,30,251,31,191,31,100,31,109,31,30,31,10,31,10,30,39,31,64,31,236,31,236,30,208,31,92,31,4,31,4,30,4,29,191,31,191,30,117,31,221,31,12,31,12,30,12,29,5,31,217,31,217,30,63,31,27,31,222,31,44,31,44,30,44,29,44,28,8,31,234,31,32,31,244,31,200,31,200,30,171,31,8,31,106,31,233,31,208,31,154,31,3,31,206,31,206,30,57,31,38,31,38,30,220,31,195,31,158,31,32,31,241,31,21,31,140,31,62,31,33,31,65,31,65,30,65,29,65,28,65,27,205,31,252,31,252,30,219,31,52,31,215,31,150,31,80,31,220,31,152,31,56,31,56,30,173,31,79,31,125,31,187,31,153,31,130,31,226,31,226,30,226,29,226,28,213,31,21,31,21,30,21,29,220,31,169,31,179,31,106,31,106,30,106,29,106,28,38,31,62,31,33,31,218,31,228,31,228,30,107,31,107,30,107,29,191,31,25,31,129,31,234,31,234,30,79,31,184,31,68,31,166,31,141,31,219,31,153,31,213,31,217,31,228,31,143,31,74,31,169,31,137,31,45,31,133,31,184,31,40,31,73,31,52,31,52,30,151,31,151,30,11,31,238,31,122,31,68,31,68,30,68,29,108,31,147,31,92,31,156,31,66,31,243,31,15,31,116,31,116,30,161,31,131,31,131,30,220,31,110,31,82,31,82,30,141,31,61,31,34,31,34,30,222,31,176,31,236,31,236,30,206,31,36,31,83,31,169,31,249,31,239,31,239,30,79,31,148,31,160,31,91,31,56,31,136,31,129,31,72,31,134,31,179,31,204,31,48,31,68,31,64,31,225,31,4,31,4,30,46,31,2,31,62,31,234,31,234,30,154,31,28,31,253,31,105,31,251,31,95,31,242,31,165,31,38,31,74,31,145,31,196,31,146,31,152,31,55,31,57,31,187,31,224,31,224,30,88,31,139,31,139,30,168,31,240,31,2,31,212,31,56,31,97,31,157,31,167,31,83,31,12,31,12,30,182,31,10,31,234,31,222,31,154,31,36,31,36,30,36,29,36,28,85,31,85,30,85,29,107,31,7,31,7,30,189,31,61,31,172,31,131,31,145,31,145,30,36,31,113,31,122,31,231,31,75,31,242,31,164,31,23,31,23,30,8,31,243,31,28,31,189,31,189,30,189,29,170,31,43,31,43,30,211,31,161,31,161,30,80,31,80,30,80,29,80,28,64,31,64,30,96,31,96,30,9,31,9,30,9,29,31,31,20,31,20,31,189,31,28,31,148,31,128,31,94,31,252,31,97,31,97,30,208,31,185,31,148,31,4,31,215,31,7,31,231,31,170,31,198,31,198,30,74,31,100,31,100,30,40,31,249,31,176,31,225,31,228,31,228,30,39,31,248,31,248,30,42,31,65,31,49,31,196,31,164,31,25,31,13,31,178,31,67,31,67,30,61,31,235,31,232,31,232,30,36,31,36,30,128,31,210,31,20,31,129,31,234,31,234,30,165,31,165,30,6,31,255,31,51,31,167,31,212,31,121,31,97,31,61,31,124,31,124,30,135,31,211,31,62,31,210,31,208,31,172,31,33,31,26,31,39,31,203,31,221,31,92,31,224,31,224,30,6,31,243,31,92,31,166,31,159,31,153,31,203,31,225,31,225,30,161,31,2,31,21,31,21,30,138,31,42,31,46,31,46,30,132,31,132,30,149,31,149,31,57,31,57,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
