-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_367 is
end project_tb_367;

architecture project_tb_arch_367 of project_tb_367 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 959;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,135,0,0,0,127,0,0,0,0,0,21,0,101,0,175,0,186,0,85,0,153,0,0,0,221,0,136,0,133,0,221,0,68,0,178,0,35,0,164,0,87,0,0,0,0,0,22,0,241,0,0,0,139,0,72,0,228,0,238,0,102,0,11,0,55,0,0,0,109,0,55,0,0,0,99,0,243,0,219,0,119,0,133,0,5,0,89,0,197,0,181,0,19,0,220,0,46,0,198,0,0,0,226,0,79,0,160,0,79,0,205,0,107,0,1,0,210,0,17,0,196,0,165,0,205,0,31,0,69,0,142,0,158,0,192,0,0,0,220,0,186,0,234,0,24,0,0,0,127,0,252,0,45,0,0,0,53,0,116,0,182,0,141,0,208,0,224,0,115,0,60,0,127,0,247,0,210,0,170,0,233,0,0,0,100,0,0,0,167,0,6,0,170,0,254,0,221,0,0,0,65,0,0,0,209,0,242,0,119,0,203,0,248,0,121,0,0,0,155,0,120,0,126,0,197,0,203,0,0,0,17,0,68,0,0,0,147,0,162,0,133,0,210,0,211,0,68,0,231,0,86,0,158,0,152,0,201,0,164,0,15,0,0,0,59,0,101,0,38,0,182,0,56,0,128,0,0,0,91,0,121,0,246,0,0,0,0,0,109,0,168,0,0,0,205,0,64,0,189,0,123,0,21,0,223,0,200,0,0,0,7,0,199,0,175,0,159,0,0,0,189,0,220,0,28,0,23,0,0,0,34,0,253,0,120,0,217,0,0,0,187,0,21,0,167,0,116,0,0,0,32,0,0,0,82,0,91,0,0,0,230,0,86,0,114,0,104,0,186,0,211,0,20,0,103,0,23,0,130,0,222,0,224,0,35,0,78,0,154,0,172,0,178,0,100,0,0,0,235,0,240,0,0,0,109,0,220,0,144,0,91,0,242,0,0,0,200,0,85,0,0,0,0,0,135,0,0,0,0,0,70,0,229,0,121,0,0,0,63,0,208,0,0,0,0,0,46,0,101,0,241,0,163,0,199,0,18,0,156,0,34,0,16,0,247,0,177,0,86,0,220,0,204,0,10,0,39,0,25,0,46,0,87,0,39,0,161,0,63,0,0,0,137,0,160,0,154,0,191,0,129,0,59,0,0,0,24,0,54,0,221,0,183,0,116,0,193,0,0,0,0,0,93,0,59,0,0,0,135,0,215,0,212,0,4,0,0,0,0,0,207,0,0,0,142,0,0,0,120,0,124,0,48,0,180,0,105,0,33,0,4,0,208,0,179,0,117,0,159,0,70,0,0,0,19,0,247,0,209,0,90,0,216,0,127,0,0,0,64,0,0,0,202,0,38,0,67,0,105,0,0,0,0,0,0,0,0,0,194,0,114,0,181,0,213,0,229,0,230,0,0,0,30,0,75,0,37,0,81,0,225,0,19,0,147,0,11,0,0,0,176,0,29,0,0,0,0,0,195,0,0,0,219,0,167,0,7,0,219,0,251,0,235,0,103,0,30,0,113,0,249,0,202,0,116,0,103,0,65,0,21,0,236,0,0,0,0,0,175,0,117,0,162,0,10,0,246,0,123,0,209,0,229,0,3,0,171,0,202,0,166,0,189,0,3,0,50,0,190,0,250,0,119,0,0,0,238,0,92,0,104,0,242,0,87,0,236,0,0,0,0,0,62,0,228,0,0,0,179,0,77,0,156,0,58,0,117,0,0,0,58,0,218,0,0,0,138,0,123,0,102,0,119,0,94,0,117,0,34,0,30,0,158,0,0,0,40,0,0,0,0,0,197,0,0,0,31,0,136,0,102,0,141,0,158,0,0,0,93,0,110,0,212,0,114,0,0,0,190,0,87,0,2,0,76,0,250,0,175,0,57,0,0,0,55,0,23,0,40,0,112,0,146,0,251,0,230,0,37,0,234,0,228,0,34,0,17,0,112,0,154,0,247,0,56,0,58,0,96,0,204,0,2,0,137,0,143,0,0,0,248,0,0,0,140,0,110,0,26,0,0,0,0,0,0,0,112,0,0,0,218,0,196,0,0,0,56,0,225,0,73,0,128,0,236,0,0,0,189,0,167,0,0,0,0,0,230,0,236,0,221,0,87,0,38,0,0,0,0,0,251,0,79,0,0,0,220,0,187,0,0,0,44,0,28,0,206,0,45,0,82,0,0,0,106,0,0,0,44,0,102,0,119,0,207,0,215,0,208,0,31,0,158,0,131,0,30,0,99,0,52,0,222,0,157,0,0,0,0,0,0,0,147,0,128,0,185,0,177,0,110,0,119,0,224,0,146,0,236,0,21,0,235,0,243,0,199,0,173,0,121,0,0,0,90,0,216,0,174,0,155,0,102,0,25,0,196,0,242,0,45,0,0,0,122,0,36,0,22,0,168,0,235,0,220,0,212,0,110,0,139,0,112,0,0,0,27,0,96,0,87,0,0,0,79,0,206,0,150,0,249,0,198,0,226,0,117,0,30,0,5,0,60,0,0,0,101,0,201,0,148,0,55,0,235,0,177,0,91,0,25,0,162,0,194,0,118,0,13,0,6,0,47,0,0,0,18,0,237,0,150,0,149,0,172,0,90,0,8,0,0,0,115,0,223,0,232,0,0,0,123,0,143,0,195,0,239,0,95,0,0,0,92,0,67,0,32,0,0,0,88,0,57,0,175,0,82,0,79,0,214,0,152,0,50,0,0,0,150,0,44,0,40,0,224,0,223,0,155,0,245,0,38,0,79,0,17,0,183,0,222,0,33,0,0,0,168,0,127,0,0,0,166,0,205,0,198,0,150,0,202,0,237,0,0,0,145,0,111,0,40,0,4,0,0,0,0,0,183,0,107,0,221,0,0,0,38,0,0,0,0,0,86,0,5,0,82,0,0,0,33,0,157,0,33,0,158,0,196,0,0,0,0,0,136,0,232,0,0,0,0,0,208,0,0,0,30,0,12,0,20,0,183,0,179,0,37,0,0,0,99,0,0,0,0,0,67,0,112,0,0,0,0,0,75,0,68,0,210,0,137,0,0,0,0,0,77,0,247,0,186,0,89,0,0,0,234,0,0,0,10,0,100,0,181,0,139,0,158,0,134,0,251,0,226,0,86,0,236,0,141,0,85,0,6,0,129,0,229,0,57,0,121,0,0,0,0,0,0,0,41,0,134,0,235,0,40,0,0,0,44,0,0,0,115,0,106,0,61,0,112,0,142,0,252,0,1,0,0,0,187,0,37,0,0,0,35,0,209,0,108,0,133,0,168,0,0,0,75,0,147,0,116,0,122,0,166,0,26,0,251,0,41,0,26,0,180,0,84,0,191,0,206,0,208,0,131,0,188,0,69,0,235,0,75,0,150,0,100,0,145,0,110,0,0,0,0,0,41,0,139,0,176,0,201,0,97,0,102,0,109,0,161,0,0,0,147,0,28,0,33,0,148,0,180,0,33,0,134,0,127,0,155,0,55,0,0,0,23,0,92,0,83,0,183,0,208,0,56,0,244,0,119,0,153,0,158,0,127,0,0,0,192,0,53,0,171,0,0,0,37,0,13,0,170,0,135,0,190,0,0,0,156,0,110,0,245,0,124,0,164,0,12,0,51,0,41,0,132,0,86,0,0,0,201,0,128,0,32,0,0,0,9,0,80,0,163,0,42,0,92,0,223,0,207,0,66,0,247,0,66,0,19,0,0,0,241,0,14,0,153,0,233,0,220,0,163,0,0,0,221,0,154,0,234,0,169,0,115,0,110,0,196,0,0,0,73,0,83,0,68,0,96,0,0,0,60,0,110,0,227,0,0,0,124,0,133,0,58,0,253,0,139,0,71,0,151,0,19,0,121,0,119,0,96,0,0,0,166,0,71,0,134,0,193,0,0,0,93,0,226,0,173,0,0,0,131,0,183,0,158,0,246,0,9,0,0,0,83,0,238,0,0,0,24,0,211,0,69,0,0,0,206,0,183,0,172,0,85,0,150,0,16,0,220,0,7,0,60,0,1,0,145,0,84,0,205,0,192,0,24,0,1,0,112,0,111,0,115,0,17,0,95,0,155,0,128,0,0,0,33,0,162,0,114,0,90,0,36,0,5,0,0,0,15,0,173,0,110,0,228,0,86,0,0,0,198,0,55,0,87,0,0,0,91,0,137,0,176,0,52,0,224,0,91,0,210,0,236,0,74,0,103,0,39,0,49,0,160,0,64,0,100,0,0,0,120,0,110,0,0,0,63,0,68,0,49,0,236,0,12,0,0,0,0,0,11,0,0,0,116,0,157,0,207,0,52,0,249,0,184,0,60,0,168,0,88,0,42,0,251,0,130,0,116,0);
signal scenario_full  : scenario_type := (0,0,135,31,135,30,127,31,127,30,127,29,21,31,101,31,175,31,186,31,85,31,153,31,153,30,221,31,136,31,133,31,221,31,68,31,178,31,35,31,164,31,87,31,87,30,87,29,22,31,241,31,241,30,139,31,72,31,228,31,238,31,102,31,11,31,55,31,55,30,109,31,55,31,55,30,99,31,243,31,219,31,119,31,133,31,5,31,89,31,197,31,181,31,19,31,220,31,46,31,198,31,198,30,226,31,79,31,160,31,79,31,205,31,107,31,1,31,210,31,17,31,196,31,165,31,205,31,31,31,69,31,142,31,158,31,192,31,192,30,220,31,186,31,234,31,24,31,24,30,127,31,252,31,45,31,45,30,53,31,116,31,182,31,141,31,208,31,224,31,115,31,60,31,127,31,247,31,210,31,170,31,233,31,233,30,100,31,100,30,167,31,6,31,170,31,254,31,221,31,221,30,65,31,65,30,209,31,242,31,119,31,203,31,248,31,121,31,121,30,155,31,120,31,126,31,197,31,203,31,203,30,17,31,68,31,68,30,147,31,162,31,133,31,210,31,211,31,68,31,231,31,86,31,158,31,152,31,201,31,164,31,15,31,15,30,59,31,101,31,38,31,182,31,56,31,128,31,128,30,91,31,121,31,246,31,246,30,246,29,109,31,168,31,168,30,205,31,64,31,189,31,123,31,21,31,223,31,200,31,200,30,7,31,199,31,175,31,159,31,159,30,189,31,220,31,28,31,23,31,23,30,34,31,253,31,120,31,217,31,217,30,187,31,21,31,167,31,116,31,116,30,32,31,32,30,82,31,91,31,91,30,230,31,86,31,114,31,104,31,186,31,211,31,20,31,103,31,23,31,130,31,222,31,224,31,35,31,78,31,154,31,172,31,178,31,100,31,100,30,235,31,240,31,240,30,109,31,220,31,144,31,91,31,242,31,242,30,200,31,85,31,85,30,85,29,135,31,135,30,135,29,70,31,229,31,121,31,121,30,63,31,208,31,208,30,208,29,46,31,101,31,241,31,163,31,199,31,18,31,156,31,34,31,16,31,247,31,177,31,86,31,220,31,204,31,10,31,39,31,25,31,46,31,87,31,39,31,161,31,63,31,63,30,137,31,160,31,154,31,191,31,129,31,59,31,59,30,24,31,54,31,221,31,183,31,116,31,193,31,193,30,193,29,93,31,59,31,59,30,135,31,215,31,212,31,4,31,4,30,4,29,207,31,207,30,142,31,142,30,120,31,124,31,48,31,180,31,105,31,33,31,4,31,208,31,179,31,117,31,159,31,70,31,70,30,19,31,247,31,209,31,90,31,216,31,127,31,127,30,64,31,64,30,202,31,38,31,67,31,105,31,105,30,105,29,105,28,105,27,194,31,114,31,181,31,213,31,229,31,230,31,230,30,30,31,75,31,37,31,81,31,225,31,19,31,147,31,11,31,11,30,176,31,29,31,29,30,29,29,195,31,195,30,219,31,167,31,7,31,219,31,251,31,235,31,103,31,30,31,113,31,249,31,202,31,116,31,103,31,65,31,21,31,236,31,236,30,236,29,175,31,117,31,162,31,10,31,246,31,123,31,209,31,229,31,3,31,171,31,202,31,166,31,189,31,3,31,50,31,190,31,250,31,119,31,119,30,238,31,92,31,104,31,242,31,87,31,236,31,236,30,236,29,62,31,228,31,228,30,179,31,77,31,156,31,58,31,117,31,117,30,58,31,218,31,218,30,138,31,123,31,102,31,119,31,94,31,117,31,34,31,30,31,158,31,158,30,40,31,40,30,40,29,197,31,197,30,31,31,136,31,102,31,141,31,158,31,158,30,93,31,110,31,212,31,114,31,114,30,190,31,87,31,2,31,76,31,250,31,175,31,57,31,57,30,55,31,23,31,40,31,112,31,146,31,251,31,230,31,37,31,234,31,228,31,34,31,17,31,112,31,154,31,247,31,56,31,58,31,96,31,204,31,2,31,137,31,143,31,143,30,248,31,248,30,140,31,110,31,26,31,26,30,26,29,26,28,112,31,112,30,218,31,196,31,196,30,56,31,225,31,73,31,128,31,236,31,236,30,189,31,167,31,167,30,167,29,230,31,236,31,221,31,87,31,38,31,38,30,38,29,251,31,79,31,79,30,220,31,187,31,187,30,44,31,28,31,206,31,45,31,82,31,82,30,106,31,106,30,44,31,102,31,119,31,207,31,215,31,208,31,31,31,158,31,131,31,30,31,99,31,52,31,222,31,157,31,157,30,157,29,157,28,147,31,128,31,185,31,177,31,110,31,119,31,224,31,146,31,236,31,21,31,235,31,243,31,199,31,173,31,121,31,121,30,90,31,216,31,174,31,155,31,102,31,25,31,196,31,242,31,45,31,45,30,122,31,36,31,22,31,168,31,235,31,220,31,212,31,110,31,139,31,112,31,112,30,27,31,96,31,87,31,87,30,79,31,206,31,150,31,249,31,198,31,226,31,117,31,30,31,5,31,60,31,60,30,101,31,201,31,148,31,55,31,235,31,177,31,91,31,25,31,162,31,194,31,118,31,13,31,6,31,47,31,47,30,18,31,237,31,150,31,149,31,172,31,90,31,8,31,8,30,115,31,223,31,232,31,232,30,123,31,143,31,195,31,239,31,95,31,95,30,92,31,67,31,32,31,32,30,88,31,57,31,175,31,82,31,79,31,214,31,152,31,50,31,50,30,150,31,44,31,40,31,224,31,223,31,155,31,245,31,38,31,79,31,17,31,183,31,222,31,33,31,33,30,168,31,127,31,127,30,166,31,205,31,198,31,150,31,202,31,237,31,237,30,145,31,111,31,40,31,4,31,4,30,4,29,183,31,107,31,221,31,221,30,38,31,38,30,38,29,86,31,5,31,82,31,82,30,33,31,157,31,33,31,158,31,196,31,196,30,196,29,136,31,232,31,232,30,232,29,208,31,208,30,30,31,12,31,20,31,183,31,179,31,37,31,37,30,99,31,99,30,99,29,67,31,112,31,112,30,112,29,75,31,68,31,210,31,137,31,137,30,137,29,77,31,247,31,186,31,89,31,89,30,234,31,234,30,10,31,100,31,181,31,139,31,158,31,134,31,251,31,226,31,86,31,236,31,141,31,85,31,6,31,129,31,229,31,57,31,121,31,121,30,121,29,121,28,41,31,134,31,235,31,40,31,40,30,44,31,44,30,115,31,106,31,61,31,112,31,142,31,252,31,1,31,1,30,187,31,37,31,37,30,35,31,209,31,108,31,133,31,168,31,168,30,75,31,147,31,116,31,122,31,166,31,26,31,251,31,41,31,26,31,180,31,84,31,191,31,206,31,208,31,131,31,188,31,69,31,235,31,75,31,150,31,100,31,145,31,110,31,110,30,110,29,41,31,139,31,176,31,201,31,97,31,102,31,109,31,161,31,161,30,147,31,28,31,33,31,148,31,180,31,33,31,134,31,127,31,155,31,55,31,55,30,23,31,92,31,83,31,183,31,208,31,56,31,244,31,119,31,153,31,158,31,127,31,127,30,192,31,53,31,171,31,171,30,37,31,13,31,170,31,135,31,190,31,190,30,156,31,110,31,245,31,124,31,164,31,12,31,51,31,41,31,132,31,86,31,86,30,201,31,128,31,32,31,32,30,9,31,80,31,163,31,42,31,92,31,223,31,207,31,66,31,247,31,66,31,19,31,19,30,241,31,14,31,153,31,233,31,220,31,163,31,163,30,221,31,154,31,234,31,169,31,115,31,110,31,196,31,196,30,73,31,83,31,68,31,96,31,96,30,60,31,110,31,227,31,227,30,124,31,133,31,58,31,253,31,139,31,71,31,151,31,19,31,121,31,119,31,96,31,96,30,166,31,71,31,134,31,193,31,193,30,93,31,226,31,173,31,173,30,131,31,183,31,158,31,246,31,9,31,9,30,83,31,238,31,238,30,24,31,211,31,69,31,69,30,206,31,183,31,172,31,85,31,150,31,16,31,220,31,7,31,60,31,1,31,145,31,84,31,205,31,192,31,24,31,1,31,112,31,111,31,115,31,17,31,95,31,155,31,128,31,128,30,33,31,162,31,114,31,90,31,36,31,5,31,5,30,15,31,173,31,110,31,228,31,86,31,86,30,198,31,55,31,87,31,87,30,91,31,137,31,176,31,52,31,224,31,91,31,210,31,236,31,74,31,103,31,39,31,49,31,160,31,64,31,100,31,100,30,120,31,110,31,110,30,63,31,68,31,49,31,236,31,12,31,12,30,12,29,11,31,11,30,116,31,157,31,207,31,52,31,249,31,184,31,60,31,168,31,88,31,42,31,251,31,130,31,116,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
