-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 597;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (138,0,0,0,153,0,197,0,59,0,0,0,93,0,28,0,0,0,55,0,18,0,216,0,0,0,0,0,66,0,143,0,38,0,137,0,0,0,0,0,212,0,0,0,178,0,222,0,80,0,252,0,0,0,71,0,236,0,121,0,22,0,177,0,0,0,97,0,28,0,228,0,141,0,143,0,152,0,230,0,52,0,0,0,53,0,211,0,12,0,242,0,46,0,62,0,250,0,78,0,0,0,0,0,177,0,184,0,146,0,17,0,137,0,13,0,90,0,12,0,0,0,148,0,164,0,126,0,65,0,43,0,94,0,132,0,231,0,28,0,0,0,201,0,23,0,137,0,237,0,42,0,51,0,29,0,250,0,98,0,115,0,0,0,127,0,43,0,0,0,0,0,198,0,107,0,115,0,146,0,235,0,8,0,221,0,0,0,115,0,77,0,225,0,0,0,179,0,156,0,213,0,0,0,93,0,127,0,232,0,93,0,0,0,0,0,0,0,0,0,0,0,37,0,40,0,45,0,0,0,103,0,0,0,222,0,218,0,102,0,0,0,122,0,187,0,0,0,152,0,89,0,48,0,233,0,198,0,42,0,0,0,0,0,32,0,0,0,23,0,78,0,201,0,158,0,239,0,70,0,4,0,0,0,235,0,143,0,122,0,78,0,141,0,109,0,121,0,52,0,183,0,63,0,150,0,115,0,150,0,140,0,221,0,4,0,233,0,238,0,209,0,129,0,56,0,0,0,219,0,82,0,17,0,160,0,34,0,44,0,78,0,254,0,216,0,228,0,0,0,0,0,245,0,0,0,185,0,42,0,234,0,0,0,15,0,0,0,224,0,2,0,0,0,20,0,232,0,56,0,150,0,95,0,24,0,189,0,154,0,126,0,51,0,68,0,0,0,0,0,107,0,177,0,0,0,44,0,181,0,0,0,225,0,0,0,0,0,252,0,122,0,174,0,96,0,151,0,57,0,72,0,155,0,87,0,167,0,25,0,228,0,78,0,115,0,0,0,0,0,9,0,40,0,114,0,81,0,180,0,254,0,91,0,151,0,98,0,8,0,148,0,97,0,157,0,125,0,105,0,165,0,246,0,199,0,89,0,131,0,124,0,3,0,163,0,116,0,110,0,205,0,241,0,251,0,164,0,131,0,18,0,0,0,229,0,85,0,196,0,0,0,26,0,34,0,0,0,49,0,133,0,212,0,78,0,14,0,26,0,154,0,167,0,132,0,173,0,0,0,196,0,44,0,25,0,213,0,247,0,18,0,112,0,232,0,0,0,0,0,135,0,245,0,23,0,90,0,90,0,51,0,183,0,133,0,163,0,0,0,0,0,39,0,213,0,0,0,198,0,181,0,70,0,0,0,17,0,58,0,106,0,255,0,202,0,17,0,71,0,251,0,0,0,121,0,153,0,124,0,27,0,0,0,0,0,165,0,171,0,233,0,0,0,45,0,196,0,240,0,0,0,0,0,0,0,0,0,193,0,65,0,70,0,105,0,130,0,187,0,162,0,208,0,130,0,36,0,144,0,37,0,178,0,239,0,0,0,77,0,0,0,143,0,211,0,10,0,0,0,0,0,103,0,0,0,194,0,100,0,110,0,106,0,245,0,232,0,147,0,3,0,6,0,0,0,0,0,20,0,187,0,106,0,193,0,2,0,240,0,198,0,172,0,48,0,109,0,242,0,232,0,159,0,80,0,22,0,51,0,236,0,33,0,251,0,0,0,180,0,239,0,105,0,196,0,0,0,0,0,247,0,45,0,122,0,83,0,35,0,0,0,181,0,193,0,91,0,27,0,241,0,73,0,0,0,181,0,210,0,88,0,60,0,23,0,96,0,78,0,136,0,0,0,115,0,98,0,237,0,95,0,0,0,244,0,130,0,106,0,32,0,0,0,82,0,85,0,20,0,0,0,81,0,242,0,91,0,0,0,0,0,92,0,0,0,165,0,115,0,123,0,202,0,123,0,122,0,142,0,0,0,71,0,0,0,110,0,232,0,0,0,59,0,239,0,171,0,195,0,95,0,10,0,158,0,131,0,146,0,0,0,131,0,50,0,38,0,0,0,0,0,246,0,0,0,117,0,102,0,53,0,252,0,0,0,31,0,40,0,192,0,32,0,202,0,192,0,20,0,0,0,180,0,10,0,125,0,207,0,249,0,0,0,73,0,0,0,140,0,107,0,198,0,0,0,63,0,110,0,113,0,10,0,39,0,250,0,0,0,104,0,90,0,218,0,141,0,21,0,47,0,0,0,35,0,160,0,211,0,53,0,77,0,52,0,241,0,193,0,165,0,202,0,183,0,202,0,115,0,149,0,134,0,207,0,91,0,82,0,240,0,0,0,74,0,90,0,195,0,63,0,26,0,42,0,0,0,13,0,24,0,84,0,0,0,102,0,104,0,0,0,96,0,135,0,53,0,196,0,0,0,0,0,93,0,255,0,54,0,247,0,101,0,127,0,0,0,210,0,194,0,0,0,0,0,216,0,21,0,60,0,29,0,0,0,108,0,232,0,65,0,243,0,31,0,156,0,0,0,52,0,252,0,156,0,3,0,0,0,162,0,49,0,195,0,182,0,245,0,252,0,57,0,20,0,163,0,215,0,0,0,20,0,113,0,0,0,55,0,0,0,49,0,19,0,200,0,125,0,0,0,149,0,39,0,93,0,116,0,52,0,198,0);
signal scenario_full  : scenario_type := (138,31,138,30,153,31,197,31,59,31,59,30,93,31,28,31,28,30,55,31,18,31,216,31,216,30,216,29,66,31,143,31,38,31,137,31,137,30,137,29,212,31,212,30,178,31,222,31,80,31,252,31,252,30,71,31,236,31,121,31,22,31,177,31,177,30,97,31,28,31,228,31,141,31,143,31,152,31,230,31,52,31,52,30,53,31,211,31,12,31,242,31,46,31,62,31,250,31,78,31,78,30,78,29,177,31,184,31,146,31,17,31,137,31,13,31,90,31,12,31,12,30,148,31,164,31,126,31,65,31,43,31,94,31,132,31,231,31,28,31,28,30,201,31,23,31,137,31,237,31,42,31,51,31,29,31,250,31,98,31,115,31,115,30,127,31,43,31,43,30,43,29,198,31,107,31,115,31,146,31,235,31,8,31,221,31,221,30,115,31,77,31,225,31,225,30,179,31,156,31,213,31,213,30,93,31,127,31,232,31,93,31,93,30,93,29,93,28,93,27,93,26,37,31,40,31,45,31,45,30,103,31,103,30,222,31,218,31,102,31,102,30,122,31,187,31,187,30,152,31,89,31,48,31,233,31,198,31,42,31,42,30,42,29,32,31,32,30,23,31,78,31,201,31,158,31,239,31,70,31,4,31,4,30,235,31,143,31,122,31,78,31,141,31,109,31,121,31,52,31,183,31,63,31,150,31,115,31,150,31,140,31,221,31,4,31,233,31,238,31,209,31,129,31,56,31,56,30,219,31,82,31,17,31,160,31,34,31,44,31,78,31,254,31,216,31,228,31,228,30,228,29,245,31,245,30,185,31,42,31,234,31,234,30,15,31,15,30,224,31,2,31,2,30,20,31,232,31,56,31,150,31,95,31,24,31,189,31,154,31,126,31,51,31,68,31,68,30,68,29,107,31,177,31,177,30,44,31,181,31,181,30,225,31,225,30,225,29,252,31,122,31,174,31,96,31,151,31,57,31,72,31,155,31,87,31,167,31,25,31,228,31,78,31,115,31,115,30,115,29,9,31,40,31,114,31,81,31,180,31,254,31,91,31,151,31,98,31,8,31,148,31,97,31,157,31,125,31,105,31,165,31,246,31,199,31,89,31,131,31,124,31,3,31,163,31,116,31,110,31,205,31,241,31,251,31,164,31,131,31,18,31,18,30,229,31,85,31,196,31,196,30,26,31,34,31,34,30,49,31,133,31,212,31,78,31,14,31,26,31,154,31,167,31,132,31,173,31,173,30,196,31,44,31,25,31,213,31,247,31,18,31,112,31,232,31,232,30,232,29,135,31,245,31,23,31,90,31,90,31,51,31,183,31,133,31,163,31,163,30,163,29,39,31,213,31,213,30,198,31,181,31,70,31,70,30,17,31,58,31,106,31,255,31,202,31,17,31,71,31,251,31,251,30,121,31,153,31,124,31,27,31,27,30,27,29,165,31,171,31,233,31,233,30,45,31,196,31,240,31,240,30,240,29,240,28,240,27,193,31,65,31,70,31,105,31,130,31,187,31,162,31,208,31,130,31,36,31,144,31,37,31,178,31,239,31,239,30,77,31,77,30,143,31,211,31,10,31,10,30,10,29,103,31,103,30,194,31,100,31,110,31,106,31,245,31,232,31,147,31,3,31,6,31,6,30,6,29,20,31,187,31,106,31,193,31,2,31,240,31,198,31,172,31,48,31,109,31,242,31,232,31,159,31,80,31,22,31,51,31,236,31,33,31,251,31,251,30,180,31,239,31,105,31,196,31,196,30,196,29,247,31,45,31,122,31,83,31,35,31,35,30,181,31,193,31,91,31,27,31,241,31,73,31,73,30,181,31,210,31,88,31,60,31,23,31,96,31,78,31,136,31,136,30,115,31,98,31,237,31,95,31,95,30,244,31,130,31,106,31,32,31,32,30,82,31,85,31,20,31,20,30,81,31,242,31,91,31,91,30,91,29,92,31,92,30,165,31,115,31,123,31,202,31,123,31,122,31,142,31,142,30,71,31,71,30,110,31,232,31,232,30,59,31,239,31,171,31,195,31,95,31,10,31,158,31,131,31,146,31,146,30,131,31,50,31,38,31,38,30,38,29,246,31,246,30,117,31,102,31,53,31,252,31,252,30,31,31,40,31,192,31,32,31,202,31,192,31,20,31,20,30,180,31,10,31,125,31,207,31,249,31,249,30,73,31,73,30,140,31,107,31,198,31,198,30,63,31,110,31,113,31,10,31,39,31,250,31,250,30,104,31,90,31,218,31,141,31,21,31,47,31,47,30,35,31,160,31,211,31,53,31,77,31,52,31,241,31,193,31,165,31,202,31,183,31,202,31,115,31,149,31,134,31,207,31,91,31,82,31,240,31,240,30,74,31,90,31,195,31,63,31,26,31,42,31,42,30,13,31,24,31,84,31,84,30,102,31,104,31,104,30,96,31,135,31,53,31,196,31,196,30,196,29,93,31,255,31,54,31,247,31,101,31,127,31,127,30,210,31,194,31,194,30,194,29,216,31,21,31,60,31,29,31,29,30,108,31,232,31,65,31,243,31,31,31,156,31,156,30,52,31,252,31,156,31,3,31,3,30,162,31,49,31,195,31,182,31,245,31,252,31,57,31,20,31,163,31,215,31,215,30,20,31,113,31,113,30,55,31,55,30,49,31,19,31,200,31,125,31,125,30,149,31,39,31,93,31,116,31,52,31,198,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
