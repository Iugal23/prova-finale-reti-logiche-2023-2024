-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_348 is
end project_tb_348;

architecture project_tb_arch_348 of project_tb_348 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 806;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (252,0,139,0,242,0,176,0,37,0,62,0,245,0,17,0,187,0,194,0,107,0,251,0,185,0,36,0,25,0,168,0,171,0,186,0,12,0,160,0,51,0,179,0,166,0,141,0,175,0,126,0,136,0,27,0,44,0,75,0,185,0,186,0,66,0,226,0,143,0,0,0,0,0,143,0,56,0,222,0,0,0,67,0,76,0,204,0,0,0,246,0,60,0,39,0,37,0,203,0,0,0,141,0,66,0,0,0,0,0,32,0,0,0,143,0,53,0,244,0,60,0,0,0,91,0,104,0,130,0,234,0,0,0,0,0,106,0,7,0,47,0,240,0,34,0,0,0,185,0,1,0,47,0,249,0,62,0,0,0,205,0,26,0,37,0,10,0,79,0,0,0,60,0,112,0,134,0,117,0,21,0,0,0,0,0,64,0,40,0,0,0,0,0,255,0,68,0,0,0,138,0,78,0,227,0,179,0,78,0,252,0,231,0,181,0,192,0,172,0,133,0,49,0,168,0,0,0,143,0,240,0,88,0,0,0,0,0,178,0,0,0,19,0,84,0,151,0,35,0,101,0,220,0,0,0,142,0,0,0,233,0,158,0,0,0,0,0,211,0,0,0,67,0,184,0,10,0,131,0,118,0,100,0,253,0,172,0,211,0,124,0,191,0,99,0,20,0,24,0,158,0,67,0,0,0,75,0,195,0,16,0,78,0,200,0,0,0,29,0,43,0,132,0,147,0,4,0,217,0,231,0,29,0,211,0,17,0,144,0,181,0,0,0,0,0,0,0,6,0,134,0,0,0,192,0,175,0,102,0,200,0,151,0,15,0,55,0,232,0,204,0,81,0,0,0,27,0,191,0,233,0,165,0,84,0,0,0,62,0,163,0,0,0,5,0,211,0,103,0,200,0,0,0,0,0,31,0,153,0,121,0,234,0,8,0,0,0,242,0,150,0,37,0,209,0,110,0,134,0,0,0,86,0,251,0,242,0,240,0,188,0,198,0,0,0,211,0,0,0,0,0,0,0,224,0,213,0,131,0,66,0,45,0,161,0,184,0,222,0,96,0,30,0,100,0,254,0,146,0,139,0,166,0,197,0,0,0,0,0,54,0,117,0,3,0,85,0,60,0,7,0,189,0,0,0,0,0,121,0,185,0,0,0,0,0,187,0,118,0,156,0,161,0,0,0,104,0,72,0,160,0,181,0,0,0,70,0,181,0,193,0,32,0,146,0,35,0,55,0,0,0,127,0,46,0,0,0,1,0,0,0,198,0,125,0,68,0,0,0,188,0,206,0,139,0,68,0,139,0,20,0,112,0,0,0,156,0,247,0,0,0,0,0,105,0,55,0,217,0,0,0,251,0,116,0,213,0,107,0,11,0,0,0,34,0,71,0,66,0,24,0,124,0,65,0,40,0,233,0,0,0,171,0,254,0,203,0,175,0,0,0,232,0,238,0,3,0,158,0,167,0,0,0,47,0,157,0,52,0,39,0,112,0,220,0,0,0,241,0,18,0,52,0,210,0,67,0,13,0,0,0,0,0,0,0,198,0,0,0,134,0,192,0,36,0,0,0,251,0,94,0,222,0,0,0,57,0,171,0,208,0,27,0,160,0,244,0,106,0,61,0,155,0,44,0,72,0,228,0,0,0,79,0,41,0,10,0,155,0,0,0,0,0,72,0,0,0,167,0,240,0,139,0,105,0,3,0,90,0,0,0,115,0,200,0,60,0,0,0,162,0,188,0,165,0,0,0,71,0,9,0,108,0,0,0,111,0,216,0,43,0,190,0,0,0,84,0,168,0,101,0,242,0,0,0,6,0,52,0,60,0,102,0,207,0,63,0,49,0,0,0,171,0,91,0,165,0,188,0,106,0,211,0,109,0,245,0,228,0,190,0,0,0,133,0,241,0,9,0,241,0,0,0,0,0,0,0,204,0,45,0,50,0,237,0,237,0,32,0,72,0,250,0,186,0,107,0,122,0,6,0,21,0,71,0,0,0,82,0,27,0,203,0,240,0,57,0,0,0,238,0,0,0,20,0,83,0,0,0,5,0,0,0,181,0,20,0,56,0,193,0,29,0,166,0,117,0,219,0,0,0,156,0,0,0,0,0,0,0,139,0,248,0,61,0,0,0,130,0,104,0,153,0,0,0,43,0,143,0,243,0,84,0,10,0,42,0,98,0,0,0,98,0,103,0,46,0,96,0,159,0,211,0,240,0,177,0,139,0,142,0,225,0,0,0,234,0,0,0,252,0,205,0,119,0,183,0,186,0,190,0,0,0,119,0,0,0,155,0,19,0,8,0,132,0,60,0,152,0,0,0,14,0,162,0,0,0,0,0,48,0,0,0,0,0,0,0,127,0,43,0,79,0,85,0,106,0,67,0,249,0,0,0,0,0,140,0,157,0,57,0,0,0,154,0,247,0,80,0,0,0,133,0,0,0,0,0,111,0,62,0,29,0,191,0,0,0,30,0,185,0,21,0,0,0,214,0,39,0,1,0,57,0,198,0,116,0,161,0,37,0,133,0,251,0,237,0,0,0,238,0,0,0,235,0,251,0,0,0,6,0,154,0,241,0,90,0,81,0,153,0,207,0,185,0,3,0,27,0,28,0,101,0,0,0,64,0,246,0,142,0,0,0,4,0,12,0,251,0,59,0,229,0,210,0,169,0,21,0,159,0,222,0,10,0,26,0,30,0,133,0,0,0,154,0,225,0,108,0,0,0,94,0,171,0,53,0,249,0,32,0,88,0,234,0,57,0,55,0,0,0,38,0,197,0,212,0,248,0,245,0,104,0,220,0,128,0,51,0,109,0,218,0,21,0,121,0,157,0,108,0,215,0,94,0,251,0,166,0,22,0,0,0,53,0,0,0,163,0,17,0,32,0,79,0,0,0,0,0,129,0,0,0,88,0,33,0,13,0,3,0,170,0,59,0,0,0,120,0,41,0,213,0,85,0,0,0,11,0,137,0,246,0,164,0,205,0,35,0,237,0,240,0,3,0,200,0,56,0,238,0,245,0,0,0,162,0,234,0,218,0,247,0,209,0,230,0,0,0,21,0,0,0,219,0,44,0,241,0,188,0,28,0,10,0,132,0,47,0,104,0,236,0,48,0,7,0,202,0,162,0,0,0,0,0,147,0,247,0,131,0,17,0,0,0,188,0,87,0,0,0,122,0,31,0,7,0,110,0,109,0,96,0,253,0,240,0,185,0,96,0,0,0,116,0,0,0,210,0,172,0,246,0,95,0,248,0,32,0,4,0,248,0,0,0,128,0,85,0,0,0,176,0,0,0,70,0,0,0,187,0,9,0,49,0,0,0,157,0,41,0,0,0,116,0,29,0,115,0,187,0,34,0,101,0,0,0,68,0,0,0,81,0,204,0,8,0,0,0,181,0,43,0,130,0,151,0,102,0,167,0,190,0,36,0,111,0,100,0,114,0,255,0,14,0,95,0,0,0,206,0,44,0,111,0,86,0,0,0,215,0,169,0,123,0,193,0,3,0,215,0,15,0,0,0,0,0,0,0,38,0,0,0,122,0,69,0,69,0,149,0,113,0,64,0,145,0,98,0,168,0,0,0,53,0,88,0,15,0,0,0,8,0,69,0,0,0,114,0,175,0);
signal scenario_full  : scenario_type := (252,31,139,31,242,31,176,31,37,31,62,31,245,31,17,31,187,31,194,31,107,31,251,31,185,31,36,31,25,31,168,31,171,31,186,31,12,31,160,31,51,31,179,31,166,31,141,31,175,31,126,31,136,31,27,31,44,31,75,31,185,31,186,31,66,31,226,31,143,31,143,30,143,29,143,31,56,31,222,31,222,30,67,31,76,31,204,31,204,30,246,31,60,31,39,31,37,31,203,31,203,30,141,31,66,31,66,30,66,29,32,31,32,30,143,31,53,31,244,31,60,31,60,30,91,31,104,31,130,31,234,31,234,30,234,29,106,31,7,31,47,31,240,31,34,31,34,30,185,31,1,31,47,31,249,31,62,31,62,30,205,31,26,31,37,31,10,31,79,31,79,30,60,31,112,31,134,31,117,31,21,31,21,30,21,29,64,31,40,31,40,30,40,29,255,31,68,31,68,30,138,31,78,31,227,31,179,31,78,31,252,31,231,31,181,31,192,31,172,31,133,31,49,31,168,31,168,30,143,31,240,31,88,31,88,30,88,29,178,31,178,30,19,31,84,31,151,31,35,31,101,31,220,31,220,30,142,31,142,30,233,31,158,31,158,30,158,29,211,31,211,30,67,31,184,31,10,31,131,31,118,31,100,31,253,31,172,31,211,31,124,31,191,31,99,31,20,31,24,31,158,31,67,31,67,30,75,31,195,31,16,31,78,31,200,31,200,30,29,31,43,31,132,31,147,31,4,31,217,31,231,31,29,31,211,31,17,31,144,31,181,31,181,30,181,29,181,28,6,31,134,31,134,30,192,31,175,31,102,31,200,31,151,31,15,31,55,31,232,31,204,31,81,31,81,30,27,31,191,31,233,31,165,31,84,31,84,30,62,31,163,31,163,30,5,31,211,31,103,31,200,31,200,30,200,29,31,31,153,31,121,31,234,31,8,31,8,30,242,31,150,31,37,31,209,31,110,31,134,31,134,30,86,31,251,31,242,31,240,31,188,31,198,31,198,30,211,31,211,30,211,29,211,28,224,31,213,31,131,31,66,31,45,31,161,31,184,31,222,31,96,31,30,31,100,31,254,31,146,31,139,31,166,31,197,31,197,30,197,29,54,31,117,31,3,31,85,31,60,31,7,31,189,31,189,30,189,29,121,31,185,31,185,30,185,29,187,31,118,31,156,31,161,31,161,30,104,31,72,31,160,31,181,31,181,30,70,31,181,31,193,31,32,31,146,31,35,31,55,31,55,30,127,31,46,31,46,30,1,31,1,30,198,31,125,31,68,31,68,30,188,31,206,31,139,31,68,31,139,31,20,31,112,31,112,30,156,31,247,31,247,30,247,29,105,31,55,31,217,31,217,30,251,31,116,31,213,31,107,31,11,31,11,30,34,31,71,31,66,31,24,31,124,31,65,31,40,31,233,31,233,30,171,31,254,31,203,31,175,31,175,30,232,31,238,31,3,31,158,31,167,31,167,30,47,31,157,31,52,31,39,31,112,31,220,31,220,30,241,31,18,31,52,31,210,31,67,31,13,31,13,30,13,29,13,28,198,31,198,30,134,31,192,31,36,31,36,30,251,31,94,31,222,31,222,30,57,31,171,31,208,31,27,31,160,31,244,31,106,31,61,31,155,31,44,31,72,31,228,31,228,30,79,31,41,31,10,31,155,31,155,30,155,29,72,31,72,30,167,31,240,31,139,31,105,31,3,31,90,31,90,30,115,31,200,31,60,31,60,30,162,31,188,31,165,31,165,30,71,31,9,31,108,31,108,30,111,31,216,31,43,31,190,31,190,30,84,31,168,31,101,31,242,31,242,30,6,31,52,31,60,31,102,31,207,31,63,31,49,31,49,30,171,31,91,31,165,31,188,31,106,31,211,31,109,31,245,31,228,31,190,31,190,30,133,31,241,31,9,31,241,31,241,30,241,29,241,28,204,31,45,31,50,31,237,31,237,31,32,31,72,31,250,31,186,31,107,31,122,31,6,31,21,31,71,31,71,30,82,31,27,31,203,31,240,31,57,31,57,30,238,31,238,30,20,31,83,31,83,30,5,31,5,30,181,31,20,31,56,31,193,31,29,31,166,31,117,31,219,31,219,30,156,31,156,30,156,29,156,28,139,31,248,31,61,31,61,30,130,31,104,31,153,31,153,30,43,31,143,31,243,31,84,31,10,31,42,31,98,31,98,30,98,31,103,31,46,31,96,31,159,31,211,31,240,31,177,31,139,31,142,31,225,31,225,30,234,31,234,30,252,31,205,31,119,31,183,31,186,31,190,31,190,30,119,31,119,30,155,31,19,31,8,31,132,31,60,31,152,31,152,30,14,31,162,31,162,30,162,29,48,31,48,30,48,29,48,28,127,31,43,31,79,31,85,31,106,31,67,31,249,31,249,30,249,29,140,31,157,31,57,31,57,30,154,31,247,31,80,31,80,30,133,31,133,30,133,29,111,31,62,31,29,31,191,31,191,30,30,31,185,31,21,31,21,30,214,31,39,31,1,31,57,31,198,31,116,31,161,31,37,31,133,31,251,31,237,31,237,30,238,31,238,30,235,31,251,31,251,30,6,31,154,31,241,31,90,31,81,31,153,31,207,31,185,31,3,31,27,31,28,31,101,31,101,30,64,31,246,31,142,31,142,30,4,31,12,31,251,31,59,31,229,31,210,31,169,31,21,31,159,31,222,31,10,31,26,31,30,31,133,31,133,30,154,31,225,31,108,31,108,30,94,31,171,31,53,31,249,31,32,31,88,31,234,31,57,31,55,31,55,30,38,31,197,31,212,31,248,31,245,31,104,31,220,31,128,31,51,31,109,31,218,31,21,31,121,31,157,31,108,31,215,31,94,31,251,31,166,31,22,31,22,30,53,31,53,30,163,31,17,31,32,31,79,31,79,30,79,29,129,31,129,30,88,31,33,31,13,31,3,31,170,31,59,31,59,30,120,31,41,31,213,31,85,31,85,30,11,31,137,31,246,31,164,31,205,31,35,31,237,31,240,31,3,31,200,31,56,31,238,31,245,31,245,30,162,31,234,31,218,31,247,31,209,31,230,31,230,30,21,31,21,30,219,31,44,31,241,31,188,31,28,31,10,31,132,31,47,31,104,31,236,31,48,31,7,31,202,31,162,31,162,30,162,29,147,31,247,31,131,31,17,31,17,30,188,31,87,31,87,30,122,31,31,31,7,31,110,31,109,31,96,31,253,31,240,31,185,31,96,31,96,30,116,31,116,30,210,31,172,31,246,31,95,31,248,31,32,31,4,31,248,31,248,30,128,31,85,31,85,30,176,31,176,30,70,31,70,30,187,31,9,31,49,31,49,30,157,31,41,31,41,30,116,31,29,31,115,31,187,31,34,31,101,31,101,30,68,31,68,30,81,31,204,31,8,31,8,30,181,31,43,31,130,31,151,31,102,31,167,31,190,31,36,31,111,31,100,31,114,31,255,31,14,31,95,31,95,30,206,31,44,31,111,31,86,31,86,30,215,31,169,31,123,31,193,31,3,31,215,31,15,31,15,30,15,29,15,28,38,31,38,30,122,31,69,31,69,31,149,31,113,31,64,31,145,31,98,31,168,31,168,30,53,31,88,31,15,31,15,30,8,31,69,31,69,30,114,31,175,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
