-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 632;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (114,0,53,0,6,0,0,0,195,0,152,0,36,0,215,0,0,0,0,0,0,0,112,0,0,0,61,0,20,0,95,0,86,0,83,0,46,0,0,0,222,0,205,0,254,0,0,0,232,0,63,0,102,0,0,0,57,0,171,0,249,0,184,0,0,0,196,0,190,0,68,0,29,0,47,0,35,0,187,0,94,0,0,0,215,0,23,0,238,0,135,0,65,0,62,0,30,0,0,0,0,0,0,0,79,0,150,0,0,0,16,0,133,0,78,0,64,0,89,0,0,0,107,0,36,0,92,0,181,0,0,0,0,0,214,0,185,0,67,0,120,0,109,0,17,0,105,0,86,0,53,0,158,0,124,0,241,0,113,0,89,0,0,0,42,0,119,0,232,0,0,0,155,0,137,0,134,0,0,0,251,0,0,0,91,0,59,0,164,0,180,0,8,0,63,0,185,0,83,0,1,0,59,0,0,0,0,0,0,0,37,0,242,0,207,0,254,0,159,0,195,0,0,0,150,0,16,0,167,0,125,0,104,0,158,0,158,0,181,0,49,0,164,0,206,0,16,0,0,0,168,0,0,0,154,0,0,0,193,0,5,0,149,0,190,0,89,0,244,0,62,0,65,0,84,0,39,0,24,0,70,0,117,0,178,0,55,0,0,0,59,0,205,0,108,0,173,0,120,0,25,0,0,0,209,0,53,0,130,0,0,0,214,0,0,0,169,0,154,0,125,0,5,0,38,0,45,0,234,0,97,0,109,0,179,0,170,0,153,0,65,0,199,0,44,0,0,0,223,0,122,0,0,0,182,0,23,0,158,0,29,0,0,0,168,0,73,0,81,0,255,0,108,0,182,0,146,0,167,0,242,0,85,0,105,0,52,0,180,0,0,0,99,0,183,0,227,0,178,0,56,0,0,0,22,0,30,0,165,0,31,0,236,0,127,0,19,0,0,0,23,0,0,0,0,0,164,0,29,0,0,0,141,0,63,0,22,0,150,0,37,0,127,0,67,0,238,0,165,0,175,0,152,0,7,0,57,0,183,0,0,0,0,0,114,0,225,0,0,0,231,0,188,0,191,0,169,0,113,0,0,0,193,0,21,0,182,0,178,0,0,0,149,0,189,0,0,0,90,0,214,0,0,0,0,0,212,0,240,0,0,0,243,0,219,0,124,0,177,0,142,0,144,0,0,0,240,0,113,0,53,0,71,0,48,0,239,0,110,0,0,0,245,0,225,0,44,0,192,0,203,0,19,0,0,0,89,0,99,0,216,0,4,0,100,0,0,0,0,0,119,0,254,0,45,0,128,0,0,0,151,0,0,0,138,0,162,0,0,0,212,0,213,0,97,0,104,0,139,0,124,0,77,0,163,0,0,0,25,0,0,0,189,0,12,0,5,0,5,0,0,0,237,0,218,0,194,0,7,0,237,0,64,0,196,0,0,0,64,0,59,0,71,0,34,0,0,0,0,0,28,0,125,0,92,0,128,0,164,0,0,0,40,0,130,0,57,0,242,0,230,0,185,0,97,0,121,0,218,0,77,0,0,0,0,0,213,0,50,0,181,0,224,0,0,0,157,0,201,0,239,0,0,0,154,0,0,0,156,0,160,0,82,0,66,0,117,0,15,0,0,0,0,0,0,0,0,0,137,0,178,0,41,0,0,0,210,0,123,0,240,0,137,0,3,0,49,0,101,0,0,0,10,0,93,0,250,0,232,0,24,0,217,0,149,0,0,0,0,0,182,0,91,0,229,0,98,0,242,0,82,0,40,0,220,0,72,0,138,0,237,0,151,0,201,0,113,0,0,0,0,0,244,0,59,0,28,0,99,0,0,0,72,0,192,0,110,0,147,0,0,0,0,0,170,0,32,0,0,0,42,0,91,0,40,0,206,0,90,0,88,0,6,0,27,0,0,0,89,0,0,0,91,0,92,0,212,0,6,0,0,0,0,0,116,0,207,0,213,0,0,0,237,0,42,0,0,0,93,0,94,0,190,0,38,0,98,0,0,0,105,0,0,0,106,0,29,0,206,0,253,0,186,0,96,0,117,0,0,0,129,0,58,0,51,0,201,0,0,0,52,0,240,0,180,0,243,0,158,0,252,0,221,0,87,0,0,0,174,0,0,0,251,0,107,0,18,0,40,0,108,0,176,0,40,0,24,0,89,0,0,0,29,0,254,0,184,0,103,0,111,0,84,0,0,0,0,0,217,0,44,0,166,0,164,0,5,0,79,0,26,0,122,0,195,0,43,0,0,0,79,0,188,0,155,0,207,0,34,0,27,0,208,0,246,0,245,0,34,0,206,0,66,0,208,0,240,0,144,0,0,0,194,0,142,0,0,0,156,0,169,0,0,0,128,0,0,0,197,0,163,0,157,0,0,0,0,0,124,0,227,0,105,0,45,0,175,0,15,0,135,0,228,0,123,0,161,0,65,0,0,0,92,0,0,0,0,0,238,0,202,0,127,0,23,0,202,0,61,0,237,0,78,0,236,0,160,0,153,0,242,0,238,0,21,0,108,0,0,0,182,0,173,0,173,0,0,0,229,0,217,0,89,0,189,0,0,0,58,0,132,0,30,0,108,0,0,0,202,0,42,0,217,0,165,0,0,0,19,0,185,0,0,0,129,0,198,0,80,0,192,0,254,0,220,0,0,0,179,0,128,0,57,0,146,0,33,0,106,0,4,0,180,0,0,0,99,0,219,0,121,0,180,0,105,0,41,0,75,0,159,0,142,0,164,0,79,0,65,0,24,0,0,0,94,0,57,0,0,0,0,0,195,0,144,0,90,0,18,0,0,0,101,0,9,0,229,0,0,0,50,0,97,0,129,0,244,0,48,0,145,0,185,0);
signal scenario_full  : scenario_type := (114,31,53,31,6,31,6,30,195,31,152,31,36,31,215,31,215,30,215,29,215,28,112,31,112,30,61,31,20,31,95,31,86,31,83,31,46,31,46,30,222,31,205,31,254,31,254,30,232,31,63,31,102,31,102,30,57,31,171,31,249,31,184,31,184,30,196,31,190,31,68,31,29,31,47,31,35,31,187,31,94,31,94,30,215,31,23,31,238,31,135,31,65,31,62,31,30,31,30,30,30,29,30,28,79,31,150,31,150,30,16,31,133,31,78,31,64,31,89,31,89,30,107,31,36,31,92,31,181,31,181,30,181,29,214,31,185,31,67,31,120,31,109,31,17,31,105,31,86,31,53,31,158,31,124,31,241,31,113,31,89,31,89,30,42,31,119,31,232,31,232,30,155,31,137,31,134,31,134,30,251,31,251,30,91,31,59,31,164,31,180,31,8,31,63,31,185,31,83,31,1,31,59,31,59,30,59,29,59,28,37,31,242,31,207,31,254,31,159,31,195,31,195,30,150,31,16,31,167,31,125,31,104,31,158,31,158,31,181,31,49,31,164,31,206,31,16,31,16,30,168,31,168,30,154,31,154,30,193,31,5,31,149,31,190,31,89,31,244,31,62,31,65,31,84,31,39,31,24,31,70,31,117,31,178,31,55,31,55,30,59,31,205,31,108,31,173,31,120,31,25,31,25,30,209,31,53,31,130,31,130,30,214,31,214,30,169,31,154,31,125,31,5,31,38,31,45,31,234,31,97,31,109,31,179,31,170,31,153,31,65,31,199,31,44,31,44,30,223,31,122,31,122,30,182,31,23,31,158,31,29,31,29,30,168,31,73,31,81,31,255,31,108,31,182,31,146,31,167,31,242,31,85,31,105,31,52,31,180,31,180,30,99,31,183,31,227,31,178,31,56,31,56,30,22,31,30,31,165,31,31,31,236,31,127,31,19,31,19,30,23,31,23,30,23,29,164,31,29,31,29,30,141,31,63,31,22,31,150,31,37,31,127,31,67,31,238,31,165,31,175,31,152,31,7,31,57,31,183,31,183,30,183,29,114,31,225,31,225,30,231,31,188,31,191,31,169,31,113,31,113,30,193,31,21,31,182,31,178,31,178,30,149,31,189,31,189,30,90,31,214,31,214,30,214,29,212,31,240,31,240,30,243,31,219,31,124,31,177,31,142,31,144,31,144,30,240,31,113,31,53,31,71,31,48,31,239,31,110,31,110,30,245,31,225,31,44,31,192,31,203,31,19,31,19,30,89,31,99,31,216,31,4,31,100,31,100,30,100,29,119,31,254,31,45,31,128,31,128,30,151,31,151,30,138,31,162,31,162,30,212,31,213,31,97,31,104,31,139,31,124,31,77,31,163,31,163,30,25,31,25,30,189,31,12,31,5,31,5,31,5,30,237,31,218,31,194,31,7,31,237,31,64,31,196,31,196,30,64,31,59,31,71,31,34,31,34,30,34,29,28,31,125,31,92,31,128,31,164,31,164,30,40,31,130,31,57,31,242,31,230,31,185,31,97,31,121,31,218,31,77,31,77,30,77,29,213,31,50,31,181,31,224,31,224,30,157,31,201,31,239,31,239,30,154,31,154,30,156,31,160,31,82,31,66,31,117,31,15,31,15,30,15,29,15,28,15,27,137,31,178,31,41,31,41,30,210,31,123,31,240,31,137,31,3,31,49,31,101,31,101,30,10,31,93,31,250,31,232,31,24,31,217,31,149,31,149,30,149,29,182,31,91,31,229,31,98,31,242,31,82,31,40,31,220,31,72,31,138,31,237,31,151,31,201,31,113,31,113,30,113,29,244,31,59,31,28,31,99,31,99,30,72,31,192,31,110,31,147,31,147,30,147,29,170,31,32,31,32,30,42,31,91,31,40,31,206,31,90,31,88,31,6,31,27,31,27,30,89,31,89,30,91,31,92,31,212,31,6,31,6,30,6,29,116,31,207,31,213,31,213,30,237,31,42,31,42,30,93,31,94,31,190,31,38,31,98,31,98,30,105,31,105,30,106,31,29,31,206,31,253,31,186,31,96,31,117,31,117,30,129,31,58,31,51,31,201,31,201,30,52,31,240,31,180,31,243,31,158,31,252,31,221,31,87,31,87,30,174,31,174,30,251,31,107,31,18,31,40,31,108,31,176,31,40,31,24,31,89,31,89,30,29,31,254,31,184,31,103,31,111,31,84,31,84,30,84,29,217,31,44,31,166,31,164,31,5,31,79,31,26,31,122,31,195,31,43,31,43,30,79,31,188,31,155,31,207,31,34,31,27,31,208,31,246,31,245,31,34,31,206,31,66,31,208,31,240,31,144,31,144,30,194,31,142,31,142,30,156,31,169,31,169,30,128,31,128,30,197,31,163,31,157,31,157,30,157,29,124,31,227,31,105,31,45,31,175,31,15,31,135,31,228,31,123,31,161,31,65,31,65,30,92,31,92,30,92,29,238,31,202,31,127,31,23,31,202,31,61,31,237,31,78,31,236,31,160,31,153,31,242,31,238,31,21,31,108,31,108,30,182,31,173,31,173,31,173,30,229,31,217,31,89,31,189,31,189,30,58,31,132,31,30,31,108,31,108,30,202,31,42,31,217,31,165,31,165,30,19,31,185,31,185,30,129,31,198,31,80,31,192,31,254,31,220,31,220,30,179,31,128,31,57,31,146,31,33,31,106,31,4,31,180,31,180,30,99,31,219,31,121,31,180,31,105,31,41,31,75,31,159,31,142,31,164,31,79,31,65,31,24,31,24,30,94,31,57,31,57,30,57,29,195,31,144,31,90,31,18,31,18,30,101,31,9,31,229,31,229,30,50,31,97,31,129,31,244,31,48,31,145,31,185,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
