-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_929 is
end project_tb_929;

architecture project_tb_arch_929 of project_tb_929 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 781;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (134,0,129,0,0,0,143,0,79,0,31,0,246,0,59,0,0,0,217,0,183,0,103,0,24,0,217,0,0,0,0,0,158,0,0,0,72,0,0,0,247,0,146,0,0,0,109,0,0,0,8,0,3,0,0,0,181,0,181,0,78,0,208,0,140,0,235,0,140,0,24,0,166,0,0,0,137,0,232,0,63,0,117,0,118,0,87,0,134,0,168,0,147,0,0,0,43,0,16,0,84,0,86,0,127,0,137,0,0,0,95,0,128,0,75,0,40,0,129,0,189,0,111,0,0,0,133,0,65,0,71,0,138,0,237,0,66,0,171,0,202,0,244,0,198,0,182,0,74,0,160,0,10,0,194,0,0,0,100,0,153,0,0,0,81,0,0,0,137,0,189,0,77,0,101,0,196,0,132,0,0,0,91,0,34,0,139,0,213,0,0,0,235,0,0,0,136,0,163,0,228,0,66,0,212,0,201,0,139,0,232,0,14,0,218,0,189,0,0,0,21,0,212,0,0,0,0,0,224,0,21,0,169,0,148,0,0,0,112,0,250,0,0,0,185,0,0,0,10,0,72,0,234,0,112,0,45,0,124,0,141,0,112,0,248,0,88,0,0,0,180,0,0,0,156,0,143,0,10,0,29,0,129,0,0,0,23,0,64,0,0,0,225,0,170,0,0,0,70,0,59,0,203,0,236,0,0,0,0,0,0,0,217,0,101,0,10,0,109,0,0,0,0,0,196,0,240,0,223,0,80,0,1,0,0,0,5,0,0,0,100,0,127,0,224,0,69,0,40,0,0,0,181,0,0,0,79,0,173,0,242,0,111,0,115,0,144,0,114,0,28,0,0,0,31,0,11,0,2,0,27,0,88,0,0,0,162,0,124,0,58,0,50,0,179,0,20,0,93,0,209,0,117,0,142,0,188,0,11,0,71,0,190,0,0,0,172,0,134,0,103,0,247,0,58,0,45,0,22,0,219,0,167,0,208,0,0,0,159,0,252,0,134,0,124,0,194,0,14,0,241,0,247,0,253,0,134,0,87,0,251,0,0,0,0,0,0,0,36,0,36,0,0,0,212,0,77,0,196,0,210,0,29,0,8,0,0,0,131,0,131,0,210,0,187,0,172,0,109,0,124,0,0,0,134,0,154,0,16,0,127,0,51,0,85,0,217,0,0,0,203,0,16,0,111,0,238,0,19,0,44,0,75,0,0,0,0,0,128,0,181,0,226,0,21,0,0,0,186,0,153,0,144,0,0,0,46,0,0,0,69,0,202,0,0,0,136,0,234,0,40,0,106,0,54,0,116,0,0,0,35,0,202,0,39,0,222,0,132,0,77,0,119,0,4,0,25,0,154,0,112,0,89,0,4,0,198,0,84,0,78,0,249,0,51,0,167,0,116,0,101,0,161,0,146,0,152,0,0,0,80,0,0,0,52,0,76,0,32,0,147,0,228,0,5,0,190,0,228,0,34,0,8,0,114,0,0,0,147,0,209,0,0,0,151,0,30,0,0,0,32,0,126,0,148,0,0,0,232,0,33,0,71,0,17,0,197,0,131,0,36,0,149,0,95,0,210,0,78,0,0,0,206,0,245,0,103,0,40,0,104,0,0,0,107,0,251,0,0,0,255,0,223,0,126,0,28,0,232,0,0,0,0,0,78,0,245,0,255,0,128,0,0,0,193,0,111,0,177,0,0,0,31,0,56,0,231,0,189,0,210,0,158,0,23,0,16,0,0,0,106,0,42,0,46,0,193,0,81,0,153,0,200,0,0,0,19,0,247,0,114,0,137,0,190,0,0,0,160,0,31,0,2,0,114,0,47,0,200,0,155,0,0,0,101,0,206,0,0,0,107,0,0,0,216,0,187,0,73,0,31,0,0,0,227,0,153,0,117,0,239,0,247,0,106,0,180,0,88,0,0,0,24,0,107,0,75,0,220,0,0,0,90,0,242,0,80,0,163,0,152,0,147,0,36,0,0,0,85,0,0,0,151,0,0,0,27,0,108,0,186,0,108,0,0,0,63,0,248,0,85,0,164,0,242,0,23,0,0,0,0,0,75,0,172,0,0,0,0,0,184,0,211,0,116,0,109,0,202,0,154,0,21,0,0,0,254,0,67,0,169,0,172,0,125,0,152,0,61,0,124,0,0,0,199,0,224,0,0,0,237,0,189,0,0,0,0,0,129,0,66,0,199,0,129,0,0,0,68,0,0,0,171,0,153,0,192,0,0,0,176,0,126,0,73,0,57,0,0,0,215,0,192,0,164,0,169,0,231,0,146,0,175,0,155,0,249,0,41,0,0,0,9,0,54,0,105,0,56,0,152,0,252,0,0,0,208,0,134,0,120,0,47,0,230,0,0,0,26,0,248,0,72,0,211,0,0,0,105,0,171,0,224,0,20,0,112,0,200,0,0,0,162,0,55,0,0,0,35,0,16,0,66,0,68,0,5,0,54,0,120,0,96,0,67,0,125,0,237,0,88,0,27,0,229,0,172,0,147,0,200,0,251,0,0,0,6,0,240,0,230,0,141,0,132,0,194,0,30,0,159,0,0,0,0,0,67,0,6,0,131,0,28,0,38,0,51,0,109,0,229,0,197,0,66,0,27,0,5,0,0,0,179,0,3,0,0,0,209,0,0,0,0,0,197,0,86,0,114,0,144,0,196,0,171,0,248,0,50,0,0,0,134,0,36,0,171,0,5,0,228,0,161,0,98,0,0,0,99,0,0,0,0,0,0,0,0,0,52,0,174,0,141,0,100,0,1,0,83,0,0,0,0,0,5,0,77,0,50,0,16,0,50,0,40,0,100,0,90,0,165,0,250,0,35,0,0,0,0,0,38,0,41,0,0,0,34,0,239,0,130,0,79,0,136,0,0,0,25,0,183,0,244,0,236,0,83,0,0,0,162,0,0,0,172,0,177,0,0,0,43,0,20,0,44,0,0,0,245,0,181,0,121,0,191,0,219,0,222,0,85,0,156,0,248,0,0,0,0,0,28,0,136,0,167,0,41,0,211,0,141,0,65,0,81,0,9,0,233,0,0,0,26,0,109,0,36,0,112,0,0,0,2,0,98,0,94,0,89,0,115,0,127,0,191,0,204,0,220,0,14,0,236,0,0,0,159,0,204,0,177,0,116,0,226,0,0,0,134,0,74,0,178,0,211,0,175,0,100,0,191,0,0,0,0,0,0,0,0,0,200,0,239,0,1,0,0,0,223,0,74,0,226,0,77,0,225,0,0,0,82,0,0,0,86,0,154,0,242,0,40,0,138,0,0,0,119,0,223,0,3,0,90,0,97,0,14,0,125,0,12,0,5,0,0,0,222,0,1,0,16,0,180,0,207,0,95,0,118,0,0,0,60,0,164,0,0,0,0,0,40,0,196,0,77,0,29,0,1,0,230,0,141,0,0,0,0,0,108,0,57,0,118,0,199,0,237,0,127,0,0,0,79,0,0,0,0,0,249,0,170,0,2,0,87,0,0,0,59,0,0,0,209,0,0,0,202,0,162,0,0,0);
signal scenario_full  : scenario_type := (134,31,129,31,129,30,143,31,79,31,31,31,246,31,59,31,59,30,217,31,183,31,103,31,24,31,217,31,217,30,217,29,158,31,158,30,72,31,72,30,247,31,146,31,146,30,109,31,109,30,8,31,3,31,3,30,181,31,181,31,78,31,208,31,140,31,235,31,140,31,24,31,166,31,166,30,137,31,232,31,63,31,117,31,118,31,87,31,134,31,168,31,147,31,147,30,43,31,16,31,84,31,86,31,127,31,137,31,137,30,95,31,128,31,75,31,40,31,129,31,189,31,111,31,111,30,133,31,65,31,71,31,138,31,237,31,66,31,171,31,202,31,244,31,198,31,182,31,74,31,160,31,10,31,194,31,194,30,100,31,153,31,153,30,81,31,81,30,137,31,189,31,77,31,101,31,196,31,132,31,132,30,91,31,34,31,139,31,213,31,213,30,235,31,235,30,136,31,163,31,228,31,66,31,212,31,201,31,139,31,232,31,14,31,218,31,189,31,189,30,21,31,212,31,212,30,212,29,224,31,21,31,169,31,148,31,148,30,112,31,250,31,250,30,185,31,185,30,10,31,72,31,234,31,112,31,45,31,124,31,141,31,112,31,248,31,88,31,88,30,180,31,180,30,156,31,143,31,10,31,29,31,129,31,129,30,23,31,64,31,64,30,225,31,170,31,170,30,70,31,59,31,203,31,236,31,236,30,236,29,236,28,217,31,101,31,10,31,109,31,109,30,109,29,196,31,240,31,223,31,80,31,1,31,1,30,5,31,5,30,100,31,127,31,224,31,69,31,40,31,40,30,181,31,181,30,79,31,173,31,242,31,111,31,115,31,144,31,114,31,28,31,28,30,31,31,11,31,2,31,27,31,88,31,88,30,162,31,124,31,58,31,50,31,179,31,20,31,93,31,209,31,117,31,142,31,188,31,11,31,71,31,190,31,190,30,172,31,134,31,103,31,247,31,58,31,45,31,22,31,219,31,167,31,208,31,208,30,159,31,252,31,134,31,124,31,194,31,14,31,241,31,247,31,253,31,134,31,87,31,251,31,251,30,251,29,251,28,36,31,36,31,36,30,212,31,77,31,196,31,210,31,29,31,8,31,8,30,131,31,131,31,210,31,187,31,172,31,109,31,124,31,124,30,134,31,154,31,16,31,127,31,51,31,85,31,217,31,217,30,203,31,16,31,111,31,238,31,19,31,44,31,75,31,75,30,75,29,128,31,181,31,226,31,21,31,21,30,186,31,153,31,144,31,144,30,46,31,46,30,69,31,202,31,202,30,136,31,234,31,40,31,106,31,54,31,116,31,116,30,35,31,202,31,39,31,222,31,132,31,77,31,119,31,4,31,25,31,154,31,112,31,89,31,4,31,198,31,84,31,78,31,249,31,51,31,167,31,116,31,101,31,161,31,146,31,152,31,152,30,80,31,80,30,52,31,76,31,32,31,147,31,228,31,5,31,190,31,228,31,34,31,8,31,114,31,114,30,147,31,209,31,209,30,151,31,30,31,30,30,32,31,126,31,148,31,148,30,232,31,33,31,71,31,17,31,197,31,131,31,36,31,149,31,95,31,210,31,78,31,78,30,206,31,245,31,103,31,40,31,104,31,104,30,107,31,251,31,251,30,255,31,223,31,126,31,28,31,232,31,232,30,232,29,78,31,245,31,255,31,128,31,128,30,193,31,111,31,177,31,177,30,31,31,56,31,231,31,189,31,210,31,158,31,23,31,16,31,16,30,106,31,42,31,46,31,193,31,81,31,153,31,200,31,200,30,19,31,247,31,114,31,137,31,190,31,190,30,160,31,31,31,2,31,114,31,47,31,200,31,155,31,155,30,101,31,206,31,206,30,107,31,107,30,216,31,187,31,73,31,31,31,31,30,227,31,153,31,117,31,239,31,247,31,106,31,180,31,88,31,88,30,24,31,107,31,75,31,220,31,220,30,90,31,242,31,80,31,163,31,152,31,147,31,36,31,36,30,85,31,85,30,151,31,151,30,27,31,108,31,186,31,108,31,108,30,63,31,248,31,85,31,164,31,242,31,23,31,23,30,23,29,75,31,172,31,172,30,172,29,184,31,211,31,116,31,109,31,202,31,154,31,21,31,21,30,254,31,67,31,169,31,172,31,125,31,152,31,61,31,124,31,124,30,199,31,224,31,224,30,237,31,189,31,189,30,189,29,129,31,66,31,199,31,129,31,129,30,68,31,68,30,171,31,153,31,192,31,192,30,176,31,126,31,73,31,57,31,57,30,215,31,192,31,164,31,169,31,231,31,146,31,175,31,155,31,249,31,41,31,41,30,9,31,54,31,105,31,56,31,152,31,252,31,252,30,208,31,134,31,120,31,47,31,230,31,230,30,26,31,248,31,72,31,211,31,211,30,105,31,171,31,224,31,20,31,112,31,200,31,200,30,162,31,55,31,55,30,35,31,16,31,66,31,68,31,5,31,54,31,120,31,96,31,67,31,125,31,237,31,88,31,27,31,229,31,172,31,147,31,200,31,251,31,251,30,6,31,240,31,230,31,141,31,132,31,194,31,30,31,159,31,159,30,159,29,67,31,6,31,131,31,28,31,38,31,51,31,109,31,229,31,197,31,66,31,27,31,5,31,5,30,179,31,3,31,3,30,209,31,209,30,209,29,197,31,86,31,114,31,144,31,196,31,171,31,248,31,50,31,50,30,134,31,36,31,171,31,5,31,228,31,161,31,98,31,98,30,99,31,99,30,99,29,99,28,99,27,52,31,174,31,141,31,100,31,1,31,83,31,83,30,83,29,5,31,77,31,50,31,16,31,50,31,40,31,100,31,90,31,165,31,250,31,35,31,35,30,35,29,38,31,41,31,41,30,34,31,239,31,130,31,79,31,136,31,136,30,25,31,183,31,244,31,236,31,83,31,83,30,162,31,162,30,172,31,177,31,177,30,43,31,20,31,44,31,44,30,245,31,181,31,121,31,191,31,219,31,222,31,85,31,156,31,248,31,248,30,248,29,28,31,136,31,167,31,41,31,211,31,141,31,65,31,81,31,9,31,233,31,233,30,26,31,109,31,36,31,112,31,112,30,2,31,98,31,94,31,89,31,115,31,127,31,191,31,204,31,220,31,14,31,236,31,236,30,159,31,204,31,177,31,116,31,226,31,226,30,134,31,74,31,178,31,211,31,175,31,100,31,191,31,191,30,191,29,191,28,191,27,200,31,239,31,1,31,1,30,223,31,74,31,226,31,77,31,225,31,225,30,82,31,82,30,86,31,154,31,242,31,40,31,138,31,138,30,119,31,223,31,3,31,90,31,97,31,14,31,125,31,12,31,5,31,5,30,222,31,1,31,16,31,180,31,207,31,95,31,118,31,118,30,60,31,164,31,164,30,164,29,40,31,196,31,77,31,29,31,1,31,230,31,141,31,141,30,141,29,108,31,57,31,118,31,199,31,237,31,127,31,127,30,79,31,79,30,79,29,249,31,170,31,2,31,87,31,87,30,59,31,59,30,209,31,209,30,202,31,162,31,162,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
