-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 206;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,189,0,105,0,191,0,157,0,82,0,78,0,68,0,0,0,41,0,187,0,183,0,0,0,55,0,0,0,98,0,202,0,16,0,242,0,88,0,68,0,0,0,100,0,127,0,0,0,140,0,0,0,189,0,184,0,178,0,117,0,201,0,0,0,170,0,246,0,54,0,0,0,25,0,83,0,156,0,75,0,135,0,85,0,26,0,212,0,34,0,204,0,50,0,0,0,114,0,104,0,140,0,137,0,174,0,154,0,47,0,255,0,237,0,4,0,254,0,56,0,89,0,42,0,17,0,174,0,242,0,7,0,126,0,97,0,81,0,0,0,248,0,76,0,144,0,252,0,203,0,42,0,36,0,103,0,40,0,216,0,222,0,0,0,0,0,0,0,0,0,144,0,0,0,77,0,196,0,58,0,67,0,121,0,159,0,117,0,100,0,78,0,153,0,242,0,167,0,0,0,212,0,134,0,99,0,51,0,0,0,94,0,214,0,95,0,0,0,0,0,0,0,8,0,44,0,160,0,86,0,7,0,198,0,90,0,105,0,31,0,235,0,246,0,218,0,152,0,200,0,56,0,92,0,209,0,0,0,0,0,0,0,83,0,240,0,133,0,125,0,180,0,58,0,0,0,70,0,249,0,42,0,0,0,118,0,0,0,0,0,119,0,194,0,249,0,237,0,154,0,124,0,158,0,38,0,246,0,0,0,1,0,192,0,183,0,166,0,173,0,31,0,0,0,21,0,255,0,210,0,131,0,224,0,240,0,174,0,0,0,54,0,225,0,199,0,158,0,206,0,159,0,182,0,37,0,37,0,114,0,3,0,118,0,0,0,190,0,191,0,155,0,109,0,145,0,215,0,105,0,0,0,172,0,163,0,0,0,158,0,0,0,68,0,22,0,63,0,0,0,121,0,0,0,0,0,0,0,156,0);
signal scenario_full  : scenario_type := (0,0,189,31,105,31,191,31,157,31,82,31,78,31,68,31,68,30,41,31,187,31,183,31,183,30,55,31,55,30,98,31,202,31,16,31,242,31,88,31,68,31,68,30,100,31,127,31,127,30,140,31,140,30,189,31,184,31,178,31,117,31,201,31,201,30,170,31,246,31,54,31,54,30,25,31,83,31,156,31,75,31,135,31,85,31,26,31,212,31,34,31,204,31,50,31,50,30,114,31,104,31,140,31,137,31,174,31,154,31,47,31,255,31,237,31,4,31,254,31,56,31,89,31,42,31,17,31,174,31,242,31,7,31,126,31,97,31,81,31,81,30,248,31,76,31,144,31,252,31,203,31,42,31,36,31,103,31,40,31,216,31,222,31,222,30,222,29,222,28,222,27,144,31,144,30,77,31,196,31,58,31,67,31,121,31,159,31,117,31,100,31,78,31,153,31,242,31,167,31,167,30,212,31,134,31,99,31,51,31,51,30,94,31,214,31,95,31,95,30,95,29,95,28,8,31,44,31,160,31,86,31,7,31,198,31,90,31,105,31,31,31,235,31,246,31,218,31,152,31,200,31,56,31,92,31,209,31,209,30,209,29,209,28,83,31,240,31,133,31,125,31,180,31,58,31,58,30,70,31,249,31,42,31,42,30,118,31,118,30,118,29,119,31,194,31,249,31,237,31,154,31,124,31,158,31,38,31,246,31,246,30,1,31,192,31,183,31,166,31,173,31,31,31,31,30,21,31,255,31,210,31,131,31,224,31,240,31,174,31,174,30,54,31,225,31,199,31,158,31,206,31,159,31,182,31,37,31,37,31,114,31,3,31,118,31,118,30,190,31,191,31,155,31,109,31,145,31,215,31,105,31,105,30,172,31,163,31,163,30,158,31,158,30,68,31,22,31,63,31,63,30,121,31,121,30,121,29,121,28,156,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
