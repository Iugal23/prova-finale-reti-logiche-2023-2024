-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 785;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (162,0,232,0,141,0,78,0,172,0,161,0,69,0,118,0,1,0,0,0,0,0,156,0,66,0,118,0,0,0,0,0,167,0,113,0,124,0,0,0,13,0,68,0,65,0,0,0,69,0,139,0,201,0,56,0,127,0,227,0,133,0,114,0,186,0,0,0,92,0,150,0,166,0,0,0,143,0,158,0,233,0,3,0,9,0,131,0,130,0,0,0,0,0,0,0,58,0,204,0,108,0,251,0,24,0,0,0,222,0,0,0,36,0,233,0,39,0,179,0,194,0,74,0,7,0,26,0,90,0,198,0,70,0,133,0,147,0,124,0,216,0,180,0,83,0,210,0,248,0,48,0,0,0,55,0,0,0,252,0,122,0,194,0,0,0,46,0,87,0,0,0,21,0,47,0,0,0,55,0,46,0,151,0,138,0,75,0,101,0,0,0,195,0,180,0,239,0,137,0,171,0,174,0,192,0,62,0,213,0,0,0,0,0,48,0,0,0,27,0,0,0,0,0,255,0,120,0,167,0,66,0,104,0,23,0,0,0,0,0,221,0,23,0,16,0,25,0,62,0,77,0,202,0,84,0,67,0,145,0,79,0,0,0,170,0,213,0,118,0,0,0,56,0,139,0,194,0,177,0,170,0,227,0,131,0,176,0,0,0,160,0,0,0,0,0,0,0,103,0,60,0,1,0,18,0,229,0,214,0,158,0,103,0,0,0,96,0,80,0,64,0,36,0,75,0,0,0,45,0,139,0,0,0,35,0,50,0,0,0,0,0,10,0,15,0,58,0,140,0,70,0,123,0,208,0,91,0,0,0,39,0,21,0,48,0,223,0,97,0,172,0,0,0,38,0,96,0,15,0,0,0,226,0,173,0,61,0,180,0,0,0,204,0,29,0,40,0,93,0,0,0,132,0,155,0,55,0,0,0,190,0,250,0,200,0,16,0,230,0,168,0,26,0,134,0,3,0,0,0,173,0,0,0,0,0,19,0,153,0,219,0,28,0,1,0,54,0,195,0,0,0,67,0,117,0,70,0,161,0,87,0,19,0,65,0,0,0,165,0,58,0,22,0,152,0,99,0,240,0,122,0,171,0,0,0,0,0,30,0,0,0,0,0,54,0,200,0,5,0,0,0,32,0,0,0,181,0,46,0,221,0,0,0,149,0,0,0,129,0,199,0,120,0,234,0,104,0,187,0,206,0,83,0,221,0,0,0,0,0,0,0,136,0,238,0,0,0,52,0,143,0,160,0,239,0,26,0,0,0,19,0,239,0,132,0,0,0,128,0,54,0,253,0,0,0,217,0,203,0,0,0,135,0,197,0,120,0,119,0,142,0,86,0,176,0,227,0,0,0,0,0,7,0,88,0,48,0,5,0,0,0,179,0,108,0,99,0,123,0,177,0,124,0,195,0,70,0,0,0,110,0,46,0,199,0,219,0,148,0,138,0,0,0,87,0,231,0,17,0,45,0,98,0,231,0,70,0,86,0,125,0,0,0,52,0,97,0,31,0,38,0,0,0,28,0,209,0,145,0,87,0,89,0,129,0,6,0,173,0,157,0,213,0,50,0,122,0,129,0,225,0,0,0,168,0,246,0,69,0,102,0,0,0,0,0,173,0,0,0,249,0,126,0,234,0,9,0,208,0,0,0,238,0,243,0,87,0,96,0,200,0,63,0,67,0,171,0,251,0,125,0,70,0,108,0,134,0,226,0,91,0,104,0,160,0,0,0,31,0,70,0,26,0,0,0,175,0,156,0,0,0,0,0,148,0,70,0,216,0,0,0,0,0,0,0,180,0,0,0,232,0,52,0,0,0,39,0,122,0,144,0,100,0,127,0,142,0,231,0,47,0,5,0,203,0,144,0,31,0,185,0,0,0,0,0,0,0,175,0,89,0,133,0,94,0,16,0,0,0,60,0,0,0,25,0,201,0,0,0,70,0,70,0,242,0,0,0,57,0,209,0,94,0,68,0,0,0,187,0,247,0,108,0,132,0,74,0,70,0,183,0,0,0,192,0,42,0,73,0,85,0,213,0,66,0,0,0,0,0,198,0,0,0,98,0,219,0,101,0,0,0,55,0,153,0,146,0,209,0,219,0,0,0,0,0,22,0,0,0,199,0,66,0,248,0,5,0,0,0,0,0,171,0,69,0,156,0,42,0,34,0,44,0,110,0,177,0,40,0,43,0,77,0,254,0,193,0,79,0,187,0,227,0,78,0,0,0,239,0,104,0,159,0,35,0,250,0,0,0,68,0,154,0,211,0,195,0,0,0,0,0,222,0,86,0,0,0,113,0,167,0,37,0,104,0,118,0,109,0,115,0,39,0,169,0,34,0,254,0,198,0,14,0,0,0,246,0,67,0,199,0,51,0,106,0,12,0,159,0,0,0,68,0,86,0,212,0,149,0,48,0,25,0,0,0,142,0,251,0,167,0,0,0,0,0,221,0,154,0,135,0,145,0,14,0,94,0,50,0,40,0,43,0,184,0,140,0,15,0,183,0,103,0,76,0,0,0,212,0,0,0,14,0,0,0,4,0,115,0,0,0,146,0,81,0,46,0,133,0,83,0,52,0,62,0,141,0,0,0,31,0,0,0,224,0,8,0,162,0,50,0,0,0,125,0,140,0,93,0,200,0,204,0,35,0,74,0,142,0,83,0,0,0,149,0,20,0,73,0,28,0,0,0,0,0,74,0,125,0,222,0,241,0,185,0,148,0,0,0,185,0,43,0,225,0,21,0,220,0,187,0,163,0,211,0,0,0,238,0,1,0,126,0,0,0,218,0,132,0,0,0,0,0,176,0,88,0,131,0,176,0,249,0,0,0,187,0,162,0,97,0,138,0,18,0,234,0,205,0,146,0,93,0,221,0,64,0,54,0,47,0,30,0,172,0,202,0,173,0,0,0,0,0,13,0,240,0,182,0,129,0,7,0,138,0,27,0,240,0,130,0,19,0,219,0,135,0,129,0,243,0,80,0,67,0,143,0,246,0,171,0,40,0,0,0,213,0,0,0,153,0,0,0,174,0,119,0,176,0,125,0,102,0,0,0,243,0,79,0,52,0,237,0,121,0,0,0,176,0,0,0,102,0,0,0,129,0,247,0,62,0,99,0,219,0,15,0,210,0,67,0,65,0,55,0,231,0,247,0,87,0,120,0,159,0,206,0,56,0,130,0,29,0,15,0,60,0,0,0,40,0,0,0,230,0,6,0,140,0,27,0,140,0,95,0,0,0,0,0,44,0,86,0,178,0,222,0,151,0,19,0,161,0,191,0,2,0,76,0,0,0,33,0,0,0,25,0,163,0,134,0,0,0,233,0,82,0,89,0,183,0,0,0,209,0,0,0,178,0,124,0,163,0,32,0,55,0,0,0,0,0,164,0,4,0,0,0,54,0,20,0,238,0,222,0,136,0,82,0,0,0,48,0,202,0,106,0,201,0,85,0,113,0,101,0,0,0,93,0,34,0,9,0,32,0,49,0,32,0,0,0,0,0,175,0,0,0,186,0,227,0,78,0,160,0,161,0,74,0);
signal scenario_full  : scenario_type := (162,31,232,31,141,31,78,31,172,31,161,31,69,31,118,31,1,31,1,30,1,29,156,31,66,31,118,31,118,30,118,29,167,31,113,31,124,31,124,30,13,31,68,31,65,31,65,30,69,31,139,31,201,31,56,31,127,31,227,31,133,31,114,31,186,31,186,30,92,31,150,31,166,31,166,30,143,31,158,31,233,31,3,31,9,31,131,31,130,31,130,30,130,29,130,28,58,31,204,31,108,31,251,31,24,31,24,30,222,31,222,30,36,31,233,31,39,31,179,31,194,31,74,31,7,31,26,31,90,31,198,31,70,31,133,31,147,31,124,31,216,31,180,31,83,31,210,31,248,31,48,31,48,30,55,31,55,30,252,31,122,31,194,31,194,30,46,31,87,31,87,30,21,31,47,31,47,30,55,31,46,31,151,31,138,31,75,31,101,31,101,30,195,31,180,31,239,31,137,31,171,31,174,31,192,31,62,31,213,31,213,30,213,29,48,31,48,30,27,31,27,30,27,29,255,31,120,31,167,31,66,31,104,31,23,31,23,30,23,29,221,31,23,31,16,31,25,31,62,31,77,31,202,31,84,31,67,31,145,31,79,31,79,30,170,31,213,31,118,31,118,30,56,31,139,31,194,31,177,31,170,31,227,31,131,31,176,31,176,30,160,31,160,30,160,29,160,28,103,31,60,31,1,31,18,31,229,31,214,31,158,31,103,31,103,30,96,31,80,31,64,31,36,31,75,31,75,30,45,31,139,31,139,30,35,31,50,31,50,30,50,29,10,31,15,31,58,31,140,31,70,31,123,31,208,31,91,31,91,30,39,31,21,31,48,31,223,31,97,31,172,31,172,30,38,31,96,31,15,31,15,30,226,31,173,31,61,31,180,31,180,30,204,31,29,31,40,31,93,31,93,30,132,31,155,31,55,31,55,30,190,31,250,31,200,31,16,31,230,31,168,31,26,31,134,31,3,31,3,30,173,31,173,30,173,29,19,31,153,31,219,31,28,31,1,31,54,31,195,31,195,30,67,31,117,31,70,31,161,31,87,31,19,31,65,31,65,30,165,31,58,31,22,31,152,31,99,31,240,31,122,31,171,31,171,30,171,29,30,31,30,30,30,29,54,31,200,31,5,31,5,30,32,31,32,30,181,31,46,31,221,31,221,30,149,31,149,30,129,31,199,31,120,31,234,31,104,31,187,31,206,31,83,31,221,31,221,30,221,29,221,28,136,31,238,31,238,30,52,31,143,31,160,31,239,31,26,31,26,30,19,31,239,31,132,31,132,30,128,31,54,31,253,31,253,30,217,31,203,31,203,30,135,31,197,31,120,31,119,31,142,31,86,31,176,31,227,31,227,30,227,29,7,31,88,31,48,31,5,31,5,30,179,31,108,31,99,31,123,31,177,31,124,31,195,31,70,31,70,30,110,31,46,31,199,31,219,31,148,31,138,31,138,30,87,31,231,31,17,31,45,31,98,31,231,31,70,31,86,31,125,31,125,30,52,31,97,31,31,31,38,31,38,30,28,31,209,31,145,31,87,31,89,31,129,31,6,31,173,31,157,31,213,31,50,31,122,31,129,31,225,31,225,30,168,31,246,31,69,31,102,31,102,30,102,29,173,31,173,30,249,31,126,31,234,31,9,31,208,31,208,30,238,31,243,31,87,31,96,31,200,31,63,31,67,31,171,31,251,31,125,31,70,31,108,31,134,31,226,31,91,31,104,31,160,31,160,30,31,31,70,31,26,31,26,30,175,31,156,31,156,30,156,29,148,31,70,31,216,31,216,30,216,29,216,28,180,31,180,30,232,31,52,31,52,30,39,31,122,31,144,31,100,31,127,31,142,31,231,31,47,31,5,31,203,31,144,31,31,31,185,31,185,30,185,29,185,28,175,31,89,31,133,31,94,31,16,31,16,30,60,31,60,30,25,31,201,31,201,30,70,31,70,31,242,31,242,30,57,31,209,31,94,31,68,31,68,30,187,31,247,31,108,31,132,31,74,31,70,31,183,31,183,30,192,31,42,31,73,31,85,31,213,31,66,31,66,30,66,29,198,31,198,30,98,31,219,31,101,31,101,30,55,31,153,31,146,31,209,31,219,31,219,30,219,29,22,31,22,30,199,31,66,31,248,31,5,31,5,30,5,29,171,31,69,31,156,31,42,31,34,31,44,31,110,31,177,31,40,31,43,31,77,31,254,31,193,31,79,31,187,31,227,31,78,31,78,30,239,31,104,31,159,31,35,31,250,31,250,30,68,31,154,31,211,31,195,31,195,30,195,29,222,31,86,31,86,30,113,31,167,31,37,31,104,31,118,31,109,31,115,31,39,31,169,31,34,31,254,31,198,31,14,31,14,30,246,31,67,31,199,31,51,31,106,31,12,31,159,31,159,30,68,31,86,31,212,31,149,31,48,31,25,31,25,30,142,31,251,31,167,31,167,30,167,29,221,31,154,31,135,31,145,31,14,31,94,31,50,31,40,31,43,31,184,31,140,31,15,31,183,31,103,31,76,31,76,30,212,31,212,30,14,31,14,30,4,31,115,31,115,30,146,31,81,31,46,31,133,31,83,31,52,31,62,31,141,31,141,30,31,31,31,30,224,31,8,31,162,31,50,31,50,30,125,31,140,31,93,31,200,31,204,31,35,31,74,31,142,31,83,31,83,30,149,31,20,31,73,31,28,31,28,30,28,29,74,31,125,31,222,31,241,31,185,31,148,31,148,30,185,31,43,31,225,31,21,31,220,31,187,31,163,31,211,31,211,30,238,31,1,31,126,31,126,30,218,31,132,31,132,30,132,29,176,31,88,31,131,31,176,31,249,31,249,30,187,31,162,31,97,31,138,31,18,31,234,31,205,31,146,31,93,31,221,31,64,31,54,31,47,31,30,31,172,31,202,31,173,31,173,30,173,29,13,31,240,31,182,31,129,31,7,31,138,31,27,31,240,31,130,31,19,31,219,31,135,31,129,31,243,31,80,31,67,31,143,31,246,31,171,31,40,31,40,30,213,31,213,30,153,31,153,30,174,31,119,31,176,31,125,31,102,31,102,30,243,31,79,31,52,31,237,31,121,31,121,30,176,31,176,30,102,31,102,30,129,31,247,31,62,31,99,31,219,31,15,31,210,31,67,31,65,31,55,31,231,31,247,31,87,31,120,31,159,31,206,31,56,31,130,31,29,31,15,31,60,31,60,30,40,31,40,30,230,31,6,31,140,31,27,31,140,31,95,31,95,30,95,29,44,31,86,31,178,31,222,31,151,31,19,31,161,31,191,31,2,31,76,31,76,30,33,31,33,30,25,31,163,31,134,31,134,30,233,31,82,31,89,31,183,31,183,30,209,31,209,30,178,31,124,31,163,31,32,31,55,31,55,30,55,29,164,31,4,31,4,30,54,31,20,31,238,31,222,31,136,31,82,31,82,30,48,31,202,31,106,31,201,31,85,31,113,31,101,31,101,30,93,31,34,31,9,31,32,31,49,31,32,31,32,30,32,29,175,31,175,30,186,31,227,31,78,31,160,31,161,31,74,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
