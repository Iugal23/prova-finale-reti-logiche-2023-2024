-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 719;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (245,0,88,0,60,0,44,0,23,0,254,0,117,0,4,0,16,0,0,0,26,0,192,0,241,0,157,0,0,0,81,0,208,0,101,0,254,0,106,0,0,0,25,0,216,0,76,0,67,0,250,0,251,0,32,0,41,0,0,0,55,0,28,0,49,0,118,0,98,0,232,0,156,0,83,0,174,0,98,0,132,0,0,0,254,0,208,0,74,0,33,0,131,0,202,0,246,0,112,0,227,0,87,0,0,0,167,0,60,0,0,0,160,0,192,0,250,0,147,0,92,0,181,0,0,0,240,0,100,0,250,0,65,0,108,0,27,0,120,0,174,0,0,0,219,0,205,0,0,0,215,0,146,0,9,0,103,0,158,0,12,0,29,0,25,0,5,0,235,0,83,0,98,0,182,0,242,0,39,0,186,0,58,0,22,0,0,0,127,0,47,0,0,0,0,0,13,0,118,0,4,0,238,0,125,0,111,0,152,0,35,0,21,0,115,0,212,0,131,0,113,0,27,0,213,0,83,0,217,0,134,0,105,0,153,0,12,0,28,0,118,0,236,0,61,0,0,0,230,0,237,0,112,0,136,0,77,0,150,0,170,0,0,0,0,0,146,0,15,0,75,0,108,0,214,0,126,0,165,0,171,0,3,0,139,0,58,0,233,0,133,0,37,0,65,0,0,0,248,0,109,0,0,0,0,0,96,0,149,0,0,0,0,0,55,0,0,0,0,0,6,0,116,0,219,0,94,0,140,0,16,0,197,0,9,0,186,0,76,0,105,0,11,0,0,0,133,0,0,0,90,0,176,0,22,0,176,0,0,0,247,0,0,0,14,0,171,0,95,0,0,0,51,0,159,0,78,0,0,0,5,0,105,0,221,0,0,0,155,0,177,0,66,0,0,0,179,0,215,0,61,0,52,0,105,0,0,0,237,0,22,0,52,0,0,0,0,0,0,0,80,0,0,0,5,0,188,0,167,0,4,0,0,0,127,0,181,0,86,0,223,0,154,0,0,0,109,0,159,0,95,0,229,0,73,0,18,0,161,0,66,0,76,0,214,0,49,0,129,0,211,0,64,0,141,0,37,0,0,0,69,0,209,0,128,0,68,0,215,0,193,0,221,0,92,0,0,0,90,0,191,0,249,0,132,0,126,0,0,0,184,0,39,0,39,0,54,0,220,0,240,0,48,0,0,0,187,0,0,0,163,0,230,0,0,0,202,0,207,0,200,0,25,0,219,0,0,0,246,0,0,0,222,0,13,0,0,0,191,0,0,0,140,0,66,0,39,0,5,0,185,0,69,0,0,0,104,0,148,0,91,0,208,0,154,0,93,0,30,0,239,0,168,0,156,0,112,0,192,0,0,0,144,0,194,0,185,0,154,0,187,0,211,0,129,0,95,0,99,0,168,0,245,0,177,0,154,0,152,0,61,0,183,0,205,0,0,0,76,0,229,0,178,0,0,0,67,0,61,0,187,0,87,0,19,0,0,0,60,0,147,0,58,0,0,0,0,0,123,0,180,0,179,0,37,0,4,0,20,0,0,0,0,0,0,0,101,0,188,0,16,0,0,0,20,0,232,0,88,0,197,0,74,0,173,0,241,0,107,0,0,0,0,0,28,0,86,0,86,0,179,0,228,0,239,0,36,0,214,0,151,0,251,0,191,0,249,0,160,0,177,0,249,0,0,0,56,0,23,0,4,0,14,0,212,0,30,0,103,0,219,0,69,0,0,0,53,0,37,0,215,0,167,0,163,0,74,0,3,0,100,0,20,0,58,0,208,0,208,0,0,0,135,0,42,0,31,0,55,0,61,0,28,0,241,0,43,0,0,0,0,0,205,0,50,0,80,0,136,0,210,0,140,0,0,0,187,0,158,0,141,0,0,0,59,0,203,0,0,0,0,0,253,0,169,0,59,0,103,0,88,0,212,0,0,0,0,0,70,0,0,0,188,0,205,0,213,0,2,0,227,0,206,0,27,0,51,0,11,0,0,0,0,0,0,0,0,0,0,0,255,0,122,0,212,0,18,0,79,0,211,0,18,0,204,0,33,0,193,0,0,0,11,0,0,0,48,0,166,0,232,0,0,0,12,0,0,0,217,0,162,0,109,0,1,0,70,0,236,0,0,0,0,0,174,0,2,0,133,0,53,0,53,0,255,0,60,0,0,0,205,0,54,0,207,0,219,0,127,0,185,0,187,0,0,0,83,0,5,0,63,0,117,0,9,0,38,0,108,0,0,0,24,0,0,0,155,0,222,0,248,0,70,0,0,0,253,0,139,0,123,0,227,0,0,0,0,0,240,0,21,0,6,0,49,0,0,0,181,0,120,0,228,0,140,0,135,0,11,0,131,0,152,0,17,0,84,0,238,0,229,0,155,0,72,0,114,0,87,0,122,0,38,0,220,0,73,0,117,0,6,0,212,0,123,0,133,0,230,0,246,0,136,0,167,0,0,0,0,0,213,0,95,0,39,0,109,0,112,0,169,0,182,0,187,0,0,0,47,0,88,0,150,0,131,0,153,0,90,0,0,0,42,0,228,0,159,0,19,0,132,0,40,0,100,0,73,0,0,0,60,0,0,0,95,0,197,0,240,0,0,0,0,0,121,0,197,0,0,0,254,0,56,0,207,0,171,0,74,0,0,0,0,0,253,0,44,0,210,0,158,0,113,0,88,0,92,0,0,0,210,0,71,0,233,0,247,0,104,0,122,0,77,0,85,0,233,0,106,0,218,0,89,0,121,0,2,0,232,0,128,0,0,0,0,0,0,0,92,0,0,0,0,0,0,0,34,0,156,0,251,0,38,0,167,0,82,0,0,0,153,0,78,0,223,0,99,0,0,0,247,0,219,0,105,0,181,0,0,0,0,0,121,0,0,0,92,0,244,0,109,0,5,0,167,0,31,0,31,0,214,0,12,0,44,0,0,0,93,0,41,0,144,0,45,0,0,0,131,0,0,0,2,0,39,0,131,0,181,0,132,0,119,0,242,0,128,0,0,0,181,0,14,0,215,0,115,0,143,0,82,0,0,0,63,0,0,0,171,0,43,0,0,0,127,0,5,0,141,0,0,0,136,0,61,0,25,0,133,0,25,0,144,0,156,0,55,0,248,0,34,0,136,0,113,0,52,0,0,0,88,0,0,0,0,0,46,0,199,0,124,0,0,0,151,0,183,0,168,0,8,0,139,0,154,0,0,0,0,0,191,0,0,0,70,0,0,0,199,0,120,0,159,0,39,0,118,0);
signal scenario_full  : scenario_type := (245,31,88,31,60,31,44,31,23,31,254,31,117,31,4,31,16,31,16,30,26,31,192,31,241,31,157,31,157,30,81,31,208,31,101,31,254,31,106,31,106,30,25,31,216,31,76,31,67,31,250,31,251,31,32,31,41,31,41,30,55,31,28,31,49,31,118,31,98,31,232,31,156,31,83,31,174,31,98,31,132,31,132,30,254,31,208,31,74,31,33,31,131,31,202,31,246,31,112,31,227,31,87,31,87,30,167,31,60,31,60,30,160,31,192,31,250,31,147,31,92,31,181,31,181,30,240,31,100,31,250,31,65,31,108,31,27,31,120,31,174,31,174,30,219,31,205,31,205,30,215,31,146,31,9,31,103,31,158,31,12,31,29,31,25,31,5,31,235,31,83,31,98,31,182,31,242,31,39,31,186,31,58,31,22,31,22,30,127,31,47,31,47,30,47,29,13,31,118,31,4,31,238,31,125,31,111,31,152,31,35,31,21,31,115,31,212,31,131,31,113,31,27,31,213,31,83,31,217,31,134,31,105,31,153,31,12,31,28,31,118,31,236,31,61,31,61,30,230,31,237,31,112,31,136,31,77,31,150,31,170,31,170,30,170,29,146,31,15,31,75,31,108,31,214,31,126,31,165,31,171,31,3,31,139,31,58,31,233,31,133,31,37,31,65,31,65,30,248,31,109,31,109,30,109,29,96,31,149,31,149,30,149,29,55,31,55,30,55,29,6,31,116,31,219,31,94,31,140,31,16,31,197,31,9,31,186,31,76,31,105,31,11,31,11,30,133,31,133,30,90,31,176,31,22,31,176,31,176,30,247,31,247,30,14,31,171,31,95,31,95,30,51,31,159,31,78,31,78,30,5,31,105,31,221,31,221,30,155,31,177,31,66,31,66,30,179,31,215,31,61,31,52,31,105,31,105,30,237,31,22,31,52,31,52,30,52,29,52,28,80,31,80,30,5,31,188,31,167,31,4,31,4,30,127,31,181,31,86,31,223,31,154,31,154,30,109,31,159,31,95,31,229,31,73,31,18,31,161,31,66,31,76,31,214,31,49,31,129,31,211,31,64,31,141,31,37,31,37,30,69,31,209,31,128,31,68,31,215,31,193,31,221,31,92,31,92,30,90,31,191,31,249,31,132,31,126,31,126,30,184,31,39,31,39,31,54,31,220,31,240,31,48,31,48,30,187,31,187,30,163,31,230,31,230,30,202,31,207,31,200,31,25,31,219,31,219,30,246,31,246,30,222,31,13,31,13,30,191,31,191,30,140,31,66,31,39,31,5,31,185,31,69,31,69,30,104,31,148,31,91,31,208,31,154,31,93,31,30,31,239,31,168,31,156,31,112,31,192,31,192,30,144,31,194,31,185,31,154,31,187,31,211,31,129,31,95,31,99,31,168,31,245,31,177,31,154,31,152,31,61,31,183,31,205,31,205,30,76,31,229,31,178,31,178,30,67,31,61,31,187,31,87,31,19,31,19,30,60,31,147,31,58,31,58,30,58,29,123,31,180,31,179,31,37,31,4,31,20,31,20,30,20,29,20,28,101,31,188,31,16,31,16,30,20,31,232,31,88,31,197,31,74,31,173,31,241,31,107,31,107,30,107,29,28,31,86,31,86,31,179,31,228,31,239,31,36,31,214,31,151,31,251,31,191,31,249,31,160,31,177,31,249,31,249,30,56,31,23,31,4,31,14,31,212,31,30,31,103,31,219,31,69,31,69,30,53,31,37,31,215,31,167,31,163,31,74,31,3,31,100,31,20,31,58,31,208,31,208,31,208,30,135,31,42,31,31,31,55,31,61,31,28,31,241,31,43,31,43,30,43,29,205,31,50,31,80,31,136,31,210,31,140,31,140,30,187,31,158,31,141,31,141,30,59,31,203,31,203,30,203,29,253,31,169,31,59,31,103,31,88,31,212,31,212,30,212,29,70,31,70,30,188,31,205,31,213,31,2,31,227,31,206,31,27,31,51,31,11,31,11,30,11,29,11,28,11,27,11,26,255,31,122,31,212,31,18,31,79,31,211,31,18,31,204,31,33,31,193,31,193,30,11,31,11,30,48,31,166,31,232,31,232,30,12,31,12,30,217,31,162,31,109,31,1,31,70,31,236,31,236,30,236,29,174,31,2,31,133,31,53,31,53,31,255,31,60,31,60,30,205,31,54,31,207,31,219,31,127,31,185,31,187,31,187,30,83,31,5,31,63,31,117,31,9,31,38,31,108,31,108,30,24,31,24,30,155,31,222,31,248,31,70,31,70,30,253,31,139,31,123,31,227,31,227,30,227,29,240,31,21,31,6,31,49,31,49,30,181,31,120,31,228,31,140,31,135,31,11,31,131,31,152,31,17,31,84,31,238,31,229,31,155,31,72,31,114,31,87,31,122,31,38,31,220,31,73,31,117,31,6,31,212,31,123,31,133,31,230,31,246,31,136,31,167,31,167,30,167,29,213,31,95,31,39,31,109,31,112,31,169,31,182,31,187,31,187,30,47,31,88,31,150,31,131,31,153,31,90,31,90,30,42,31,228,31,159,31,19,31,132,31,40,31,100,31,73,31,73,30,60,31,60,30,95,31,197,31,240,31,240,30,240,29,121,31,197,31,197,30,254,31,56,31,207,31,171,31,74,31,74,30,74,29,253,31,44,31,210,31,158,31,113,31,88,31,92,31,92,30,210,31,71,31,233,31,247,31,104,31,122,31,77,31,85,31,233,31,106,31,218,31,89,31,121,31,2,31,232,31,128,31,128,30,128,29,128,28,92,31,92,30,92,29,92,28,34,31,156,31,251,31,38,31,167,31,82,31,82,30,153,31,78,31,223,31,99,31,99,30,247,31,219,31,105,31,181,31,181,30,181,29,121,31,121,30,92,31,244,31,109,31,5,31,167,31,31,31,31,31,214,31,12,31,44,31,44,30,93,31,41,31,144,31,45,31,45,30,131,31,131,30,2,31,39,31,131,31,181,31,132,31,119,31,242,31,128,31,128,30,181,31,14,31,215,31,115,31,143,31,82,31,82,30,63,31,63,30,171,31,43,31,43,30,127,31,5,31,141,31,141,30,136,31,61,31,25,31,133,31,25,31,144,31,156,31,55,31,248,31,34,31,136,31,113,31,52,31,52,30,88,31,88,30,88,29,46,31,199,31,124,31,124,30,151,31,183,31,168,31,8,31,139,31,154,31,154,30,154,29,191,31,191,30,70,31,70,30,199,31,120,31,159,31,39,31,118,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
