-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 376;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (154,0,183,0,243,0,144,0,104,0,97,0,0,0,252,0,18,0,0,0,131,0,122,0,210,0,46,0,41,0,87,0,0,0,0,0,200,0,123,0,97,0,172,0,246,0,72,0,90,0,103,0,209,0,96,0,0,0,119,0,43,0,12,0,243,0,192,0,0,0,204,0,47,0,180,0,176,0,249,0,187,0,244,0,0,0,192,0,87,0,187,0,7,0,133,0,222,0,240,0,20,0,0,0,50,0,178,0,110,0,0,0,106,0,116,0,47,0,230,0,84,0,0,0,42,0,0,0,186,0,0,0,145,0,14,0,212,0,0,0,44,0,0,0,199,0,213,0,80,0,23,0,0,0,211,0,0,0,10,0,240,0,0,0,131,0,88,0,109,0,0,0,0,0,98,0,225,0,30,0,141,0,83,0,213,0,97,0,212,0,12,0,0,0,100,0,212,0,75,0,56,0,127,0,0,0,0,0,135,0,9,0,155,0,212,0,170,0,0,0,86,0,125,0,0,0,0,0,25,0,0,0,178,0,0,0,82,0,209,0,0,0,0,0,251,0,0,0,158,0,217,0,129,0,10,0,168,0,205,0,13,0,124,0,57,0,0,0,152,0,243,0,0,0,169,0,124,0,229,0,0,0,3,0,0,0,247,0,80,0,254,0,171,0,137,0,199,0,85,0,0,0,82,0,126,0,0,0,0,0,177,0,212,0,82,0,0,0,28,0,85,0,230,0,0,0,127,0,90,0,243,0,0,0,195,0,164,0,0,0,0,0,43,0,255,0,13,0,179,0,80,0,88,0,59,0,0,0,190,0,0,0,80,0,0,0,128,0,193,0,129,0,181,0,206,0,42,0,52,0,67,0,106,0,33,0,0,0,100,0,0,0,83,0,209,0,77,0,223,0,0,0,0,0,116,0,0,0,0,0,247,0,0,0,0,0,232,0,205,0,144,0,167,0,29,0,0,0,0,0,0,0,0,0,80,0,161,0,93,0,42,0,0,0,177,0,4,0,188,0,0,0,123,0,81,0,0,0,252,0,67,0,62,0,0,0,221,0,64,0,198,0,0,0,235,0,124,0,111,0,10,0,116,0,0,0,187,0,134,0,0,0,252,0,254,0,67,0,0,0,74,0,0,0,244,0,104,0,82,0,178,0,55,0,93,0,120,0,55,0,24,0,157,0,110,0,0,0,29,0,134,0,253,0,0,0,221,0,75,0,51,0,208,0,98,0,222,0,236,0,118,0,171,0,17,0,0,0,117,0,103,0,142,0,0,0,122,0,170,0,76,0,56,0,42,0,238,0,176,0,210,0,223,0,5,0,26,0,82,0,184,0,106,0,0,0,199,0,134,0,166,0,28,0,141,0,185,0,71,0,218,0,140,0,147,0,62,0,52,0,237,0,86,0,189,0,255,0,0,0,111,0,42,0,82,0,253,0,202,0,0,0,42,0,215,0,88,0,129,0,203,0,8,0,57,0,0,0,181,0,79,0,0,0,146,0,0,0,0,0,24,0,150,0,230,0,124,0,173,0,42,0,0,0,53,0,41,0,133,0,159,0,179,0,131,0,0,0,10,0,245,0,231,0,0,0,103,0,126,0,196,0,164,0,112,0,45,0,205,0,138,0,251,0,163,0,184,0,70,0,0,0,203,0,79,0,237,0,129,0,1,0,0,0,102,0,0,0,93,0,159,0);
signal scenario_full  : scenario_type := (154,31,183,31,243,31,144,31,104,31,97,31,97,30,252,31,18,31,18,30,131,31,122,31,210,31,46,31,41,31,87,31,87,30,87,29,200,31,123,31,97,31,172,31,246,31,72,31,90,31,103,31,209,31,96,31,96,30,119,31,43,31,12,31,243,31,192,31,192,30,204,31,47,31,180,31,176,31,249,31,187,31,244,31,244,30,192,31,87,31,187,31,7,31,133,31,222,31,240,31,20,31,20,30,50,31,178,31,110,31,110,30,106,31,116,31,47,31,230,31,84,31,84,30,42,31,42,30,186,31,186,30,145,31,14,31,212,31,212,30,44,31,44,30,199,31,213,31,80,31,23,31,23,30,211,31,211,30,10,31,240,31,240,30,131,31,88,31,109,31,109,30,109,29,98,31,225,31,30,31,141,31,83,31,213,31,97,31,212,31,12,31,12,30,100,31,212,31,75,31,56,31,127,31,127,30,127,29,135,31,9,31,155,31,212,31,170,31,170,30,86,31,125,31,125,30,125,29,25,31,25,30,178,31,178,30,82,31,209,31,209,30,209,29,251,31,251,30,158,31,217,31,129,31,10,31,168,31,205,31,13,31,124,31,57,31,57,30,152,31,243,31,243,30,169,31,124,31,229,31,229,30,3,31,3,30,247,31,80,31,254,31,171,31,137,31,199,31,85,31,85,30,82,31,126,31,126,30,126,29,177,31,212,31,82,31,82,30,28,31,85,31,230,31,230,30,127,31,90,31,243,31,243,30,195,31,164,31,164,30,164,29,43,31,255,31,13,31,179,31,80,31,88,31,59,31,59,30,190,31,190,30,80,31,80,30,128,31,193,31,129,31,181,31,206,31,42,31,52,31,67,31,106,31,33,31,33,30,100,31,100,30,83,31,209,31,77,31,223,31,223,30,223,29,116,31,116,30,116,29,247,31,247,30,247,29,232,31,205,31,144,31,167,31,29,31,29,30,29,29,29,28,29,27,80,31,161,31,93,31,42,31,42,30,177,31,4,31,188,31,188,30,123,31,81,31,81,30,252,31,67,31,62,31,62,30,221,31,64,31,198,31,198,30,235,31,124,31,111,31,10,31,116,31,116,30,187,31,134,31,134,30,252,31,254,31,67,31,67,30,74,31,74,30,244,31,104,31,82,31,178,31,55,31,93,31,120,31,55,31,24,31,157,31,110,31,110,30,29,31,134,31,253,31,253,30,221,31,75,31,51,31,208,31,98,31,222,31,236,31,118,31,171,31,17,31,17,30,117,31,103,31,142,31,142,30,122,31,170,31,76,31,56,31,42,31,238,31,176,31,210,31,223,31,5,31,26,31,82,31,184,31,106,31,106,30,199,31,134,31,166,31,28,31,141,31,185,31,71,31,218,31,140,31,147,31,62,31,52,31,237,31,86,31,189,31,255,31,255,30,111,31,42,31,82,31,253,31,202,31,202,30,42,31,215,31,88,31,129,31,203,31,8,31,57,31,57,30,181,31,79,31,79,30,146,31,146,30,146,29,24,31,150,31,230,31,124,31,173,31,42,31,42,30,53,31,41,31,133,31,159,31,179,31,131,31,131,30,10,31,245,31,231,31,231,30,103,31,126,31,196,31,164,31,112,31,45,31,205,31,138,31,251,31,163,31,184,31,70,31,70,30,203,31,79,31,237,31,129,31,1,31,1,30,102,31,102,30,93,31,159,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
