-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_93 is
end project_tb_93;

architecture project_tb_arch_93 of project_tb_93 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 591;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (253,0,32,0,7,0,135,0,165,0,9,0,220,0,0,0,0,0,128,0,241,0,209,0,149,0,69,0,0,0,95,0,38,0,108,0,50,0,70,0,144,0,96,0,246,0,72,0,60,0,0,0,0,0,62,0,21,0,21,0,82,0,75,0,0,0,41,0,13,0,235,0,0,0,170,0,178,0,253,0,0,0,33,0,44,0,97,0,96,0,30,0,0,0,249,0,35,0,87,0,124,0,56,0,60,0,203,0,0,0,182,0,0,0,19,0,107,0,0,0,6,0,22,0,121,0,0,0,121,0,138,0,7,0,61,0,112,0,104,0,245,0,0,0,246,0,190,0,0,0,163,0,68,0,144,0,0,0,208,0,0,0,0,0,0,0,231,0,144,0,0,0,134,0,37,0,1,0,116,0,64,0,144,0,0,0,41,0,128,0,245,0,92,0,232,0,94,0,0,0,122,0,0,0,81,0,126,0,154,0,105,0,65,0,210,0,226,0,157,0,53,0,132,0,25,0,56,0,84,0,5,0,82,0,72,0,176,0,112,0,0,0,221,0,67,0,0,0,199,0,24,0,0,0,0,0,213,0,194,0,0,0,201,0,0,0,126,0,164,0,19,0,0,0,85,0,0,0,38,0,220,0,57,0,1,0,169,0,19,0,80,0,15,0,68,0,162,0,0,0,59,0,0,0,160,0,180,0,185,0,22,0,4,0,89,0,160,0,148,0,90,0,0,0,60,0,0,0,91,0,0,0,242,0,17,0,59,0,63,0,162,0,245,0,4,0,0,0,0,0,229,0,139,0,175,0,18,0,0,0,119,0,56,0,66,0,83,0,117,0,111,0,10,0,116,0,173,0,231,0,230,0,0,0,209,0,44,0,224,0,28,0,122,0,121,0,90,0,83,0,37,0,0,0,248,0,0,0,179,0,198,0,0,0,149,0,101,0,133,0,32,0,132,0,38,0,0,0,33,0,34,0,36,0,97,0,0,0,237,0,0,0,0,0,28,0,23,0,20,0,31,0,0,0,120,0,129,0,42,0,146,0,19,0,0,0,233,0,44,0,14,0,129,0,242,0,74,0,17,0,119,0,247,0,0,0,180,0,12,0,203,0,52,0,54,0,166,0,175,0,115,0,25,0,204,0,232,0,0,0,0,0,0,0,222,0,81,0,42,0,118,0,161,0,136,0,83,0,185,0,58,0,209,0,56,0,99,0,184,0,71,0,52,0,49,0,0,0,100,0,8,0,0,0,199,0,0,0,0,0,46,0,0,0,0,0,9,0,0,0,77,0,251,0,32,0,0,0,26,0,128,0,136,0,200,0,0,0,13,0,56,0,169,0,235,0,142,0,80,0,39,0,55,0,70,0,0,0,46,0,152,0,237,0,13,0,161,0,0,0,0,0,0,0,236,0,94,0,214,0,113,0,78,0,177,0,137,0,159,0,149,0,43,0,118,0,243,0,89,0,146,0,62,0,1,0,0,0,19,0,145,0,140,0,85,0,181,0,234,0,0,0,46,0,97,0,194,0,234,0,0,0,110,0,180,0,0,0,179,0,0,0,86,0,195,0,234,0,193,0,15,0,64,0,205,0,185,0,11,0,204,0,70,0,160,0,0,0,72,0,80,0,28,0,200,0,117,0,169,0,154,0,1,0,244,0,95,0,53,0,23,0,246,0,21,0,224,0,153,0,238,0,250,0,216,0,112,0,82,0,54,0,131,0,159,0,0,0,196,0,206,0,80,0,0,0,0,0,147,0,0,0,173,0,176,0,249,0,124,0,0,0,64,0,218,0,92,0,164,0,199,0,184,0,104,0,49,0,70,0,228,0,77,0,0,0,145,0,0,0,0,0,209,0,63,0,180,0,68,0,21,0,185,0,170,0,160,0,226,0,148,0,101,0,251,0,130,0,228,0,199,0,157,0,164,0,0,0,0,0,49,0,217,0,69,0,22,0,26,0,228,0,5,0,133,0,144,0,101,0,238,0,0,0,219,0,209,0,177,0,40,0,148,0,0,0,196,0,0,0,128,0,154,0,122,0,236,0,0,0,20,0,43,0,126,0,0,0,0,0,198,0,0,0,249,0,146,0,0,0,249,0,0,0,31,0,0,0,245,0,0,0,90,0,250,0,0,0,192,0,0,0,0,0,103,0,25,0,13,0,172,0,30,0,219,0,195,0,39,0,28,0,164,0,0,0,0,0,20,0,239,0,6,0,0,0,197,0,97,0,172,0,0,0,99,0,255,0,52,0,0,0,123,0,18,0,123,0,93,0,89,0,30,0,252,0,0,0,32,0,51,0,157,0,162,0,184,0,8,0,185,0,199,0,231,0,95,0,217,0,193,0,176,0,92,0,0,0,218,0,0,0,247,0,12,0,69,0,149,0,0,0,0,0,68,0,9,0,0,0,240,0,165,0,38,0,66,0,199,0,156,0,10,0,33,0,130,0,125,0,0,0,238,0,0,0,243,0,131,0,251,0,0,0,130,0,115,0,162,0,190,0,0,0,0,0,0,0,243,0,101,0,165,0,222,0,222,0,81,0,0,0,0,0,200,0,150,0,85,0,173,0,113,0,110,0,90,0,62,0,129,0,255,0,122,0,240,0,226,0,210,0,112,0,232,0,128,0,35,0,83,0,0,0,41,0,215,0,201,0,153,0);
signal scenario_full  : scenario_type := (253,31,32,31,7,31,135,31,165,31,9,31,220,31,220,30,220,29,128,31,241,31,209,31,149,31,69,31,69,30,95,31,38,31,108,31,50,31,70,31,144,31,96,31,246,31,72,31,60,31,60,30,60,29,62,31,21,31,21,31,82,31,75,31,75,30,41,31,13,31,235,31,235,30,170,31,178,31,253,31,253,30,33,31,44,31,97,31,96,31,30,31,30,30,249,31,35,31,87,31,124,31,56,31,60,31,203,31,203,30,182,31,182,30,19,31,107,31,107,30,6,31,22,31,121,31,121,30,121,31,138,31,7,31,61,31,112,31,104,31,245,31,245,30,246,31,190,31,190,30,163,31,68,31,144,31,144,30,208,31,208,30,208,29,208,28,231,31,144,31,144,30,134,31,37,31,1,31,116,31,64,31,144,31,144,30,41,31,128,31,245,31,92,31,232,31,94,31,94,30,122,31,122,30,81,31,126,31,154,31,105,31,65,31,210,31,226,31,157,31,53,31,132,31,25,31,56,31,84,31,5,31,82,31,72,31,176,31,112,31,112,30,221,31,67,31,67,30,199,31,24,31,24,30,24,29,213,31,194,31,194,30,201,31,201,30,126,31,164,31,19,31,19,30,85,31,85,30,38,31,220,31,57,31,1,31,169,31,19,31,80,31,15,31,68,31,162,31,162,30,59,31,59,30,160,31,180,31,185,31,22,31,4,31,89,31,160,31,148,31,90,31,90,30,60,31,60,30,91,31,91,30,242,31,17,31,59,31,63,31,162,31,245,31,4,31,4,30,4,29,229,31,139,31,175,31,18,31,18,30,119,31,56,31,66,31,83,31,117,31,111,31,10,31,116,31,173,31,231,31,230,31,230,30,209,31,44,31,224,31,28,31,122,31,121,31,90,31,83,31,37,31,37,30,248,31,248,30,179,31,198,31,198,30,149,31,101,31,133,31,32,31,132,31,38,31,38,30,33,31,34,31,36,31,97,31,97,30,237,31,237,30,237,29,28,31,23,31,20,31,31,31,31,30,120,31,129,31,42,31,146,31,19,31,19,30,233,31,44,31,14,31,129,31,242,31,74,31,17,31,119,31,247,31,247,30,180,31,12,31,203,31,52,31,54,31,166,31,175,31,115,31,25,31,204,31,232,31,232,30,232,29,232,28,222,31,81,31,42,31,118,31,161,31,136,31,83,31,185,31,58,31,209,31,56,31,99,31,184,31,71,31,52,31,49,31,49,30,100,31,8,31,8,30,199,31,199,30,199,29,46,31,46,30,46,29,9,31,9,30,77,31,251,31,32,31,32,30,26,31,128,31,136,31,200,31,200,30,13,31,56,31,169,31,235,31,142,31,80,31,39,31,55,31,70,31,70,30,46,31,152,31,237,31,13,31,161,31,161,30,161,29,161,28,236,31,94,31,214,31,113,31,78,31,177,31,137,31,159,31,149,31,43,31,118,31,243,31,89,31,146,31,62,31,1,31,1,30,19,31,145,31,140,31,85,31,181,31,234,31,234,30,46,31,97,31,194,31,234,31,234,30,110,31,180,31,180,30,179,31,179,30,86,31,195,31,234,31,193,31,15,31,64,31,205,31,185,31,11,31,204,31,70,31,160,31,160,30,72,31,80,31,28,31,200,31,117,31,169,31,154,31,1,31,244,31,95,31,53,31,23,31,246,31,21,31,224,31,153,31,238,31,250,31,216,31,112,31,82,31,54,31,131,31,159,31,159,30,196,31,206,31,80,31,80,30,80,29,147,31,147,30,173,31,176,31,249,31,124,31,124,30,64,31,218,31,92,31,164,31,199,31,184,31,104,31,49,31,70,31,228,31,77,31,77,30,145,31,145,30,145,29,209,31,63,31,180,31,68,31,21,31,185,31,170,31,160,31,226,31,148,31,101,31,251,31,130,31,228,31,199,31,157,31,164,31,164,30,164,29,49,31,217,31,69,31,22,31,26,31,228,31,5,31,133,31,144,31,101,31,238,31,238,30,219,31,209,31,177,31,40,31,148,31,148,30,196,31,196,30,128,31,154,31,122,31,236,31,236,30,20,31,43,31,126,31,126,30,126,29,198,31,198,30,249,31,146,31,146,30,249,31,249,30,31,31,31,30,245,31,245,30,90,31,250,31,250,30,192,31,192,30,192,29,103,31,25,31,13,31,172,31,30,31,219,31,195,31,39,31,28,31,164,31,164,30,164,29,20,31,239,31,6,31,6,30,197,31,97,31,172,31,172,30,99,31,255,31,52,31,52,30,123,31,18,31,123,31,93,31,89,31,30,31,252,31,252,30,32,31,51,31,157,31,162,31,184,31,8,31,185,31,199,31,231,31,95,31,217,31,193,31,176,31,92,31,92,30,218,31,218,30,247,31,12,31,69,31,149,31,149,30,149,29,68,31,9,31,9,30,240,31,165,31,38,31,66,31,199,31,156,31,10,31,33,31,130,31,125,31,125,30,238,31,238,30,243,31,131,31,251,31,251,30,130,31,115,31,162,31,190,31,190,30,190,29,190,28,243,31,101,31,165,31,222,31,222,31,81,31,81,30,81,29,200,31,150,31,85,31,173,31,113,31,110,31,90,31,62,31,129,31,255,31,122,31,240,31,226,31,210,31,112,31,232,31,128,31,35,31,83,31,83,30,41,31,215,31,201,31,153,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
