-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 882;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,139,0,252,0,53,0,98,0,97,0,245,0,0,0,184,0,136,0,197,0,35,0,0,0,33,0,27,0,0,0,0,0,8,0,78,0,0,0,0,0,102,0,32,0,23,0,54,0,104,0,13,0,0,0,0,0,161,0,0,0,0,0,5,0,73,0,243,0,246,0,189,0,101,0,123,0,103,0,85,0,74,0,230,0,0,0,168,0,0,0,221,0,112,0,230,0,127,0,138,0,0,0,24,0,81,0,36,0,0,0,0,0,81,0,0,0,0,0,5,0,127,0,22,0,115,0,85,0,0,0,126,0,0,0,167,0,0,0,0,0,114,0,78,0,163,0,79,0,104,0,21,0,30,0,236,0,238,0,57,0,173,0,22,0,138,0,213,0,167,0,0,0,0,0,0,0,50,0,246,0,61,0,17,0,38,0,69,0,234,0,0,0,90,0,234,0,232,0,184,0,199,0,94,0,0,0,217,0,60,0,75,0,209,0,99,0,50,0,0,0,122,0,64,0,170,0,24,0,135,0,232,0,22,0,97,0,101,0,0,0,83,0,178,0,0,0,213,0,0,0,0,0,0,0,44,0,0,0,0,0,76,0,246,0,177,0,146,0,210,0,212,0,151,0,0,0,136,0,195,0,72,0,38,0,249,0,6,0,41,0,41,0,162,0,203,0,192,0,0,0,0,0,215,0,184,0,238,0,23,0,143,0,240,0,93,0,127,0,158,0,19,0,5,0,161,0,50,0,105,0,80,0,140,0,118,0,0,0,168,0,12,0,40,0,33,0,108,0,151,0,0,0,44,0,105,0,95,0,179,0,95,0,58,0,221,0,64,0,131,0,89,0,17,0,243,0,0,0,216,0,112,0,0,0,226,0,184,0,210,0,167,0,0,0,53,0,41,0,150,0,178,0,36,0,51,0,243,0,128,0,130,0,230,0,151,0,103,0,115,0,77,0,0,0,0,0,149,0,80,0,0,0,33,0,237,0,18,0,2,0,220,0,130,0,163,0,36,0,206,0,113,0,0,0,0,0,20,0,159,0,173,0,37,0,184,0,14,0,34,0,171,0,0,0,0,0,0,0,83,0,22,0,46,0,170,0,0,0,175,0,171,0,188,0,200,0,106,0,0,0,214,0,72,0,224,0,0,0,149,0,194,0,145,0,193,0,39,0,92,0,13,0,24,0,13,0,45,0,0,0,201,0,91,0,17,0,123,0,234,0,0,0,219,0,203,0,0,0,31,0,219,0,173,0,170,0,197,0,0,0,193,0,108,0,0,0,0,0,0,0,169,0,237,0,64,0,235,0,39,0,50,0,52,0,190,0,17,0,7,0,0,0,0,0,171,0,206,0,246,0,90,0,106,0,0,0,10,0,78,0,0,0,160,0,192,0,0,0,17,0,200,0,103,0,28,0,25,0,41,0,151,0,220,0,45,0,84,0,103,0,168,0,0,0,144,0,0,0,205,0,174,0,0,0,230,0,218,0,157,0,0,0,109,0,0,0,229,0,105,0,87,0,227,0,0,0,0,0,224,0,166,0,43,0,12,0,2,0,81,0,0,0,60,0,41,0,60,0,236,0,112,0,57,0,148,0,0,0,178,0,193,0,53,0,128,0,247,0,149,0,0,0,0,0,91,0,38,0,210,0,192,0,118,0,0,0,0,0,108,0,86,0,208,0,50,0,32,0,211,0,0,0,94,0,138,0,159,0,206,0,7,0,41,0,134,0,30,0,250,0,0,0,231,0,167,0,0,0,242,0,224,0,36,0,191,0,153,0,189,0,163,0,247,0,86,0,219,0,0,0,231,0,0,0,207,0,217,0,108,0,29,0,0,0,251,0,27,0,2,0,0,0,5,0,0,0,0,0,102,0,86,0,19,0,138,0,17,0,0,0,4,0,168,0,149,0,56,0,89,0,207,0,41,0,147,0,95,0,243,0,197,0,157,0,122,0,33,0,201,0,0,0,0,0,0,0,92,0,195,0,54,0,36,0,231,0,3,0,222,0,144,0,177,0,140,0,0,0,0,0,221,0,141,0,2,0,232,0,164,0,76,0,220,0,179,0,19,0,179,0,39,0,197,0,194,0,0,0,105,0,208,0,124,0,26,0,143,0,172,0,133,0,55,0,22,0,0,0,0,0,28,0,123,0,100,0,122,0,208,0,161,0,168,0,189,0,37,0,0,0,68,0,0,0,157,0,137,0,0,0,16,0,233,0,150,0,236,0,0,0,0,0,8,0,255,0,0,0,135,0,122,0,232,0,0,0,0,0,0,0,204,0,57,0,225,0,98,0,141,0,163,0,55,0,32,0,0,0,0,0,19,0,0,0,0,0,81,0,177,0,133,0,0,0,0,0,187,0,157,0,200,0,147,0,129,0,0,0,0,0,37,0,188,0,255,0,44,0,126,0,184,0,11,0,106,0,21,0,84,0,184,0,0,0,0,0,190,0,169,0,249,0,0,0,100,0,0,0,207,0,2,0,144,0,140,0,147,0,176,0,93,0,212,0,86,0,22,0,0,0,157,0,114,0,125,0,154,0,39,0,1,0,29,0,235,0,217,0,127,0,160,0,0,0,0,0,75,0,154,0,75,0,249,0,124,0,25,0,98,0,223,0,0,0,238,0,163,0,246,0,0,0,191,0,191,0,0,0,8,0,204,0,120,0,115,0,123,0,0,0,177,0,0,0,0,0,0,0,81,0,0,0,62,0,0,0,236,0,150,0,0,0,0,0,56,0,63,0,63,0,0,0,122,0,205,0,77,0,21,0,82,0,108,0,102,0,242,0,0,0,14,0,81,0,0,0,228,0,23,0,107,0,82,0,14,0,141,0,193,0,93,0,114,0,0,0,209,0,56,0,0,0,199,0,58,0,83,0,65,0,54,0,0,0,44,0,65,0,245,0,106,0,0,0,0,0,0,0,65,0,67,0,115,0,250,0,41,0,41,0,157,0,196,0,0,0,221,0,0,0,202,0,216,0,0,0,57,0,188,0,136,0,237,0,113,0,162,0,147,0,226,0,67,0,229,0,253,0,94,0,0,0,0,0,231,0,68,0,174,0,157,0,130,0,248,0,36,0,0,0,9,0,162,0,86,0,0,0,167,0,218,0,200,0,165,0,52,0,0,0,177,0,172,0,122,0,204,0,100,0,188,0,112,0,159,0,0,0,243,0,0,0,0,0,160,0,244,0,0,0,10,0,237,0,162,0,0,0,0,0,121,0,223,0,20,0,221,0,0,0,126,0,135,0,0,0,125,0,234,0,0,0,195,0,161,0,253,0,45,0,199,0,133,0,252,0,238,0,124,0,32,0,80,0,222,0,210,0,90,0,20,0,119,0,138,0,244,0,0,0,0,0,103,0,55,0,140,0,106,0,0,0,94,0,46,0,179,0,228,0,20,0,61,0,10,0,197,0,20,0,190,0,20,0,0,0,0,0,90,0,78,0,208,0,240,0,8,0,192,0,0,0,42,0,34,0,4,0,0,0,0,0,0,0,131,0,230,0,0,0,143,0,98,0,0,0,210,0,203,0,210,0,38,0,240,0,210,0,130,0,1,0,51,0,70,0,110,0,0,0,57,0,156,0,58,0,0,0,187,0,117,0,186,0,158,0,198,0,0,0,25,0,0,0,46,0,117,0,82,0,0,0,249,0,228,0,211,0,0,0,186,0,0,0,251,0,165,0,117,0,244,0,44,0,254,0,56,0,167,0,123,0,163,0,0,0,203,0,221,0,26,0,0,0,138,0,136,0,97,0,85,0,228,0,242,0,73,0,232,0,17,0,111,0,0,0,184,0,127,0,74,0,1,0,25,0,57,0,121,0,234,0,57,0,121,0,79,0,103,0,68,0,133,0,252,0,191,0,39,0,240,0,0,0,117,0,71,0,182,0,80,0,4,0,0,0,117,0,79,0,94,0,166,0,78,0,153,0,163,0,0,0,0,0,0,0,132,0,125,0,64,0);
signal scenario_full  : scenario_type := (0,0,139,31,252,31,53,31,98,31,97,31,245,31,245,30,184,31,136,31,197,31,35,31,35,30,33,31,27,31,27,30,27,29,8,31,78,31,78,30,78,29,102,31,32,31,23,31,54,31,104,31,13,31,13,30,13,29,161,31,161,30,161,29,5,31,73,31,243,31,246,31,189,31,101,31,123,31,103,31,85,31,74,31,230,31,230,30,168,31,168,30,221,31,112,31,230,31,127,31,138,31,138,30,24,31,81,31,36,31,36,30,36,29,81,31,81,30,81,29,5,31,127,31,22,31,115,31,85,31,85,30,126,31,126,30,167,31,167,30,167,29,114,31,78,31,163,31,79,31,104,31,21,31,30,31,236,31,238,31,57,31,173,31,22,31,138,31,213,31,167,31,167,30,167,29,167,28,50,31,246,31,61,31,17,31,38,31,69,31,234,31,234,30,90,31,234,31,232,31,184,31,199,31,94,31,94,30,217,31,60,31,75,31,209,31,99,31,50,31,50,30,122,31,64,31,170,31,24,31,135,31,232,31,22,31,97,31,101,31,101,30,83,31,178,31,178,30,213,31,213,30,213,29,213,28,44,31,44,30,44,29,76,31,246,31,177,31,146,31,210,31,212,31,151,31,151,30,136,31,195,31,72,31,38,31,249,31,6,31,41,31,41,31,162,31,203,31,192,31,192,30,192,29,215,31,184,31,238,31,23,31,143,31,240,31,93,31,127,31,158,31,19,31,5,31,161,31,50,31,105,31,80,31,140,31,118,31,118,30,168,31,12,31,40,31,33,31,108,31,151,31,151,30,44,31,105,31,95,31,179,31,95,31,58,31,221,31,64,31,131,31,89,31,17,31,243,31,243,30,216,31,112,31,112,30,226,31,184,31,210,31,167,31,167,30,53,31,41,31,150,31,178,31,36,31,51,31,243,31,128,31,130,31,230,31,151,31,103,31,115,31,77,31,77,30,77,29,149,31,80,31,80,30,33,31,237,31,18,31,2,31,220,31,130,31,163,31,36,31,206,31,113,31,113,30,113,29,20,31,159,31,173,31,37,31,184,31,14,31,34,31,171,31,171,30,171,29,171,28,83,31,22,31,46,31,170,31,170,30,175,31,171,31,188,31,200,31,106,31,106,30,214,31,72,31,224,31,224,30,149,31,194,31,145,31,193,31,39,31,92,31,13,31,24,31,13,31,45,31,45,30,201,31,91,31,17,31,123,31,234,31,234,30,219,31,203,31,203,30,31,31,219,31,173,31,170,31,197,31,197,30,193,31,108,31,108,30,108,29,108,28,169,31,237,31,64,31,235,31,39,31,50,31,52,31,190,31,17,31,7,31,7,30,7,29,171,31,206,31,246,31,90,31,106,31,106,30,10,31,78,31,78,30,160,31,192,31,192,30,17,31,200,31,103,31,28,31,25,31,41,31,151,31,220,31,45,31,84,31,103,31,168,31,168,30,144,31,144,30,205,31,174,31,174,30,230,31,218,31,157,31,157,30,109,31,109,30,229,31,105,31,87,31,227,31,227,30,227,29,224,31,166,31,43,31,12,31,2,31,81,31,81,30,60,31,41,31,60,31,236,31,112,31,57,31,148,31,148,30,178,31,193,31,53,31,128,31,247,31,149,31,149,30,149,29,91,31,38,31,210,31,192,31,118,31,118,30,118,29,108,31,86,31,208,31,50,31,32,31,211,31,211,30,94,31,138,31,159,31,206,31,7,31,41,31,134,31,30,31,250,31,250,30,231,31,167,31,167,30,242,31,224,31,36,31,191,31,153,31,189,31,163,31,247,31,86,31,219,31,219,30,231,31,231,30,207,31,217,31,108,31,29,31,29,30,251,31,27,31,2,31,2,30,5,31,5,30,5,29,102,31,86,31,19,31,138,31,17,31,17,30,4,31,168,31,149,31,56,31,89,31,207,31,41,31,147,31,95,31,243,31,197,31,157,31,122,31,33,31,201,31,201,30,201,29,201,28,92,31,195,31,54,31,36,31,231,31,3,31,222,31,144,31,177,31,140,31,140,30,140,29,221,31,141,31,2,31,232,31,164,31,76,31,220,31,179,31,19,31,179,31,39,31,197,31,194,31,194,30,105,31,208,31,124,31,26,31,143,31,172,31,133,31,55,31,22,31,22,30,22,29,28,31,123,31,100,31,122,31,208,31,161,31,168,31,189,31,37,31,37,30,68,31,68,30,157,31,137,31,137,30,16,31,233,31,150,31,236,31,236,30,236,29,8,31,255,31,255,30,135,31,122,31,232,31,232,30,232,29,232,28,204,31,57,31,225,31,98,31,141,31,163,31,55,31,32,31,32,30,32,29,19,31,19,30,19,29,81,31,177,31,133,31,133,30,133,29,187,31,157,31,200,31,147,31,129,31,129,30,129,29,37,31,188,31,255,31,44,31,126,31,184,31,11,31,106,31,21,31,84,31,184,31,184,30,184,29,190,31,169,31,249,31,249,30,100,31,100,30,207,31,2,31,144,31,140,31,147,31,176,31,93,31,212,31,86,31,22,31,22,30,157,31,114,31,125,31,154,31,39,31,1,31,29,31,235,31,217,31,127,31,160,31,160,30,160,29,75,31,154,31,75,31,249,31,124,31,25,31,98,31,223,31,223,30,238,31,163,31,246,31,246,30,191,31,191,31,191,30,8,31,204,31,120,31,115,31,123,31,123,30,177,31,177,30,177,29,177,28,81,31,81,30,62,31,62,30,236,31,150,31,150,30,150,29,56,31,63,31,63,31,63,30,122,31,205,31,77,31,21,31,82,31,108,31,102,31,242,31,242,30,14,31,81,31,81,30,228,31,23,31,107,31,82,31,14,31,141,31,193,31,93,31,114,31,114,30,209,31,56,31,56,30,199,31,58,31,83,31,65,31,54,31,54,30,44,31,65,31,245,31,106,31,106,30,106,29,106,28,65,31,67,31,115,31,250,31,41,31,41,31,157,31,196,31,196,30,221,31,221,30,202,31,216,31,216,30,57,31,188,31,136,31,237,31,113,31,162,31,147,31,226,31,67,31,229,31,253,31,94,31,94,30,94,29,231,31,68,31,174,31,157,31,130,31,248,31,36,31,36,30,9,31,162,31,86,31,86,30,167,31,218,31,200,31,165,31,52,31,52,30,177,31,172,31,122,31,204,31,100,31,188,31,112,31,159,31,159,30,243,31,243,30,243,29,160,31,244,31,244,30,10,31,237,31,162,31,162,30,162,29,121,31,223,31,20,31,221,31,221,30,126,31,135,31,135,30,125,31,234,31,234,30,195,31,161,31,253,31,45,31,199,31,133,31,252,31,238,31,124,31,32,31,80,31,222,31,210,31,90,31,20,31,119,31,138,31,244,31,244,30,244,29,103,31,55,31,140,31,106,31,106,30,94,31,46,31,179,31,228,31,20,31,61,31,10,31,197,31,20,31,190,31,20,31,20,30,20,29,90,31,78,31,208,31,240,31,8,31,192,31,192,30,42,31,34,31,4,31,4,30,4,29,4,28,131,31,230,31,230,30,143,31,98,31,98,30,210,31,203,31,210,31,38,31,240,31,210,31,130,31,1,31,51,31,70,31,110,31,110,30,57,31,156,31,58,31,58,30,187,31,117,31,186,31,158,31,198,31,198,30,25,31,25,30,46,31,117,31,82,31,82,30,249,31,228,31,211,31,211,30,186,31,186,30,251,31,165,31,117,31,244,31,44,31,254,31,56,31,167,31,123,31,163,31,163,30,203,31,221,31,26,31,26,30,138,31,136,31,97,31,85,31,228,31,242,31,73,31,232,31,17,31,111,31,111,30,184,31,127,31,74,31,1,31,25,31,57,31,121,31,234,31,57,31,121,31,79,31,103,31,68,31,133,31,252,31,191,31,39,31,240,31,240,30,117,31,71,31,182,31,80,31,4,31,4,30,117,31,79,31,94,31,166,31,78,31,153,31,163,31,163,30,163,29,163,28,132,31,125,31,64,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
