-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_567 is
end project_tb_567;

architecture project_tb_arch_567 of project_tb_567 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 771;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (239,0,153,0,53,0,116,0,232,0,13,0,56,0,0,0,38,0,172,0,16,0,0,0,0,0,166,0,192,0,156,0,170,0,165,0,133,0,204,0,132,0,39,0,121,0,131,0,146,0,0,0,217,0,211,0,249,0,225,0,17,0,221,0,206,0,19,0,254,0,0,0,74,0,81,0,174,0,86,0,93,0,146,0,32,0,48,0,163,0,220,0,69,0,140,0,231,0,43,0,40,0,65,0,148,0,129,0,160,0,189,0,109,0,67,0,5,0,47,0,25,0,208,0,182,0,209,0,29,0,177,0,0,0,81,0,0,0,232,0,210,0,0,0,52,0,0,0,228,0,252,0,0,0,0,0,166,0,22,0,189,0,52,0,221,0,20,0,21,0,0,0,222,0,194,0,0,0,89,0,137,0,241,0,0,0,227,0,69,0,168,0,0,0,14,0,118,0,143,0,0,0,122,0,202,0,99,0,173,0,0,0,38,0,57,0,0,0,0,0,106,0,120,0,190,0,92,0,201,0,190,0,202,0,128,0,197,0,45,0,0,0,0,0,153,0,230,0,0,0,0,0,102,0,0,0,180,0,129,0,223,0,103,0,0,0,0,0,122,0,150,0,77,0,128,0,200,0,14,0,84,0,0,0,94,0,90,0,0,0,248,0,0,0,99,0,143,0,246,0,38,0,0,0,43,0,51,0,130,0,82,0,218,0,104,0,0,0,251,0,107,0,0,0,64,0,0,0,0,0,0,0,219,0,213,0,178,0,52,0,148,0,0,0,92,0,106,0,0,0,90,0,115,0,185,0,119,0,49,0,176,0,244,0,176,0,0,0,239,0,130,0,232,0,96,0,201,0,174,0,74,0,254,0,138,0,114,0,157,0,171,0,170,0,64,0,242,0,35,0,213,0,156,0,192,0,129,0,0,0,224,0,6,0,95,0,120,0,165,0,86,0,0,0,0,0,230,0,29,0,0,0,219,0,8,0,251,0,0,0,81,0,103,0,103,0,7,0,164,0,32,0,0,0,0,0,163,0,0,0,0,0,20,0,89,0,186,0,117,0,0,0,244,0,167,0,192,0,201,0,218,0,102,0,231,0,186,0,74,0,125,0,0,0,163,0,0,0,47,0,0,0,71,0,231,0,83,0,247,0,0,0,163,0,219,0,154,0,67,0,242,0,0,0,98,0,152,0,41,0,0,0,80,0,149,0,63,0,185,0,0,0,0,0,167,0,162,0,170,0,167,0,0,0,0,0,179,0,115,0,0,0,127,0,249,0,175,0,4,0,176,0,3,0,140,0,0,0,1,0,0,0,212,0,108,0,10,0,184,0,27,0,156,0,0,0,0,0,0,0,46,0,230,0,22,0,218,0,0,0,0,0,183,0,0,0,0,0,200,0,196,0,60,0,36,0,59,0,0,0,243,0,63,0,175,0,0,0,46,0,146,0,54,0,147,0,85,0,250,0,238,0,140,0,226,0,0,0,224,0,237,0,44,0,222,0,0,0,174,0,218,0,208,0,77,0,187,0,251,0,0,0,147,0,116,0,157,0,28,0,0,0,86,0,88,0,128,0,124,0,92,0,53,0,106,0,98,0,0,0,243,0,37,0,241,0,109,0,171,0,164,0,113,0,117,0,87,0,57,0,78,0,134,0,88,0,137,0,196,0,0,0,84,0,29,0,0,0,120,0,56,0,184,0,135,0,55,0,192,0,37,0,0,0,88,0,170,0,155,0,48,0,0,0,38,0,66,0,16,0,14,0,0,0,150,0,211,0,223,0,139,0,228,0,228,0,84,0,3,0,119,0,185,0,0,0,0,0,43,0,0,0,155,0,117,0,0,0,70,0,167,0,194,0,99,0,184,0,0,0,0,0,79,0,158,0,109,0,9,0,68,0,0,0,0,0,13,0,11,0,0,0,8,0,234,0,144,0,26,0,111,0,51,0,0,0,234,0,47,0,238,0,143,0,147,0,215,0,4,0,17,0,0,0,117,0,244,0,233,0,0,0,116,0,6,0,79,0,232,0,0,0,0,0,183,0,162,0,213,0,126,0,122,0,76,0,181,0,212,0,0,0,63,0,13,0,242,0,6,0,160,0,215,0,93,0,91,0,20,0,143,0,87,0,0,0,214,0,6,0,118,0,199,0,42,0,102,0,65,0,72,0,89,0,205,0,205,0,73,0,0,0,101,0,214,0,105,0,166,0,196,0,136,0,244,0,87,0,0,0,124,0,182,0,91,0,109,0,64,0,0,0,0,0,187,0,215,0,12,0,234,0,190,0,177,0,138,0,0,0,163,0,21,0,76,0,56,0,172,0,235,0,28,0,63,0,104,0,0,0,5,0,21,0,0,0,92,0,117,0,50,0,100,0,0,0,97,0,98,0,13,0,68,0,0,0,86,0,114,0,204,0,0,0,213,0,26,0,0,0,76,0,193,0,0,0,84,0,13,0,41,0,0,0,0,0,93,0,110,0,69,0,40,0,202,0,45,0,244,0,0,0,149,0,111,0,108,0,0,0,38,0,0,0,0,0,164,0,97,0,0,0,0,0,114,0,146,0,0,0,9,0,145,0,101,0,73,0,187,0,249,0,248,0,0,0,65,0,69,0,0,0,210,0,41,0,235,0,173,0,0,0,99,0,66,0,4,0,193,0,201,0,170,0,40,0,147,0,88,0,217,0,44,0,208,0,0,0,199,0,117,0,1,0,105,0,91,0,134,0,83,0,253,0,0,0,93,0,137,0,235,0,176,0,19,0,0,0,249,0,205,0,113,0,22,0,251,0,215,0,177,0,173,0,0,0,41,0,169,0,163,0,239,0,180,0,235,0,0,0,207,0,220,0,0,0,19,0,191,0,153,0,141,0,102,0,57,0,216,0,71,0,33,0,0,0,201,0,74,0,25,0,53,0,241,0,53,0,213,0,0,0,0,0,18,0,144,0,8,0,249,0,208,0,65,0,237,0,234,0,46,0,53,0,52,0,121,0,68,0,65,0,187,0,0,0,171,0,166,0,0,0,193,0,0,0,202,0,133,0,0,0,0,0,232,0,183,0,211,0,76,0,0,0,177,0,17,0,252,0,92,0,70,0,69,0,86,0,253,0,189,0,136,0,35,0,22,0,0,0,253,0,117,0,0,0,41,0,122,0,38,0,139,0,7,0,179,0,200,0,0,0,156,0,0,0,207,0,193,0,0,0,164,0,0,0,0,0,0,0,0,0,112,0,223,0,0,0,0,0,0,0,119,0,229,0,61,0,69,0,0,0,183,0,0,0,18,0,105,0,44,0,0,0,199,0,164,0,206,0,110,0,186,0,0,0,227,0,0,0,157,0,60,0,10,0,23,0,130,0,165,0,211,0,21,0,212,0,114,0,95,0,55,0,217,0,0,0,0,0,127,0,41,0,1,0,120,0,238,0,98,0,241,0,167,0,0,0,80,0,100,0,166,0,68,0,0,0,0,0,165,0);
signal scenario_full  : scenario_type := (239,31,153,31,53,31,116,31,232,31,13,31,56,31,56,30,38,31,172,31,16,31,16,30,16,29,166,31,192,31,156,31,170,31,165,31,133,31,204,31,132,31,39,31,121,31,131,31,146,31,146,30,217,31,211,31,249,31,225,31,17,31,221,31,206,31,19,31,254,31,254,30,74,31,81,31,174,31,86,31,93,31,146,31,32,31,48,31,163,31,220,31,69,31,140,31,231,31,43,31,40,31,65,31,148,31,129,31,160,31,189,31,109,31,67,31,5,31,47,31,25,31,208,31,182,31,209,31,29,31,177,31,177,30,81,31,81,30,232,31,210,31,210,30,52,31,52,30,228,31,252,31,252,30,252,29,166,31,22,31,189,31,52,31,221,31,20,31,21,31,21,30,222,31,194,31,194,30,89,31,137,31,241,31,241,30,227,31,69,31,168,31,168,30,14,31,118,31,143,31,143,30,122,31,202,31,99,31,173,31,173,30,38,31,57,31,57,30,57,29,106,31,120,31,190,31,92,31,201,31,190,31,202,31,128,31,197,31,45,31,45,30,45,29,153,31,230,31,230,30,230,29,102,31,102,30,180,31,129,31,223,31,103,31,103,30,103,29,122,31,150,31,77,31,128,31,200,31,14,31,84,31,84,30,94,31,90,31,90,30,248,31,248,30,99,31,143,31,246,31,38,31,38,30,43,31,51,31,130,31,82,31,218,31,104,31,104,30,251,31,107,31,107,30,64,31,64,30,64,29,64,28,219,31,213,31,178,31,52,31,148,31,148,30,92,31,106,31,106,30,90,31,115,31,185,31,119,31,49,31,176,31,244,31,176,31,176,30,239,31,130,31,232,31,96,31,201,31,174,31,74,31,254,31,138,31,114,31,157,31,171,31,170,31,64,31,242,31,35,31,213,31,156,31,192,31,129,31,129,30,224,31,6,31,95,31,120,31,165,31,86,31,86,30,86,29,230,31,29,31,29,30,219,31,8,31,251,31,251,30,81,31,103,31,103,31,7,31,164,31,32,31,32,30,32,29,163,31,163,30,163,29,20,31,89,31,186,31,117,31,117,30,244,31,167,31,192,31,201,31,218,31,102,31,231,31,186,31,74,31,125,31,125,30,163,31,163,30,47,31,47,30,71,31,231,31,83,31,247,31,247,30,163,31,219,31,154,31,67,31,242,31,242,30,98,31,152,31,41,31,41,30,80,31,149,31,63,31,185,31,185,30,185,29,167,31,162,31,170,31,167,31,167,30,167,29,179,31,115,31,115,30,127,31,249,31,175,31,4,31,176,31,3,31,140,31,140,30,1,31,1,30,212,31,108,31,10,31,184,31,27,31,156,31,156,30,156,29,156,28,46,31,230,31,22,31,218,31,218,30,218,29,183,31,183,30,183,29,200,31,196,31,60,31,36,31,59,31,59,30,243,31,63,31,175,31,175,30,46,31,146,31,54,31,147,31,85,31,250,31,238,31,140,31,226,31,226,30,224,31,237,31,44,31,222,31,222,30,174,31,218,31,208,31,77,31,187,31,251,31,251,30,147,31,116,31,157,31,28,31,28,30,86,31,88,31,128,31,124,31,92,31,53,31,106,31,98,31,98,30,243,31,37,31,241,31,109,31,171,31,164,31,113,31,117,31,87,31,57,31,78,31,134,31,88,31,137,31,196,31,196,30,84,31,29,31,29,30,120,31,56,31,184,31,135,31,55,31,192,31,37,31,37,30,88,31,170,31,155,31,48,31,48,30,38,31,66,31,16,31,14,31,14,30,150,31,211,31,223,31,139,31,228,31,228,31,84,31,3,31,119,31,185,31,185,30,185,29,43,31,43,30,155,31,117,31,117,30,70,31,167,31,194,31,99,31,184,31,184,30,184,29,79,31,158,31,109,31,9,31,68,31,68,30,68,29,13,31,11,31,11,30,8,31,234,31,144,31,26,31,111,31,51,31,51,30,234,31,47,31,238,31,143,31,147,31,215,31,4,31,17,31,17,30,117,31,244,31,233,31,233,30,116,31,6,31,79,31,232,31,232,30,232,29,183,31,162,31,213,31,126,31,122,31,76,31,181,31,212,31,212,30,63,31,13,31,242,31,6,31,160,31,215,31,93,31,91,31,20,31,143,31,87,31,87,30,214,31,6,31,118,31,199,31,42,31,102,31,65,31,72,31,89,31,205,31,205,31,73,31,73,30,101,31,214,31,105,31,166,31,196,31,136,31,244,31,87,31,87,30,124,31,182,31,91,31,109,31,64,31,64,30,64,29,187,31,215,31,12,31,234,31,190,31,177,31,138,31,138,30,163,31,21,31,76,31,56,31,172,31,235,31,28,31,63,31,104,31,104,30,5,31,21,31,21,30,92,31,117,31,50,31,100,31,100,30,97,31,98,31,13,31,68,31,68,30,86,31,114,31,204,31,204,30,213,31,26,31,26,30,76,31,193,31,193,30,84,31,13,31,41,31,41,30,41,29,93,31,110,31,69,31,40,31,202,31,45,31,244,31,244,30,149,31,111,31,108,31,108,30,38,31,38,30,38,29,164,31,97,31,97,30,97,29,114,31,146,31,146,30,9,31,145,31,101,31,73,31,187,31,249,31,248,31,248,30,65,31,69,31,69,30,210,31,41,31,235,31,173,31,173,30,99,31,66,31,4,31,193,31,201,31,170,31,40,31,147,31,88,31,217,31,44,31,208,31,208,30,199,31,117,31,1,31,105,31,91,31,134,31,83,31,253,31,253,30,93,31,137,31,235,31,176,31,19,31,19,30,249,31,205,31,113,31,22,31,251,31,215,31,177,31,173,31,173,30,41,31,169,31,163,31,239,31,180,31,235,31,235,30,207,31,220,31,220,30,19,31,191,31,153,31,141,31,102,31,57,31,216,31,71,31,33,31,33,30,201,31,74,31,25,31,53,31,241,31,53,31,213,31,213,30,213,29,18,31,144,31,8,31,249,31,208,31,65,31,237,31,234,31,46,31,53,31,52,31,121,31,68,31,65,31,187,31,187,30,171,31,166,31,166,30,193,31,193,30,202,31,133,31,133,30,133,29,232,31,183,31,211,31,76,31,76,30,177,31,17,31,252,31,92,31,70,31,69,31,86,31,253,31,189,31,136,31,35,31,22,31,22,30,253,31,117,31,117,30,41,31,122,31,38,31,139,31,7,31,179,31,200,31,200,30,156,31,156,30,207,31,193,31,193,30,164,31,164,30,164,29,164,28,164,27,112,31,223,31,223,30,223,29,223,28,119,31,229,31,61,31,69,31,69,30,183,31,183,30,18,31,105,31,44,31,44,30,199,31,164,31,206,31,110,31,186,31,186,30,227,31,227,30,157,31,60,31,10,31,23,31,130,31,165,31,211,31,21,31,212,31,114,31,95,31,55,31,217,31,217,30,217,29,127,31,41,31,1,31,120,31,238,31,98,31,241,31,167,31,167,30,80,31,100,31,166,31,68,31,68,30,68,29,165,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
