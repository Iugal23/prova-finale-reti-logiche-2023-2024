-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_143 is
end project_tb_143;

architecture project_tb_arch_143 of project_tb_143 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 172;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,216,0,107,0,180,0,141,0,0,0,0,0,168,0,229,0,6,0,217,0,240,0,253,0,247,0,28,0,134,0,144,0,37,0,163,0,219,0,197,0,232,0,199,0,252,0,90,0,81,0,239,0,247,0,83,0,192,0,50,0,0,0,120,0,87,0,233,0,47,0,184,0,54,0,160,0,0,0,245,0,186,0,122,0,0,0,166,0,4,0,119,0,0,0,160,0,94,0,144,0,229,0,36,0,0,0,35,0,76,0,139,0,66,0,127,0,203,0,27,0,76,0,241,0,158,0,117,0,144,0,209,0,25,0,129,0,0,0,0,0,238,0,183,0,99,0,0,0,0,0,34,0,191,0,156,0,169,0,217,0,50,0,96,0,0,0,86,0,200,0,1,0,41,0,23,0,0,0,211,0,195,0,93,0,204,0,253,0,0,0,54,0,0,0,168,0,251,0,79,0,195,0,157,0,78,0,0,0,47,0,0,0,0,0,90,0,161,0,221,0,16,0,0,0,0,0,85,0,0,0,71,0,224,0,169,0,156,0,94,0,16,0,106,0,155,0,0,0,164,0,0,0,37,0,150,0,0,0,235,0,80,0,209,0,21,0,77,0,191,0,70,0,85,0,225,0,90,0,23,0,2,0,0,0,153,0,222,0,9,0,0,0,123,0,0,0,168,0,137,0,150,0,99,0,69,0,199,0,121,0,174,0,125,0,0,0,0,0,43,0,216,0,193,0,0,0,44,0,7,0,28,0,6,0,141,0,0,0,99,0,0,0);
signal scenario_full  : scenario_type := (0,0,216,31,107,31,180,31,141,31,141,30,141,29,168,31,229,31,6,31,217,31,240,31,253,31,247,31,28,31,134,31,144,31,37,31,163,31,219,31,197,31,232,31,199,31,252,31,90,31,81,31,239,31,247,31,83,31,192,31,50,31,50,30,120,31,87,31,233,31,47,31,184,31,54,31,160,31,160,30,245,31,186,31,122,31,122,30,166,31,4,31,119,31,119,30,160,31,94,31,144,31,229,31,36,31,36,30,35,31,76,31,139,31,66,31,127,31,203,31,27,31,76,31,241,31,158,31,117,31,144,31,209,31,25,31,129,31,129,30,129,29,238,31,183,31,99,31,99,30,99,29,34,31,191,31,156,31,169,31,217,31,50,31,96,31,96,30,86,31,200,31,1,31,41,31,23,31,23,30,211,31,195,31,93,31,204,31,253,31,253,30,54,31,54,30,168,31,251,31,79,31,195,31,157,31,78,31,78,30,47,31,47,30,47,29,90,31,161,31,221,31,16,31,16,30,16,29,85,31,85,30,71,31,224,31,169,31,156,31,94,31,16,31,106,31,155,31,155,30,164,31,164,30,37,31,150,31,150,30,235,31,80,31,209,31,21,31,77,31,191,31,70,31,85,31,225,31,90,31,23,31,2,31,2,30,153,31,222,31,9,31,9,30,123,31,123,30,168,31,137,31,150,31,99,31,69,31,199,31,121,31,174,31,125,31,125,30,125,29,43,31,216,31,193,31,193,30,44,31,7,31,28,31,6,31,141,31,141,30,99,31,99,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
