-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 652;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (61,0,181,0,0,0,0,0,0,0,191,0,28,0,133,0,65,0,0,0,30,0,0,0,111,0,0,0,157,0,97,0,0,0,19,0,0,0,242,0,33,0,110,0,0,0,159,0,245,0,38,0,250,0,120,0,99,0,178,0,0,0,28,0,177,0,85,0,162,0,217,0,232,0,205,0,78,0,229,0,166,0,141,0,75,0,0,0,68,0,141,0,0,0,77,0,69,0,170,0,99,0,120,0,7,0,84,0,0,0,72,0,0,0,0,0,183,0,22,0,238,0,24,0,199,0,0,0,148,0,136,0,87,0,0,0,32,0,0,0,63,0,0,0,6,0,207,0,0,0,58,0,177,0,225,0,157,0,17,0,24,0,77,0,220,0,0,0,203,0,190,0,56,0,0,0,32,0,200,0,188,0,26,0,59,0,0,0,244,0,145,0,185,0,20,0,63,0,202,0,28,0,0,0,123,0,23,0,174,0,157,0,250,0,0,0,107,0,197,0,0,0,41,0,234,0,137,0,0,0,10,0,76,0,168,0,204,0,0,0,88,0,239,0,0,0,122,0,0,0,104,0,25,0,85,0,186,0,99,0,146,0,205,0,131,0,56,0,153,0,5,0,252,0,67,0,234,0,98,0,228,0,191,0,0,0,200,0,0,0,128,0,117,0,0,0,209,0,28,0,20,0,0,0,0,0,224,0,32,0,205,0,248,0,0,0,17,0,162,0,111,0,0,0,0,0,249,0,0,0,0,0,78,0,32,0,0,0,110,0,234,0,0,0,39,0,156,0,187,0,0,0,241,0,249,0,202,0,52,0,148,0,211,0,34,0,66,0,0,0,0,0,0,0,237,0,187,0,50,0,0,0,0,0,149,0,0,0,170,0,254,0,140,0,134,0,232,0,0,0,16,0,247,0,0,0,80,0,0,0,2,0,94,0,40,0,115,0,20,0,0,0,111,0,0,0,143,0,211,0,0,0,174,0,58,0,114,0,222,0,47,0,0,0,130,0,0,0,0,0,65,0,148,0,0,0,135,0,184,0,11,0,107,0,232,0,169,0,0,0,0,0,134,0,164,0,28,0,0,0,64,0,35,0,255,0,128,0,0,0,192,0,162,0,148,0,85,0,241,0,250,0,75,0,10,0,217,0,0,0,0,0,23,0,0,0,0,0,211,0,67,0,0,0,0,0,238,0,197,0,0,0,202,0,225,0,0,0,45,0,140,0,223,0,202,0,0,0,102,0,198,0,0,0,125,0,0,0,22,0,0,0,157,0,249,0,0,0,225,0,168,0,33,0,223,0,55,0,69,0,91,0,145,0,196,0,54,0,0,0,20,0,116,0,103,0,237,0,84,0,49,0,0,0,175,0,80,0,170,0,140,0,129,0,240,0,16,0,0,0,0,0,0,0,123,0,80,0,149,0,4,0,0,0,0,0,66,0,12,0,241,0,0,0,95,0,0,0,97,0,168,0,120,0,27,0,164,0,0,0,0,0,88,0,0,0,226,0,227,0,101,0,196,0,194,0,216,0,207,0,124,0,98,0,0,0,118,0,169,0,159,0,58,0,100,0,140,0,246,0,255,0,0,0,0,0,161,0,153,0,99,0,76,0,0,0,180,0,2,0,210,0,226,0,0,0,85,0,23,0,241,0,58,0,0,0,77,0,185,0,181,0,55,0,165,0,10,0,92,0,222,0,123,0,197,0,0,0,150,0,242,0,0,0,52,0,131,0,49,0,89,0,17,0,37,0,121,0,45,0,0,0,41,0,166,0,175,0,71,0,232,0,18,0,82,0,224,0,229,0,0,0,128,0,89,0,186,0,180,0,80,0,184,0,66,0,0,0,55,0,169,0,98,0,210,0,0,0,252,0,82,0,55,0,19,0,0,0,0,0,2,0,142,0,54,0,193,0,187,0,0,0,0,0,0,0,81,0,0,0,52,0,10,0,154,0,132,0,38,0,63,0,25,0,0,0,0,0,66,0,227,0,112,0,92,0,176,0,196,0,0,0,246,0,113,0,206,0,90,0,125,0,0,0,161,0,182,0,115,0,80,0,25,0,126,0,155,0,75,0,167,0,67,0,0,0,148,0,149,0,0,0,186,0,170,0,156,0,34,0,57,0,221,0,104,0,97,0,105,0,0,0,218,0,16,0,22,0,254,0,187,0,21,0,6,0,0,0,23,0,130,0,80,0,84,0,0,0,186,0,167,0,96,0,107,0,232,0,198,0,89,0,171,0,0,0,105,0,9,0,101,0,167,0,239,0,30,0,179,0,96,0,192,0,127,0,198,0,30,0,160,0,0,0,237,0,229,0,209,0,107,0,0,0,120,0,205,0,101,0,128,0,0,0,223,0,228,0,19,0,0,0,137,0,0,0,0,0,175,0,166,0,233,0,189,0,136,0,201,0,146,0,134,0,226,0,239,0,0,0,243,0,153,0,0,0,100,0,0,0,113,0,223,0,0,0,228,0,147,0,73,0,63,0,87,0,75,0,82,0,0,0,0,0,0,0,0,0,29,0,97,0,159,0,0,0,119,0,74,0,247,0,135,0,17,0,191,0,255,0,39,0,220,0,76,0,122,0,118,0,29,0,229,0,125,0,46,0,121,0,0,0,125,0,0,0,241,0,233,0,228,0,55,0,44,0,230,0,244,0,0,0,64,0,88,0,89,0,224,0,54,0,193,0,170,0,29,0,107,0,0,0,153,0,180,0,220,0,53,0,30,0,48,0,0,0,0,0,226,0,61,0,18,0,168,0,230,0,128,0,104,0,138,0,245,0,199,0,226,0,12,0,0,0,0,0,0,0,174,0,0,0,17,0,0,0,0,0,200,0,0,0,108,0,117,0,0,0,50,0,19,0,61,0,33,0,64,0,30,0,0,0,76,0,209,0,0,0,13,0,102,0,79,0,184,0,163,0,128,0,86,0,0,0);
signal scenario_full  : scenario_type := (61,31,181,31,181,30,181,29,181,28,191,31,28,31,133,31,65,31,65,30,30,31,30,30,111,31,111,30,157,31,97,31,97,30,19,31,19,30,242,31,33,31,110,31,110,30,159,31,245,31,38,31,250,31,120,31,99,31,178,31,178,30,28,31,177,31,85,31,162,31,217,31,232,31,205,31,78,31,229,31,166,31,141,31,75,31,75,30,68,31,141,31,141,30,77,31,69,31,170,31,99,31,120,31,7,31,84,31,84,30,72,31,72,30,72,29,183,31,22,31,238,31,24,31,199,31,199,30,148,31,136,31,87,31,87,30,32,31,32,30,63,31,63,30,6,31,207,31,207,30,58,31,177,31,225,31,157,31,17,31,24,31,77,31,220,31,220,30,203,31,190,31,56,31,56,30,32,31,200,31,188,31,26,31,59,31,59,30,244,31,145,31,185,31,20,31,63,31,202,31,28,31,28,30,123,31,23,31,174,31,157,31,250,31,250,30,107,31,197,31,197,30,41,31,234,31,137,31,137,30,10,31,76,31,168,31,204,31,204,30,88,31,239,31,239,30,122,31,122,30,104,31,25,31,85,31,186,31,99,31,146,31,205,31,131,31,56,31,153,31,5,31,252,31,67,31,234,31,98,31,228,31,191,31,191,30,200,31,200,30,128,31,117,31,117,30,209,31,28,31,20,31,20,30,20,29,224,31,32,31,205,31,248,31,248,30,17,31,162,31,111,31,111,30,111,29,249,31,249,30,249,29,78,31,32,31,32,30,110,31,234,31,234,30,39,31,156,31,187,31,187,30,241,31,249,31,202,31,52,31,148,31,211,31,34,31,66,31,66,30,66,29,66,28,237,31,187,31,50,31,50,30,50,29,149,31,149,30,170,31,254,31,140,31,134,31,232,31,232,30,16,31,247,31,247,30,80,31,80,30,2,31,94,31,40,31,115,31,20,31,20,30,111,31,111,30,143,31,211,31,211,30,174,31,58,31,114,31,222,31,47,31,47,30,130,31,130,30,130,29,65,31,148,31,148,30,135,31,184,31,11,31,107,31,232,31,169,31,169,30,169,29,134,31,164,31,28,31,28,30,64,31,35,31,255,31,128,31,128,30,192,31,162,31,148,31,85,31,241,31,250,31,75,31,10,31,217,31,217,30,217,29,23,31,23,30,23,29,211,31,67,31,67,30,67,29,238,31,197,31,197,30,202,31,225,31,225,30,45,31,140,31,223,31,202,31,202,30,102,31,198,31,198,30,125,31,125,30,22,31,22,30,157,31,249,31,249,30,225,31,168,31,33,31,223,31,55,31,69,31,91,31,145,31,196,31,54,31,54,30,20,31,116,31,103,31,237,31,84,31,49,31,49,30,175,31,80,31,170,31,140,31,129,31,240,31,16,31,16,30,16,29,16,28,123,31,80,31,149,31,4,31,4,30,4,29,66,31,12,31,241,31,241,30,95,31,95,30,97,31,168,31,120,31,27,31,164,31,164,30,164,29,88,31,88,30,226,31,227,31,101,31,196,31,194,31,216,31,207,31,124,31,98,31,98,30,118,31,169,31,159,31,58,31,100,31,140,31,246,31,255,31,255,30,255,29,161,31,153,31,99,31,76,31,76,30,180,31,2,31,210,31,226,31,226,30,85,31,23,31,241,31,58,31,58,30,77,31,185,31,181,31,55,31,165,31,10,31,92,31,222,31,123,31,197,31,197,30,150,31,242,31,242,30,52,31,131,31,49,31,89,31,17,31,37,31,121,31,45,31,45,30,41,31,166,31,175,31,71,31,232,31,18,31,82,31,224,31,229,31,229,30,128,31,89,31,186,31,180,31,80,31,184,31,66,31,66,30,55,31,169,31,98,31,210,31,210,30,252,31,82,31,55,31,19,31,19,30,19,29,2,31,142,31,54,31,193,31,187,31,187,30,187,29,187,28,81,31,81,30,52,31,10,31,154,31,132,31,38,31,63,31,25,31,25,30,25,29,66,31,227,31,112,31,92,31,176,31,196,31,196,30,246,31,113,31,206,31,90,31,125,31,125,30,161,31,182,31,115,31,80,31,25,31,126,31,155,31,75,31,167,31,67,31,67,30,148,31,149,31,149,30,186,31,170,31,156,31,34,31,57,31,221,31,104,31,97,31,105,31,105,30,218,31,16,31,22,31,254,31,187,31,21,31,6,31,6,30,23,31,130,31,80,31,84,31,84,30,186,31,167,31,96,31,107,31,232,31,198,31,89,31,171,31,171,30,105,31,9,31,101,31,167,31,239,31,30,31,179,31,96,31,192,31,127,31,198,31,30,31,160,31,160,30,237,31,229,31,209,31,107,31,107,30,120,31,205,31,101,31,128,31,128,30,223,31,228,31,19,31,19,30,137,31,137,30,137,29,175,31,166,31,233,31,189,31,136,31,201,31,146,31,134,31,226,31,239,31,239,30,243,31,153,31,153,30,100,31,100,30,113,31,223,31,223,30,228,31,147,31,73,31,63,31,87,31,75,31,82,31,82,30,82,29,82,28,82,27,29,31,97,31,159,31,159,30,119,31,74,31,247,31,135,31,17,31,191,31,255,31,39,31,220,31,76,31,122,31,118,31,29,31,229,31,125,31,46,31,121,31,121,30,125,31,125,30,241,31,233,31,228,31,55,31,44,31,230,31,244,31,244,30,64,31,88,31,89,31,224,31,54,31,193,31,170,31,29,31,107,31,107,30,153,31,180,31,220,31,53,31,30,31,48,31,48,30,48,29,226,31,61,31,18,31,168,31,230,31,128,31,104,31,138,31,245,31,199,31,226,31,12,31,12,30,12,29,12,28,174,31,174,30,17,31,17,30,17,29,200,31,200,30,108,31,117,31,117,30,50,31,19,31,61,31,33,31,64,31,30,31,30,30,76,31,209,31,209,30,13,31,102,31,79,31,184,31,163,31,128,31,86,31,86,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
