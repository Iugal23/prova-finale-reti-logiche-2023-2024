-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 321;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (164,0,62,0,226,0,210,0,149,0,184,0,50,0,0,0,20,0,254,0,104,0,119,0,22,0,0,0,205,0,143,0,82,0,81,0,151,0,0,0,225,0,66,0,70,0,150,0,166,0,9,0,64,0,0,0,27,0,148,0,129,0,201,0,44,0,84,0,6,0,0,0,150,0,245,0,62,0,196,0,122,0,171,0,99,0,140,0,174,0,0,0,136,0,80,0,236,0,41,0,214,0,242,0,198,0,202,0,202,0,139,0,0,0,0,0,250,0,0,0,0,0,74,0,186,0,0,0,0,0,234,0,49,0,0,0,165,0,95,0,194,0,0,0,56,0,148,0,120,0,0,0,109,0,166,0,180,0,222,0,145,0,34,0,249,0,141,0,0,0,169,0,211,0,164,0,82,0,0,0,208,0,57,0,176,0,216,0,202,0,98,0,118,0,164,0,130,0,0,0,188,0,138,0,197,0,75,0,0,0,0,0,37,0,0,0,0,0,0,0,112,0,239,0,0,0,239,0,248,0,81,0,178,0,49,0,106,0,142,0,69,0,82,0,109,0,139,0,34,0,0,0,136,0,253,0,0,0,202,0,213,0,169,0,124,0,62,0,171,0,0,0,254,0,0,0,166,0,141,0,91,0,0,0,59,0,101,0,179,0,58,0,218,0,0,0,136,0,1,0,2,0,0,0,212,0,69,0,111,0,186,0,175,0,6,0,39,0,0,0,0,0,22,0,0,0,127,0,0,0,216,0,0,0,36,0,198,0,0,0,190,0,0,0,24,0,0,0,0,0,151,0,212,0,197,0,188,0,0,0,0,0,0,0,248,0,222,0,78,0,147,0,93,0,153,0,198,0,0,0,183,0,187,0,187,0,21,0,78,0,182,0,0,0,0,0,111,0,54,0,76,0,0,0,114,0,146,0,159,0,10,0,0,0,21,0,191,0,215,0,172,0,0,0,0,0,57,0,119,0,31,0,108,0,38,0,147,0,186,0,90,0,0,0,34,0,16,0,221,0,200,0,0,0,69,0,190,0,147,0,0,0,0,0,234,0,121,0,0,0,121,0,105,0,170,0,57,0,140,0,242,0,191,0,2,0,232,0,88,0,184,0,0,0,35,0,111,0,4,0,186,0,0,0,193,0,208,0,93,0,102,0,132,0,159,0,32,0,212,0,121,0,36,0,250,0,9,0,158,0,222,0,4,0,124,0,104,0,63,0,201,0,141,0,0,0,0,0,233,0,15,0,151,0,77,0,0,0,178,0,0,0,57,0,143,0,164,0,0,0,0,0,184,0,211,0,245,0,241,0,0,0,169,0,25,0,96,0,171,0,122,0,37,0,13,0,26,0,159,0,144,0,77,0,46,0,29,0,44,0,255,0,193,0,0,0,31,0,0,0,18,0,0,0,158,0,216,0,152,0,197,0,87,0,53,0,195,0,0,0,0,0);
signal scenario_full  : scenario_type := (164,31,62,31,226,31,210,31,149,31,184,31,50,31,50,30,20,31,254,31,104,31,119,31,22,31,22,30,205,31,143,31,82,31,81,31,151,31,151,30,225,31,66,31,70,31,150,31,166,31,9,31,64,31,64,30,27,31,148,31,129,31,201,31,44,31,84,31,6,31,6,30,150,31,245,31,62,31,196,31,122,31,171,31,99,31,140,31,174,31,174,30,136,31,80,31,236,31,41,31,214,31,242,31,198,31,202,31,202,31,139,31,139,30,139,29,250,31,250,30,250,29,74,31,186,31,186,30,186,29,234,31,49,31,49,30,165,31,95,31,194,31,194,30,56,31,148,31,120,31,120,30,109,31,166,31,180,31,222,31,145,31,34,31,249,31,141,31,141,30,169,31,211,31,164,31,82,31,82,30,208,31,57,31,176,31,216,31,202,31,98,31,118,31,164,31,130,31,130,30,188,31,138,31,197,31,75,31,75,30,75,29,37,31,37,30,37,29,37,28,112,31,239,31,239,30,239,31,248,31,81,31,178,31,49,31,106,31,142,31,69,31,82,31,109,31,139,31,34,31,34,30,136,31,253,31,253,30,202,31,213,31,169,31,124,31,62,31,171,31,171,30,254,31,254,30,166,31,141,31,91,31,91,30,59,31,101,31,179,31,58,31,218,31,218,30,136,31,1,31,2,31,2,30,212,31,69,31,111,31,186,31,175,31,6,31,39,31,39,30,39,29,22,31,22,30,127,31,127,30,216,31,216,30,36,31,198,31,198,30,190,31,190,30,24,31,24,30,24,29,151,31,212,31,197,31,188,31,188,30,188,29,188,28,248,31,222,31,78,31,147,31,93,31,153,31,198,31,198,30,183,31,187,31,187,31,21,31,78,31,182,31,182,30,182,29,111,31,54,31,76,31,76,30,114,31,146,31,159,31,10,31,10,30,21,31,191,31,215,31,172,31,172,30,172,29,57,31,119,31,31,31,108,31,38,31,147,31,186,31,90,31,90,30,34,31,16,31,221,31,200,31,200,30,69,31,190,31,147,31,147,30,147,29,234,31,121,31,121,30,121,31,105,31,170,31,57,31,140,31,242,31,191,31,2,31,232,31,88,31,184,31,184,30,35,31,111,31,4,31,186,31,186,30,193,31,208,31,93,31,102,31,132,31,159,31,32,31,212,31,121,31,36,31,250,31,9,31,158,31,222,31,4,31,124,31,104,31,63,31,201,31,141,31,141,30,141,29,233,31,15,31,151,31,77,31,77,30,178,31,178,30,57,31,143,31,164,31,164,30,164,29,184,31,211,31,245,31,241,31,241,30,169,31,25,31,96,31,171,31,122,31,37,31,13,31,26,31,159,31,144,31,77,31,46,31,29,31,44,31,255,31,193,31,193,30,31,31,31,30,18,31,18,30,158,31,216,31,152,31,197,31,87,31,53,31,195,31,195,30,195,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
