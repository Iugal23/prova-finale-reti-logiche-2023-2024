-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 260;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (188,0,214,0,0,0,30,0,0,0,82,0,25,0,59,0,37,0,177,0,0,0,238,0,239,0,78,0,245,0,37,0,138,0,149,0,201,0,0,0,196,0,239,0,203,0,180,0,23,0,92,0,91,0,34,0,38,0,236,0,117,0,0,0,209,0,245,0,11,0,0,0,120,0,119,0,0,0,255,0,0,0,48,0,167,0,215,0,0,0,252,0,187,0,235,0,0,0,109,0,0,0,112,0,46,0,144,0,0,0,124,0,0,0,145,0,97,0,93,0,33,0,110,0,231,0,87,0,179,0,45,0,184,0,138,0,131,0,0,0,59,0,148,0,0,0,77,0,160,0,254,0,33,0,253,0,213,0,130,0,84,0,237,0,115,0,0,0,8,0,0,0,242,0,19,0,45,0,103,0,0,0,0,0,0,0,191,0,66,0,116,0,45,0,219,0,0,0,235,0,71,0,187,0,0,0,0,0,16,0,228,0,217,0,0,0,215,0,245,0,168,0,168,0,208,0,4,0,0,0,250,0,52,0,0,0,0,0,0,0,249,0,0,0,0,0,0,0,114,0,32,0,0,0,130,0,0,0,27,0,52,0,229,0,0,0,207,0,121,0,70,0,0,0,218,0,15,0,161,0,149,0,0,0,210,0,229,0,0,0,0,0,216,0,0,0,105,0,177,0,95,0,59,0,40,0,157,0,121,0,15,0,139,0,217,0,240,0,60,0,0,0,231,0,213,0,0,0,0,0,194,0,76,0,6,0,32,0,0,0,171,0,123,0,193,0,197,0,122,0,39,0,221,0,242,0,152,0,181,0,123,0,40,0,191,0,25,0,230,0,0,0,0,0,64,0,193,0,9,0,47,0,217,0,35,0,53,0,113,0,0,0,92,0,179,0,129,0,209,0,95,0,83,0,0,0,0,0,216,0,0,0,213,0,250,0,193,0,189,0,0,0,47,0,146,0,44,0,100,0,165,0,182,0,125,0,182,0,242,0,11,0,171,0,0,0,235,0,0,0,81,0,118,0,129,0,0,0,75,0,224,0,245,0,176,0,109,0,146,0,109,0,0,0,0,0,87,0,199,0,102,0,109,0,240,0,0,0,0,0,17,0,179,0,142,0,228,0,213,0,0,0,135,0,0,0,0,0,250,0,81,0,115,0,153,0,62,0,172,0);
signal scenario_full  : scenario_type := (188,31,214,31,214,30,30,31,30,30,82,31,25,31,59,31,37,31,177,31,177,30,238,31,239,31,78,31,245,31,37,31,138,31,149,31,201,31,201,30,196,31,239,31,203,31,180,31,23,31,92,31,91,31,34,31,38,31,236,31,117,31,117,30,209,31,245,31,11,31,11,30,120,31,119,31,119,30,255,31,255,30,48,31,167,31,215,31,215,30,252,31,187,31,235,31,235,30,109,31,109,30,112,31,46,31,144,31,144,30,124,31,124,30,145,31,97,31,93,31,33,31,110,31,231,31,87,31,179,31,45,31,184,31,138,31,131,31,131,30,59,31,148,31,148,30,77,31,160,31,254,31,33,31,253,31,213,31,130,31,84,31,237,31,115,31,115,30,8,31,8,30,242,31,19,31,45,31,103,31,103,30,103,29,103,28,191,31,66,31,116,31,45,31,219,31,219,30,235,31,71,31,187,31,187,30,187,29,16,31,228,31,217,31,217,30,215,31,245,31,168,31,168,31,208,31,4,31,4,30,250,31,52,31,52,30,52,29,52,28,249,31,249,30,249,29,249,28,114,31,32,31,32,30,130,31,130,30,27,31,52,31,229,31,229,30,207,31,121,31,70,31,70,30,218,31,15,31,161,31,149,31,149,30,210,31,229,31,229,30,229,29,216,31,216,30,105,31,177,31,95,31,59,31,40,31,157,31,121,31,15,31,139,31,217,31,240,31,60,31,60,30,231,31,213,31,213,30,213,29,194,31,76,31,6,31,32,31,32,30,171,31,123,31,193,31,197,31,122,31,39,31,221,31,242,31,152,31,181,31,123,31,40,31,191,31,25,31,230,31,230,30,230,29,64,31,193,31,9,31,47,31,217,31,35,31,53,31,113,31,113,30,92,31,179,31,129,31,209,31,95,31,83,31,83,30,83,29,216,31,216,30,213,31,250,31,193,31,189,31,189,30,47,31,146,31,44,31,100,31,165,31,182,31,125,31,182,31,242,31,11,31,171,31,171,30,235,31,235,30,81,31,118,31,129,31,129,30,75,31,224,31,245,31,176,31,109,31,146,31,109,31,109,30,109,29,87,31,199,31,102,31,109,31,240,31,240,30,240,29,17,31,179,31,142,31,228,31,213,31,213,30,135,31,135,30,135,29,250,31,81,31,115,31,153,31,62,31,172,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
