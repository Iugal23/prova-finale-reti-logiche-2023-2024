-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_859 is
end project_tb_859;

architecture project_tb_arch_859 of project_tb_859 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 513;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (189,0,19,0,226,0,160,0,172,0,0,0,225,0,0,0,0,0,198,0,129,0,108,0,56,0,0,0,119,0,254,0,230,0,0,0,197,0,250,0,175,0,144,0,157,0,121,0,85,0,245,0,240,0,154,0,170,0,74,0,117,0,79,0,105,0,80,0,80,0,221,0,196,0,189,0,72,0,70,0,103,0,47,0,122,0,94,0,163,0,163,0,20,0,248,0,227,0,62,0,161,0,232,0,254,0,0,0,0,0,93,0,16,0,14,0,92,0,166,0,2,0,0,0,202,0,18,0,240,0,0,0,73,0,0,0,0,0,250,0,0,0,0,0,0,0,199,0,95,0,153,0,251,0,209,0,68,0,29,0,0,0,87,0,77,0,194,0,254,0,250,0,251,0,223,0,53,0,119,0,122,0,230,0,239,0,3,0,44,0,182,0,53,0,148,0,231,0,118,0,70,0,0,0,141,0,112,0,48,0,74,0,19,0,229,0,128,0,20,0,93,0,130,0,103,0,199,0,221,0,10,0,163,0,230,0,216,0,175,0,82,0,0,0,240,0,241,0,0,0,0,0,77,0,102,0,4,0,0,0,0,0,55,0,180,0,68,0,0,0,82,0,144,0,52,0,14,0,68,0,138,0,204,0,230,0,99,0,18,0,16,0,22,0,0,0,124,0,214,0,205,0,0,0,67,0,83,0,111,0,209,0,197,0,225,0,46,0,197,0,185,0,0,0,124,0,0,0,0,0,200,0,176,0,118,0,220,0,0,0,251,0,156,0,75,0,0,0,106,0,69,0,73,0,126,0,196,0,213,0,0,0,10,0,164,0,204,0,170,0,236,0,158,0,142,0,240,0,0,0,30,0,246,0,19,0,244,0,0,0,115,0,60,0,0,0,0,0,22,0,222,0,0,0,112,0,124,0,37,0,63,0,91,0,0,0,188,0,95,0,89,0,223,0,13,0,0,0,150,0,189,0,150,0,134,0,9,0,252,0,155,0,157,0,73,0,0,0,176,0,154,0,204,0,48,0,28,0,10,0,145,0,57,0,0,0,186,0,0,0,111,0,115,0,147,0,34,0,115,0,162,0,246,0,154,0,54,0,129,0,0,0,0,0,206,0,213,0,206,0,159,0,145,0,68,0,64,0,14,0,135,0,59,0,0,0,195,0,149,0,59,0,144,0,88,0,0,0,153,0,221,0,189,0,0,0,183,0,36,0,130,0,240,0,8,0,88,0,174,0,0,0,0,0,78,0,132,0,208,0,238,0,215,0,251,0,223,0,96,0,0,0,177,0,222,0,181,0,211,0,234,0,129,0,33,0,0,0,230,0,0,0,23,0,0,0,181,0,218,0,93,0,214,0,105,0,0,0,210,0,147,0,0,0,123,0,74,0,172,0,0,0,64,0,72,0,0,0,36,0,0,0,214,0,31,0,107,0,138,0,0,0,9,0,59,0,250,0,150,0,58,0,0,0,172,0,0,0,77,0,151,0,0,0,0,0,206,0,122,0,106,0,0,0,25,0,73,0,52,0,0,0,23,0,0,0,0,0,176,0,13,0,105,0,232,0,0,0,2,0,106,0,253,0,0,0,0,0,0,0,251,0,139,0,204,0,0,0,141,0,239,0,0,0,0,0,222,0,54,0,88,0,197,0,113,0,134,0,221,0,216,0,59,0,183,0,91,0,78,0,0,0,162,0,0,0,1,0,51,0,214,0,70,0,183,0,4,0,247,0,0,0,0,0,0,0,5,0,245,0,107,0,0,0,86,0,15,0,0,0,0,0,240,0,82,0,62,0,0,0,89,0,120,0,124,0,22,0,0,0,251,0,0,0,0,0,165,0,255,0,30,0,118,0,109,0,0,0,115,0,182,0,150,0,129,0,110,0,11,0,0,0,220,0,0,0,111,0,202,0,0,0,83,0,159,0,236,0,237,0,59,0,0,0,96,0,194,0,107,0,0,0,155,0,24,0,53,0,97,0,127,0,7,0,160,0,100,0,243,0,0,0,174,0,77,0,36,0,216,0,30,0,98,0,198,0,0,0,3,0,0,0,242,0,17,0,0,0,48,0,255,0,161,0,238,0,129,0,84,0,109,0,0,0,146,0,0,0,152,0,43,0,168,0,69,0,7,0,0,0,97,0,0,0,147,0,224,0,41,0,21,0,0,0,94,0,0,0,127,0,78,0,0,0,123,0,239,0,11,0,103,0,148,0,103,0,114,0,48,0,18,0,0,0,10,0,155,0,64,0,0,0,216,0,84,0,145,0,219,0,175,0,168,0,238,0,0,0,0,0,0,0,0,0,0,0);
signal scenario_full  : scenario_type := (189,31,19,31,226,31,160,31,172,31,172,30,225,31,225,30,225,29,198,31,129,31,108,31,56,31,56,30,119,31,254,31,230,31,230,30,197,31,250,31,175,31,144,31,157,31,121,31,85,31,245,31,240,31,154,31,170,31,74,31,117,31,79,31,105,31,80,31,80,31,221,31,196,31,189,31,72,31,70,31,103,31,47,31,122,31,94,31,163,31,163,31,20,31,248,31,227,31,62,31,161,31,232,31,254,31,254,30,254,29,93,31,16,31,14,31,92,31,166,31,2,31,2,30,202,31,18,31,240,31,240,30,73,31,73,30,73,29,250,31,250,30,250,29,250,28,199,31,95,31,153,31,251,31,209,31,68,31,29,31,29,30,87,31,77,31,194,31,254,31,250,31,251,31,223,31,53,31,119,31,122,31,230,31,239,31,3,31,44,31,182,31,53,31,148,31,231,31,118,31,70,31,70,30,141,31,112,31,48,31,74,31,19,31,229,31,128,31,20,31,93,31,130,31,103,31,199,31,221,31,10,31,163,31,230,31,216,31,175,31,82,31,82,30,240,31,241,31,241,30,241,29,77,31,102,31,4,31,4,30,4,29,55,31,180,31,68,31,68,30,82,31,144,31,52,31,14,31,68,31,138,31,204,31,230,31,99,31,18,31,16,31,22,31,22,30,124,31,214,31,205,31,205,30,67,31,83,31,111,31,209,31,197,31,225,31,46,31,197,31,185,31,185,30,124,31,124,30,124,29,200,31,176,31,118,31,220,31,220,30,251,31,156,31,75,31,75,30,106,31,69,31,73,31,126,31,196,31,213,31,213,30,10,31,164,31,204,31,170,31,236,31,158,31,142,31,240,31,240,30,30,31,246,31,19,31,244,31,244,30,115,31,60,31,60,30,60,29,22,31,222,31,222,30,112,31,124,31,37,31,63,31,91,31,91,30,188,31,95,31,89,31,223,31,13,31,13,30,150,31,189,31,150,31,134,31,9,31,252,31,155,31,157,31,73,31,73,30,176,31,154,31,204,31,48,31,28,31,10,31,145,31,57,31,57,30,186,31,186,30,111,31,115,31,147,31,34,31,115,31,162,31,246,31,154,31,54,31,129,31,129,30,129,29,206,31,213,31,206,31,159,31,145,31,68,31,64,31,14,31,135,31,59,31,59,30,195,31,149,31,59,31,144,31,88,31,88,30,153,31,221,31,189,31,189,30,183,31,36,31,130,31,240,31,8,31,88,31,174,31,174,30,174,29,78,31,132,31,208,31,238,31,215,31,251,31,223,31,96,31,96,30,177,31,222,31,181,31,211,31,234,31,129,31,33,31,33,30,230,31,230,30,23,31,23,30,181,31,218,31,93,31,214,31,105,31,105,30,210,31,147,31,147,30,123,31,74,31,172,31,172,30,64,31,72,31,72,30,36,31,36,30,214,31,31,31,107,31,138,31,138,30,9,31,59,31,250,31,150,31,58,31,58,30,172,31,172,30,77,31,151,31,151,30,151,29,206,31,122,31,106,31,106,30,25,31,73,31,52,31,52,30,23,31,23,30,23,29,176,31,13,31,105,31,232,31,232,30,2,31,106,31,253,31,253,30,253,29,253,28,251,31,139,31,204,31,204,30,141,31,239,31,239,30,239,29,222,31,54,31,88,31,197,31,113,31,134,31,221,31,216,31,59,31,183,31,91,31,78,31,78,30,162,31,162,30,1,31,51,31,214,31,70,31,183,31,4,31,247,31,247,30,247,29,247,28,5,31,245,31,107,31,107,30,86,31,15,31,15,30,15,29,240,31,82,31,62,31,62,30,89,31,120,31,124,31,22,31,22,30,251,31,251,30,251,29,165,31,255,31,30,31,118,31,109,31,109,30,115,31,182,31,150,31,129,31,110,31,11,31,11,30,220,31,220,30,111,31,202,31,202,30,83,31,159,31,236,31,237,31,59,31,59,30,96,31,194,31,107,31,107,30,155,31,24,31,53,31,97,31,127,31,7,31,160,31,100,31,243,31,243,30,174,31,77,31,36,31,216,31,30,31,98,31,198,31,198,30,3,31,3,30,242,31,17,31,17,30,48,31,255,31,161,31,238,31,129,31,84,31,109,31,109,30,146,31,146,30,152,31,43,31,168,31,69,31,7,31,7,30,97,31,97,30,147,31,224,31,41,31,21,31,21,30,94,31,94,30,127,31,78,31,78,30,123,31,239,31,11,31,103,31,148,31,103,31,114,31,48,31,18,31,18,30,10,31,155,31,64,31,64,30,216,31,84,31,145,31,219,31,175,31,168,31,238,31,238,30,238,29,238,28,238,27,238,26);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
