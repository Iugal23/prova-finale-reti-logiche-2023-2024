-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 263;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,0,0,58,0,216,0,0,0,168,0,192,0,0,0,50,0,94,0,23,0,19,0,58,0,75,0,0,0,2,0,0,0,0,0,201,0,115,0,133,0,163,0,219,0,131,0,0,0,242,0,10,0,78,0,49,0,127,0,0,0,0,0,0,0,0,0,80,0,169,0,107,0,211,0,65,0,99,0,249,0,56,0,62,0,0,0,0,0,0,0,233,0,226,0,99,0,141,0,206,0,0,0,44,0,0,0,159,0,168,0,115,0,99,0,43,0,0,0,211,0,244,0,48,0,134,0,170,0,62,0,120,0,245,0,137,0,89,0,10,0,235,0,110,0,243,0,236,0,67,0,232,0,6,0,23,0,153,0,170,0,0,0,213,0,151,0,41,0,238,0,0,0,34,0,0,0,0,0,0,0,150,0,18,0,80,0,19,0,0,0,0,0,53,0,185,0,209,0,0,0,103,0,218,0,32,0,192,0,172,0,22,0,49,0,0,0,103,0,0,0,57,0,9,0,60,0,0,0,168,0,191,0,24,0,0,0,94,0,251,0,126,0,41,0,47,0,0,0,235,0,122,0,86,0,226,0,160,0,0,0,3,0,153,0,174,0,144,0,136,0,0,0,52,0,78,0,0,0,176,0,0,0,0,0,248,0,145,0,129,0,0,0,0,0,181,0,57,0,5,0,44,0,176,0,0,0,3,0,0,0,142,0,0,0,68,0,140,0,0,0,0,0,132,0,0,0,223,0,149,0,246,0,116,0,75,0,234,0,0,0,8,0,46,0,181,0,151,0,110,0,183,0,109,0,0,0,79,0,231,0,138,0,160,0,0,0,50,0,74,0,148,0,200,0,19,0,222,0,140,0,241,0,180,0,252,0,189,0,166,0,140,0,216,0,234,0,112,0,9,0,132,0,0,0,149,0,230,0,104,0,0,0,0,0,0,0,243,0,105,0,58,0,107,0,155,0,84,0,99,0,0,0,241,0,233,0,50,0,97,0,184,0,203,0,2,0,0,0,0,0,246,0,61,0,241,0,22,0,0,0,144,0,35,0,67,0,185,0,52,0,121,0,0,0,143,0,215,0,85,0,218,0,0,0,114,0,69,0,0,0,0,0,132,0,0,0,80,0,100,0,38,0,198,0,167,0,212,0,250,0,0,0,252,0,50,0,45,0,126,0,246,0);
signal scenario_full  : scenario_type := (0,0,0,0,0,0,58,31,216,31,216,30,168,31,192,31,192,30,50,31,94,31,23,31,19,31,58,31,75,31,75,30,2,31,2,30,2,29,201,31,115,31,133,31,163,31,219,31,131,31,131,30,242,31,10,31,78,31,49,31,127,31,127,30,127,29,127,28,127,27,80,31,169,31,107,31,211,31,65,31,99,31,249,31,56,31,62,31,62,30,62,29,62,28,233,31,226,31,99,31,141,31,206,31,206,30,44,31,44,30,159,31,168,31,115,31,99,31,43,31,43,30,211,31,244,31,48,31,134,31,170,31,62,31,120,31,245,31,137,31,89,31,10,31,235,31,110,31,243,31,236,31,67,31,232,31,6,31,23,31,153,31,170,31,170,30,213,31,151,31,41,31,238,31,238,30,34,31,34,30,34,29,34,28,150,31,18,31,80,31,19,31,19,30,19,29,53,31,185,31,209,31,209,30,103,31,218,31,32,31,192,31,172,31,22,31,49,31,49,30,103,31,103,30,57,31,9,31,60,31,60,30,168,31,191,31,24,31,24,30,94,31,251,31,126,31,41,31,47,31,47,30,235,31,122,31,86,31,226,31,160,31,160,30,3,31,153,31,174,31,144,31,136,31,136,30,52,31,78,31,78,30,176,31,176,30,176,29,248,31,145,31,129,31,129,30,129,29,181,31,57,31,5,31,44,31,176,31,176,30,3,31,3,30,142,31,142,30,68,31,140,31,140,30,140,29,132,31,132,30,223,31,149,31,246,31,116,31,75,31,234,31,234,30,8,31,46,31,181,31,151,31,110,31,183,31,109,31,109,30,79,31,231,31,138,31,160,31,160,30,50,31,74,31,148,31,200,31,19,31,222,31,140,31,241,31,180,31,252,31,189,31,166,31,140,31,216,31,234,31,112,31,9,31,132,31,132,30,149,31,230,31,104,31,104,30,104,29,104,28,243,31,105,31,58,31,107,31,155,31,84,31,99,31,99,30,241,31,233,31,50,31,97,31,184,31,203,31,2,31,2,30,2,29,246,31,61,31,241,31,22,31,22,30,144,31,35,31,67,31,185,31,52,31,121,31,121,30,143,31,215,31,85,31,218,31,218,30,114,31,69,31,69,30,69,29,132,31,132,30,80,31,100,31,38,31,198,31,167,31,212,31,250,31,250,30,252,31,50,31,45,31,126,31,246,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
