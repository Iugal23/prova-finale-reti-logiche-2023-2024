-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 733;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (246,0,153,0,246,0,89,0,206,0,136,0,0,0,0,0,126,0,87,0,150,0,203,0,109,0,0,0,0,0,243,0,36,0,184,0,0,0,0,0,104,0,0,0,0,0,194,0,11,0,61,0,167,0,143,0,137,0,0,0,0,0,0,0,107,0,114,0,125,0,162,0,0,0,104,0,124,0,0,0,0,0,206,0,42,0,171,0,183,0,44,0,119,0,46,0,0,0,86,0,58,0,223,0,67,0,70,0,99,0,124,0,164,0,127,0,232,0,240,0,114,0,0,0,93,0,161,0,24,0,201,0,141,0,42,0,162,0,223,0,107,0,93,0,0,0,181,0,0,0,0,0,0,0,203,0,80,0,11,0,254,0,0,0,112,0,114,0,220,0,223,0,0,0,0,0,0,0,3,0,189,0,249,0,60,0,202,0,232,0,119,0,52,0,0,0,76,0,101,0,153,0,196,0,24,0,180,0,120,0,5,0,111,0,221,0,0,0,0,0,198,0,98,0,248,0,118,0,202,0,124,0,0,0,52,0,86,0,162,0,52,0,75,0,108,0,158,0,224,0,125,0,234,0,35,0,0,0,34,0,0,0,83,0,99,0,80,0,0,0,192,0,69,0,4,0,132,0,34,0,128,0,36,0,23,0,221,0,8,0,63,0,230,0,54,0,23,0,134,0,105,0,194,0,128,0,52,0,135,0,32,0,228,0,211,0,31,0,128,0,146,0,61,0,0,0,163,0,200,0,32,0,102,0,0,0,82,0,185,0,41,0,0,0,0,0,0,0,55,0,1,0,192,0,24,0,0,0,158,0,85,0,0,0,0,0,189,0,49,0,189,0,17,0,244,0,104,0,0,0,99,0,101,0,163,0,0,0,31,0,194,0,99,0,0,0,140,0,107,0,198,0,75,0,58,0,229,0,36,0,176,0,124,0,0,0,229,0,0,0,0,0,0,0,41,0,147,0,0,0,184,0,62,0,114,0,93,0,223,0,125,0,0,0,180,0,234,0,74,0,219,0,251,0,0,0,0,0,42,0,58,0,62,0,242,0,165,0,0,0,222,0,0,0,30,0,28,0,0,0,0,0,70,0,123,0,0,0,0,0,170,0,0,0,157,0,71,0,91,0,166,0,130,0,107,0,42,0,190,0,212,0,0,0,114,0,2,0,194,0,223,0,162,0,0,0,95,0,45,0,249,0,0,0,121,0,49,0,154,0,191,0,73,0,16,0,65,0,249,0,7,0,215,0,187,0,162,0,194,0,205,0,38,0,0,0,0,0,225,0,90,0,115,0,0,0,0,0,195,0,73,0,85,0,0,0,35,0,107,0,0,0,162,0,76,0,116,0,238,0,42,0,0,0,126,0,129,0,0,0,120,0,129,0,154,0,86,0,0,0,157,0,0,0,141,0,112,0,191,0,160,0,0,0,204,0,252,0,215,0,136,0,56,0,0,0,85,0,74,0,43,0,141,0,22,0,0,0,67,0,177,0,21,0,0,0,229,0,0,0,244,0,94,0,61,0,221,0,123,0,110,0,58,0,0,0,216,0,0,0,174,0,151,0,125,0,0,0,0,0,230,0,208,0,107,0,0,0,44,0,0,0,197,0,0,0,106,0,240,0,0,0,52,0,195,0,37,0,45,0,16,0,89,0,0,0,144,0,183,0,64,0,147,0,138,0,30,0,193,0,141,0,113,0,60,0,246,0,234,0,0,0,0,0,134,0,206,0,214,0,0,0,0,0,194,0,0,0,149,0,0,0,246,0,0,0,36,0,78,0,87,0,0,0,0,0,77,0,37,0,151,0,65,0,180,0,177,0,80,0,45,0,204,0,251,0,228,0,140,0,42,0,252,0,0,0,96,0,26,0,164,0,210,0,216,0,0,0,125,0,119,0,194,0,0,0,109,0,107,0,0,0,0,0,0,0,77,0,56,0,117,0,163,0,139,0,80,0,46,0,0,0,217,0,120,0,0,0,244,0,210,0,10,0,0,0,27,0,0,0,38,0,242,0,245,0,57,0,80,0,20,0,167,0,0,0,197,0,191,0,188,0,229,0,99,0,27,0,248,0,39,0,86,0,131,0,220,0,0,0,239,0,0,0,250,0,133,0,130,0,96,0,79,0,103,0,94,0,157,0,0,0,94,0,33,0,0,0,223,0,164,0,162,0,94,0,230,0,242,0,121,0,195,0,34,0,0,0,235,0,255,0,147,0,159,0,227,0,149,0,246,0,135,0,132,0,64,0,153,0,100,0,60,0,130,0,4,0,152,0,116,0,38,0,191,0,248,0,104,0,125,0,111,0,248,0,0,0,65,0,49,0,200,0,43,0,34,0,124,0,154,0,12,0,79,0,234,0,172,0,40,0,46,0,171,0,123,0,82,0,19,0,169,0,0,0,0,0,197,0,106,0,150,0,213,0,121,0,31,0,122,0,24,0,176,0,92,0,237,0,184,0,18,0,212,0,0,0,109,0,249,0,51,0,0,0,47,0,216,0,0,0,126,0,0,0,59,0,177,0,240,0,136,0,53,0,135,0,244,0,0,0,136,0,0,0,67,0,142,0,0,0,140,0,46,0,0,0,120,0,25,0,0,0,19,0,0,0,221,0,162,0,99,0,240,0,79,0,244,0,142,0,207,0,0,0,128,0,0,0,190,0,0,0,0,0,140,0,79,0,70,0,145,0,220,0,182,0,29,0,129,0,231,0,156,0,0,0,164,0,0,0,235,0,26,0,0,0,132,0,78,0,0,0,0,0,0,0,173,0,32,0,26,0,0,0,152,0,81,0,97,0,35,0,31,0,208,0,184,0,139,0,48,0,86,0,34,0,0,0,197,0,174,0,141,0,0,0,0,0,1,0,3,0,70,0,0,0,116,0,62,0,134,0,52,0,185,0,44,0,96,0,116,0,0,0,96,0,0,0,191,0,109,0,23,0,218,0,149,0,135,0,155,0,135,0,0,0,153,0,0,0,0,0,161,0,112,0,219,0,0,0,5,0,0,0,100,0,6,0,47,0,6,0,220,0,172,0,41,0,176,0,93,0,0,0,180,0,10,0,0,0,123,0,0,0,0,0,39,0,128,0,78,0,86,0,0,0,162,0,145,0,231,0,0,0,27,0,121,0,137,0,0,0,11,0,144,0,9,0,2,0,5,0,252,0,6,0,65,0,76,0,0,0,0,0,246,0,110,0,73,0,221,0,231,0,234,0,182,0,180,0,0,0,218,0,0,0,220,0,86,0,149,0,97,0,74,0,40,0,31,0,180,0,198,0,0,0,124,0,244,0,242,0,42,0);
signal scenario_full  : scenario_type := (246,31,153,31,246,31,89,31,206,31,136,31,136,30,136,29,126,31,87,31,150,31,203,31,109,31,109,30,109,29,243,31,36,31,184,31,184,30,184,29,104,31,104,30,104,29,194,31,11,31,61,31,167,31,143,31,137,31,137,30,137,29,137,28,107,31,114,31,125,31,162,31,162,30,104,31,124,31,124,30,124,29,206,31,42,31,171,31,183,31,44,31,119,31,46,31,46,30,86,31,58,31,223,31,67,31,70,31,99,31,124,31,164,31,127,31,232,31,240,31,114,31,114,30,93,31,161,31,24,31,201,31,141,31,42,31,162,31,223,31,107,31,93,31,93,30,181,31,181,30,181,29,181,28,203,31,80,31,11,31,254,31,254,30,112,31,114,31,220,31,223,31,223,30,223,29,223,28,3,31,189,31,249,31,60,31,202,31,232,31,119,31,52,31,52,30,76,31,101,31,153,31,196,31,24,31,180,31,120,31,5,31,111,31,221,31,221,30,221,29,198,31,98,31,248,31,118,31,202,31,124,31,124,30,52,31,86,31,162,31,52,31,75,31,108,31,158,31,224,31,125,31,234,31,35,31,35,30,34,31,34,30,83,31,99,31,80,31,80,30,192,31,69,31,4,31,132,31,34,31,128,31,36,31,23,31,221,31,8,31,63,31,230,31,54,31,23,31,134,31,105,31,194,31,128,31,52,31,135,31,32,31,228,31,211,31,31,31,128,31,146,31,61,31,61,30,163,31,200,31,32,31,102,31,102,30,82,31,185,31,41,31,41,30,41,29,41,28,55,31,1,31,192,31,24,31,24,30,158,31,85,31,85,30,85,29,189,31,49,31,189,31,17,31,244,31,104,31,104,30,99,31,101,31,163,31,163,30,31,31,194,31,99,31,99,30,140,31,107,31,198,31,75,31,58,31,229,31,36,31,176,31,124,31,124,30,229,31,229,30,229,29,229,28,41,31,147,31,147,30,184,31,62,31,114,31,93,31,223,31,125,31,125,30,180,31,234,31,74,31,219,31,251,31,251,30,251,29,42,31,58,31,62,31,242,31,165,31,165,30,222,31,222,30,30,31,28,31,28,30,28,29,70,31,123,31,123,30,123,29,170,31,170,30,157,31,71,31,91,31,166,31,130,31,107,31,42,31,190,31,212,31,212,30,114,31,2,31,194,31,223,31,162,31,162,30,95,31,45,31,249,31,249,30,121,31,49,31,154,31,191,31,73,31,16,31,65,31,249,31,7,31,215,31,187,31,162,31,194,31,205,31,38,31,38,30,38,29,225,31,90,31,115,31,115,30,115,29,195,31,73,31,85,31,85,30,35,31,107,31,107,30,162,31,76,31,116,31,238,31,42,31,42,30,126,31,129,31,129,30,120,31,129,31,154,31,86,31,86,30,157,31,157,30,141,31,112,31,191,31,160,31,160,30,204,31,252,31,215,31,136,31,56,31,56,30,85,31,74,31,43,31,141,31,22,31,22,30,67,31,177,31,21,31,21,30,229,31,229,30,244,31,94,31,61,31,221,31,123,31,110,31,58,31,58,30,216,31,216,30,174,31,151,31,125,31,125,30,125,29,230,31,208,31,107,31,107,30,44,31,44,30,197,31,197,30,106,31,240,31,240,30,52,31,195,31,37,31,45,31,16,31,89,31,89,30,144,31,183,31,64,31,147,31,138,31,30,31,193,31,141,31,113,31,60,31,246,31,234,31,234,30,234,29,134,31,206,31,214,31,214,30,214,29,194,31,194,30,149,31,149,30,246,31,246,30,36,31,78,31,87,31,87,30,87,29,77,31,37,31,151,31,65,31,180,31,177,31,80,31,45,31,204,31,251,31,228,31,140,31,42,31,252,31,252,30,96,31,26,31,164,31,210,31,216,31,216,30,125,31,119,31,194,31,194,30,109,31,107,31,107,30,107,29,107,28,77,31,56,31,117,31,163,31,139,31,80,31,46,31,46,30,217,31,120,31,120,30,244,31,210,31,10,31,10,30,27,31,27,30,38,31,242,31,245,31,57,31,80,31,20,31,167,31,167,30,197,31,191,31,188,31,229,31,99,31,27,31,248,31,39,31,86,31,131,31,220,31,220,30,239,31,239,30,250,31,133,31,130,31,96,31,79,31,103,31,94,31,157,31,157,30,94,31,33,31,33,30,223,31,164,31,162,31,94,31,230,31,242,31,121,31,195,31,34,31,34,30,235,31,255,31,147,31,159,31,227,31,149,31,246,31,135,31,132,31,64,31,153,31,100,31,60,31,130,31,4,31,152,31,116,31,38,31,191,31,248,31,104,31,125,31,111,31,248,31,248,30,65,31,49,31,200,31,43,31,34,31,124,31,154,31,12,31,79,31,234,31,172,31,40,31,46,31,171,31,123,31,82,31,19,31,169,31,169,30,169,29,197,31,106,31,150,31,213,31,121,31,31,31,122,31,24,31,176,31,92,31,237,31,184,31,18,31,212,31,212,30,109,31,249,31,51,31,51,30,47,31,216,31,216,30,126,31,126,30,59,31,177,31,240,31,136,31,53,31,135,31,244,31,244,30,136,31,136,30,67,31,142,31,142,30,140,31,46,31,46,30,120,31,25,31,25,30,19,31,19,30,221,31,162,31,99,31,240,31,79,31,244,31,142,31,207,31,207,30,128,31,128,30,190,31,190,30,190,29,140,31,79,31,70,31,145,31,220,31,182,31,29,31,129,31,231,31,156,31,156,30,164,31,164,30,235,31,26,31,26,30,132,31,78,31,78,30,78,29,78,28,173,31,32,31,26,31,26,30,152,31,81,31,97,31,35,31,31,31,208,31,184,31,139,31,48,31,86,31,34,31,34,30,197,31,174,31,141,31,141,30,141,29,1,31,3,31,70,31,70,30,116,31,62,31,134,31,52,31,185,31,44,31,96,31,116,31,116,30,96,31,96,30,191,31,109,31,23,31,218,31,149,31,135,31,155,31,135,31,135,30,153,31,153,30,153,29,161,31,112,31,219,31,219,30,5,31,5,30,100,31,6,31,47,31,6,31,220,31,172,31,41,31,176,31,93,31,93,30,180,31,10,31,10,30,123,31,123,30,123,29,39,31,128,31,78,31,86,31,86,30,162,31,145,31,231,31,231,30,27,31,121,31,137,31,137,30,11,31,144,31,9,31,2,31,5,31,252,31,6,31,65,31,76,31,76,30,76,29,246,31,110,31,73,31,221,31,231,31,234,31,182,31,180,31,180,30,218,31,218,30,220,31,86,31,149,31,97,31,74,31,40,31,31,31,180,31,198,31,198,30,124,31,244,31,242,31,42,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
