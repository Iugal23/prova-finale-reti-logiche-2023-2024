-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 798;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (197,0,148,0,241,0,31,0,148,0,226,0,90,0,0,0,174,0,0,0,208,0,114,0,218,0,44,0,176,0,93,0,230,0,127,0,0,0,0,0,21,0,0,0,200,0,27,0,215,0,146,0,162,0,124,0,194,0,0,0,158,0,201,0,49,0,191,0,214,0,0,0,116,0,0,0,31,0,69,0,251,0,36,0,154,0,193,0,147,0,108,0,47,0,120,0,141,0,122,0,0,0,104,0,44,0,64,0,200,0,10,0,200,0,56,0,0,0,0,0,221,0,0,0,0,0,214,0,226,0,0,0,89,0,39,0,34,0,218,0,0,0,213,0,222,0,0,0,157,0,105,0,189,0,208,0,117,0,86,0,211,0,162,0,0,0,0,0,187,0,228,0,81,0,249,0,0,0,234,0,0,0,0,0,181,0,179,0,70,0,85,0,11,0,111,0,23,0,197,0,201,0,161,0,38,0,0,0,168,0,0,0,52,0,0,0,47,0,236,0,27,0,0,0,209,0,235,0,187,0,71,0,0,0,151,0,104,0,101,0,160,0,0,0,22,0,41,0,3,0,250,0,24,0,147,0,203,0,183,0,186,0,0,0,0,0,251,0,125,0,253,0,11,0,28,0,136,0,212,0,172,0,126,0,0,0,216,0,187,0,204,0,0,0,29,0,90,0,205,0,36,0,0,0,30,0,65,0,177,0,193,0,64,0,232,0,234,0,58,0,188,0,0,0,132,0,104,0,166,0,92,0,175,0,0,0,0,0,131,0,101,0,0,0,0,0,84,0,232,0,142,0,41,0,0,0,10,0,218,0,48,0,0,0,76,0,76,0,120,0,0,0,122,0,98,0,0,0,145,0,101,0,198,0,156,0,76,0,21,0,244,0,0,0,0,0,229,0,251,0,44,0,29,0,249,0,127,0,179,0,0,0,82,0,70,0,216,0,60,0,243,0,90,0,183,0,219,0,219,0,66,0,190,0,178,0,0,0,134,0,185,0,243,0,12,0,129,0,207,0,105,0,184,0,118,0,0,0,93,0,232,0,59,0,23,0,12,0,114,0,189,0,63,0,88,0,153,0,16,0,0,0,87,0,17,0,203,0,178,0,0,0,187,0,213,0,207,0,3,0,233,0,130,0,105,0,7,0,58,0,46,0,221,0,131,0,136,0,121,0,0,0,0,0,104,0,86,0,57,0,0,0,0,0,227,0,156,0,0,0,0,0,67,0,2,0,151,0,174,0,0,0,79,0,141,0,175,0,12,0,235,0,122,0,49,0,212,0,0,0,128,0,199,0,0,0,96,0,251,0,78,0,222,0,33,0,244,0,152,0,157,0,199,0,107,0,0,0,173,0,0,0,78,0,84,0,0,0,48,0,0,0,171,0,0,0,246,0,178,0,213,0,182,0,221,0,235,0,200,0,50,0,128,0,0,0,208,0,180,0,61,0,0,0,239,0,124,0,0,0,157,0,12,0,250,0,42,0,146,0,163,0,19,0,0,0,75,0,0,0,120,0,162,0,128,0,106,0,0,0,0,0,56,0,220,0,250,0,13,0,79,0,0,0,114,0,0,0,166,0,86,0,72,0,133,0,130,0,208,0,214,0,203,0,15,0,155,0,218,0,0,0,74,0,0,0,155,0,175,0,239,0,147,0,126,0,0,0,0,0,0,0,83,0,128,0,0,0,136,0,178,0,249,0,186,0,93,0,108,0,7,0,111,0,31,0,179,0,154,0,15,0,199,0,34,0,0,0,0,0,42,0,190,0,243,0,248,0,132,0,2,0,204,0,105,0,0,0,191,0,102,0,48,0,227,0,34,0,0,0,106,0,183,0,0,0,166,0,7,0,0,0,0,0,50,0,90,0,171,0,0,0,255,0,209,0,65,0,11,0,0,0,80,0,36,0,87,0,177,0,0,0,108,0,233,0,174,0,0,0,99,0,5,0,236,0,14,0,95,0,121,0,0,0,104,0,144,0,234,0,0,0,129,0,0,0,76,0,235,0,89,0,247,0,0,0,0,0,76,0,17,0,0,0,192,0,0,0,251,0,252,0,0,0,0,0,0,0,109,0,185,0,0,0,148,0,15,0,0,0,106,0,0,0,0,0,0,0,115,0,41,0,58,0,85,0,221,0,141,0,159,0,237,0,33,0,204,0,0,0,68,0,0,0,148,0,132,0,1,0,102,0,0,0,105,0,0,0,70,0,67,0,0,0,18,0,233,0,218,0,0,0,0,0,0,0,70,0,51,0,39,0,158,0,16,0,30,0,0,0,139,0,0,0,63,0,4,0,0,0,156,0,171,0,92,0,0,0,136,0,85,0,5,0,57,0,184,0,197,0,42,0,0,0,223,0,222,0,0,0,0,0,0,0,122,0,136,0,0,0,140,0,0,0,147,0,13,0,24,0,61,0,118,0,159,0,0,0,0,0,41,0,49,0,0,0,77,0,169,0,86,0,183,0,101,0,195,0,240,0,171,0,128,0,200,0,0,0,233,0,133,0,136,0,242,0,14,0,97,0,223,0,153,0,186,0,4,0,0,0,80,0,15,0,219,0,0,0,169,0,0,0,17,0,108,0,13,0,220,0,115,0,142,0,68,0,27,0,77,0,0,0,151,0,155,0,250,0,94,0,44,0,0,0,38,0,253,0,95,0,1,0,121,0,229,0,0,0,153,0,115,0,211,0,191,0,194,0,0,0,94,0,85,0,0,0,29,0,56,0,0,0,220,0,206,0,219,0,212,0,213,0,50,0,72,0,0,0,177,0,153,0,237,0,118,0,224,0,207,0,248,0,84,0,249,0,128,0,218,0,225,0,106,0,106,0,0,0,105,0,0,0,204,0,83,0,78,0,207,0,0,0,50,0,110,0,225,0,17,0,0,0,190,0,17,0,0,0,42,0,55,0,247,0,190,0,235,0,249,0,0,0,241,0,146,0,189,0,135,0,121,0,128,0,43,0,102,0,246,0,42,0,146,0,0,0,136,0,33,0,201,0,10,0,101,0,77,0,18,0,30,0,232,0,0,0,22,0,27,0,145,0,150,0,16,0,210,0,237,0,163,0,242,0,136,0,0,0,0,0,120,0,141,0,19,0,122,0,25,0,217,0,0,0,142,0,8,0,13,0,15,0,0,0,204,0,140,0,136,0,72,0,0,0,0,0,0,0,178,0,131,0,203,0,111,0,171,0,115,0,78,0,0,0,0,0,7,0,28,0,84,0,0,0,0,0,133,0,39,0,226,0,0,0,156,0,127,0,67,0,114,0,190,0,27,0,17,0,242,0,239,0,254,0,127,0,0,0,154,0,190,0,176,0,204,0,42,0,119,0,0,0,135,0,17,0,0,0,66,0,252,0,213,0,81,0,95,0,194,0,149,0,0,0,102,0,134,0,127,0,73,0,0,0,242,0,11,0,143,0,155,0,75,0,156,0,74,0,203,0,159,0,94,0,0,0,187,0,0,0,72,0,35,0,55,0,0,0,5,0,23,0,128,0,123,0,42,0,13,0,59,0,52,0,165,0,162,0,160,0,125,0,27,0,0,0,135,0,96,0,0,0,51,0,2,0,90,0,0,0,172,0,84,0,63,0);
signal scenario_full  : scenario_type := (197,31,148,31,241,31,31,31,148,31,226,31,90,31,90,30,174,31,174,30,208,31,114,31,218,31,44,31,176,31,93,31,230,31,127,31,127,30,127,29,21,31,21,30,200,31,27,31,215,31,146,31,162,31,124,31,194,31,194,30,158,31,201,31,49,31,191,31,214,31,214,30,116,31,116,30,31,31,69,31,251,31,36,31,154,31,193,31,147,31,108,31,47,31,120,31,141,31,122,31,122,30,104,31,44,31,64,31,200,31,10,31,200,31,56,31,56,30,56,29,221,31,221,30,221,29,214,31,226,31,226,30,89,31,39,31,34,31,218,31,218,30,213,31,222,31,222,30,157,31,105,31,189,31,208,31,117,31,86,31,211,31,162,31,162,30,162,29,187,31,228,31,81,31,249,31,249,30,234,31,234,30,234,29,181,31,179,31,70,31,85,31,11,31,111,31,23,31,197,31,201,31,161,31,38,31,38,30,168,31,168,30,52,31,52,30,47,31,236,31,27,31,27,30,209,31,235,31,187,31,71,31,71,30,151,31,104,31,101,31,160,31,160,30,22,31,41,31,3,31,250,31,24,31,147,31,203,31,183,31,186,31,186,30,186,29,251,31,125,31,253,31,11,31,28,31,136,31,212,31,172,31,126,31,126,30,216,31,187,31,204,31,204,30,29,31,90,31,205,31,36,31,36,30,30,31,65,31,177,31,193,31,64,31,232,31,234,31,58,31,188,31,188,30,132,31,104,31,166,31,92,31,175,31,175,30,175,29,131,31,101,31,101,30,101,29,84,31,232,31,142,31,41,31,41,30,10,31,218,31,48,31,48,30,76,31,76,31,120,31,120,30,122,31,98,31,98,30,145,31,101,31,198,31,156,31,76,31,21,31,244,31,244,30,244,29,229,31,251,31,44,31,29,31,249,31,127,31,179,31,179,30,82,31,70,31,216,31,60,31,243,31,90,31,183,31,219,31,219,31,66,31,190,31,178,31,178,30,134,31,185,31,243,31,12,31,129,31,207,31,105,31,184,31,118,31,118,30,93,31,232,31,59,31,23,31,12,31,114,31,189,31,63,31,88,31,153,31,16,31,16,30,87,31,17,31,203,31,178,31,178,30,187,31,213,31,207,31,3,31,233,31,130,31,105,31,7,31,58,31,46,31,221,31,131,31,136,31,121,31,121,30,121,29,104,31,86,31,57,31,57,30,57,29,227,31,156,31,156,30,156,29,67,31,2,31,151,31,174,31,174,30,79,31,141,31,175,31,12,31,235,31,122,31,49,31,212,31,212,30,128,31,199,31,199,30,96,31,251,31,78,31,222,31,33,31,244,31,152,31,157,31,199,31,107,31,107,30,173,31,173,30,78,31,84,31,84,30,48,31,48,30,171,31,171,30,246,31,178,31,213,31,182,31,221,31,235,31,200,31,50,31,128,31,128,30,208,31,180,31,61,31,61,30,239,31,124,31,124,30,157,31,12,31,250,31,42,31,146,31,163,31,19,31,19,30,75,31,75,30,120,31,162,31,128,31,106,31,106,30,106,29,56,31,220,31,250,31,13,31,79,31,79,30,114,31,114,30,166,31,86,31,72,31,133,31,130,31,208,31,214,31,203,31,15,31,155,31,218,31,218,30,74,31,74,30,155,31,175,31,239,31,147,31,126,31,126,30,126,29,126,28,83,31,128,31,128,30,136,31,178,31,249,31,186,31,93,31,108,31,7,31,111,31,31,31,179,31,154,31,15,31,199,31,34,31,34,30,34,29,42,31,190,31,243,31,248,31,132,31,2,31,204,31,105,31,105,30,191,31,102,31,48,31,227,31,34,31,34,30,106,31,183,31,183,30,166,31,7,31,7,30,7,29,50,31,90,31,171,31,171,30,255,31,209,31,65,31,11,31,11,30,80,31,36,31,87,31,177,31,177,30,108,31,233,31,174,31,174,30,99,31,5,31,236,31,14,31,95,31,121,31,121,30,104,31,144,31,234,31,234,30,129,31,129,30,76,31,235,31,89,31,247,31,247,30,247,29,76,31,17,31,17,30,192,31,192,30,251,31,252,31,252,30,252,29,252,28,109,31,185,31,185,30,148,31,15,31,15,30,106,31,106,30,106,29,106,28,115,31,41,31,58,31,85,31,221,31,141,31,159,31,237,31,33,31,204,31,204,30,68,31,68,30,148,31,132,31,1,31,102,31,102,30,105,31,105,30,70,31,67,31,67,30,18,31,233,31,218,31,218,30,218,29,218,28,70,31,51,31,39,31,158,31,16,31,30,31,30,30,139,31,139,30,63,31,4,31,4,30,156,31,171,31,92,31,92,30,136,31,85,31,5,31,57,31,184,31,197,31,42,31,42,30,223,31,222,31,222,30,222,29,222,28,122,31,136,31,136,30,140,31,140,30,147,31,13,31,24,31,61,31,118,31,159,31,159,30,159,29,41,31,49,31,49,30,77,31,169,31,86,31,183,31,101,31,195,31,240,31,171,31,128,31,200,31,200,30,233,31,133,31,136,31,242,31,14,31,97,31,223,31,153,31,186,31,4,31,4,30,80,31,15,31,219,31,219,30,169,31,169,30,17,31,108,31,13,31,220,31,115,31,142,31,68,31,27,31,77,31,77,30,151,31,155,31,250,31,94,31,44,31,44,30,38,31,253,31,95,31,1,31,121,31,229,31,229,30,153,31,115,31,211,31,191,31,194,31,194,30,94,31,85,31,85,30,29,31,56,31,56,30,220,31,206,31,219,31,212,31,213,31,50,31,72,31,72,30,177,31,153,31,237,31,118,31,224,31,207,31,248,31,84,31,249,31,128,31,218,31,225,31,106,31,106,31,106,30,105,31,105,30,204,31,83,31,78,31,207,31,207,30,50,31,110,31,225,31,17,31,17,30,190,31,17,31,17,30,42,31,55,31,247,31,190,31,235,31,249,31,249,30,241,31,146,31,189,31,135,31,121,31,128,31,43,31,102,31,246,31,42,31,146,31,146,30,136,31,33,31,201,31,10,31,101,31,77,31,18,31,30,31,232,31,232,30,22,31,27,31,145,31,150,31,16,31,210,31,237,31,163,31,242,31,136,31,136,30,136,29,120,31,141,31,19,31,122,31,25,31,217,31,217,30,142,31,8,31,13,31,15,31,15,30,204,31,140,31,136,31,72,31,72,30,72,29,72,28,178,31,131,31,203,31,111,31,171,31,115,31,78,31,78,30,78,29,7,31,28,31,84,31,84,30,84,29,133,31,39,31,226,31,226,30,156,31,127,31,67,31,114,31,190,31,27,31,17,31,242,31,239,31,254,31,127,31,127,30,154,31,190,31,176,31,204,31,42,31,119,31,119,30,135,31,17,31,17,30,66,31,252,31,213,31,81,31,95,31,194,31,149,31,149,30,102,31,134,31,127,31,73,31,73,30,242,31,11,31,143,31,155,31,75,31,156,31,74,31,203,31,159,31,94,31,94,30,187,31,187,30,72,31,35,31,55,31,55,30,5,31,23,31,128,31,123,31,42,31,13,31,59,31,52,31,165,31,162,31,160,31,125,31,27,31,27,30,135,31,96,31,96,30,51,31,2,31,90,31,90,30,172,31,84,31,63,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
