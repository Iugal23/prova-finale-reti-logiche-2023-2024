-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1017;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (88,0,88,0,242,0,220,0,168,0,0,0,32,0,15,0,244,0,0,0,201,0,0,0,213,0,156,0,157,0,10,0,223,0,0,0,22,0,0,0,166,0,38,0,140,0,152,0,36,0,93,0,194,0,12,0,168,0,168,0,130,0,145,0,80,0,190,0,164,0,8,0,192,0,109,0,227,0,11,0,240,0,60,0,19,0,0,0,172,0,0,0,100,0,31,0,210,0,112,0,103,0,156,0,0,0,27,0,115,0,201,0,235,0,230,0,166,0,175,0,120,0,63,0,0,0,147,0,34,0,43,0,197,0,16,0,153,0,251,0,51,0,0,0,197,0,84,0,196,0,0,0,185,0,80,0,74,0,0,0,191,0,165,0,0,0,22,0,237,0,214,0,32,0,0,0,95,0,90,0,0,0,0,0,205,0,0,0,0,0,35,0,52,0,248,0,51,0,16,0,154,0,43,0,59,0,0,0,219,0,227,0,65,0,30,0,209,0,113,0,213,0,7,0,241,0,189,0,41,0,229,0,124,0,98,0,206,0,244,0,235,0,225,0,101,0,217,0,0,0,218,0,106,0,95,0,0,0,229,0,132,0,73,0,0,0,191,0,134,0,129,0,135,0,0,0,99,0,171,0,249,0,199,0,0,0,0,0,200,0,125,0,246,0,2,0,159,0,0,0,156,0,217,0,71,0,229,0,0,0,215,0,0,0,198,0,201,0,0,0,75,0,56,0,170,0,170,0,43,0,60,0,36,0,0,0,153,0,64,0,89,0,163,0,0,0,140,0,32,0,155,0,55,0,238,0,115,0,137,0,106,0,75,0,0,0,187,0,8,0,159,0,112,0,52,0,181,0,0,0,216,0,188,0,227,0,110,0,154,0,189,0,0,0,0,0,0,0,0,0,0,0,115,0,244,0,61,0,48,0,90,0,223,0,0,0,144,0,150,0,113,0,43,0,171,0,0,0,190,0,0,0,5,0,0,0,159,0,8,0,223,0,154,0,36,0,196,0,153,0,78,0,218,0,25,0,25,0,0,0,185,0,169,0,179,0,0,0,172,0,26,0,235,0,183,0,151,0,225,0,65,0,252,0,77,0,250,0,61,0,0,0,44,0,164,0,231,0,136,0,35,0,64,0,0,0,56,0,46,0,57,0,108,0,0,0,139,0,226,0,185,0,40,0,134,0,133,0,0,0,0,0,52,0,82,0,42,0,178,0,215,0,230,0,63,0,185,0,1,0,0,0,189,0,20,0,235,0,0,0,163,0,0,0,0,0,0,0,195,0,7,0,47,0,12,0,1,0,44,0,124,0,138,0,124,0,0,0,221,0,215,0,0,0,210,0,207,0,0,0,0,0,0,0,187,0,245,0,155,0,123,0,114,0,115,0,124,0,197,0,126,0,94,0,122,0,136,0,136,0,161,0,50,0,253,0,0,0,172,0,196,0,0,0,92,0,113,0,193,0,0,0,244,0,86,0,196,0,10,0,101,0,0,0,225,0,0,0,150,0,91,0,0,0,132,0,132,0,210,0,193,0,239,0,245,0,78,0,28,0,189,0,78,0,144,0,122,0,145,0,76,0,226,0,36,0,0,0,105,0,201,0,155,0,212,0,250,0,234,0,183,0,163,0,199,0,43,0,242,0,151,0,56,0,245,0,103,0,60,0,188,0,0,0,0,0,49,0,121,0,145,0,0,0,0,0,0,0,140,0,0,0,2,0,34,0,157,0,125,0,53,0,228,0,235,0,155,0,189,0,0,0,149,0,142,0,183,0,153,0,33,0,48,0,0,0,38,0,8,0,175,0,25,0,39,0,233,0,215,0,189,0,0,0,0,0,135,0,18,0,44,0,197,0,0,0,128,0,0,0,64,0,47,0,246,0,58,0,0,0,213,0,54,0,103,0,174,0,173,0,177,0,0,0,212,0,183,0,196,0,114,0,78,0,0,0,232,0,209,0,49,0,87,0,212,0,26,0,229,0,12,0,0,0,14,0,162,0,16,0,175,0,198,0,0,0,79,0,70,0,216,0,249,0,0,0,21,0,201,0,255,0,94,0,0,0,194,0,57,0,0,0,5,0,66,0,2,0,210,0,5,0,20,0,0,0,67,0,27,0,90,0,182,0,197,0,149,0,249,0,178,0,191,0,0,0,0,0,190,0,0,0,0,0,0,0,147,0,0,0,48,0,67,0,147,0,223,0,69,0,148,0,107,0,227,0,30,0,45,0,26,0,146,0,138,0,108,0,29,0,198,0,0,0,157,0,228,0,124,0,16,0,238,0,8,0,31,0,157,0,164,0,104,0,0,0,93,0,16,0,0,0,225,0,180,0,0,0,137,0,21,0,227,0,22,0,78,0,126,0,0,0,0,0,100,0,245,0,184,0,200,0,60,0,167,0,56,0,186,0,23,0,0,0,223,0,105,0,197,0,120,0,116,0,75,0,157,0,47,0,0,0,149,0,189,0,0,0,106,0,234,0,165,0,78,0,0,0,30,0,117,0,16,0,70,0,72,0,193,0,36,0,251,0,0,0,227,0,0,0,0,0,159,0,66,0,184,0,76,0,18,0,85,0,103,0,37,0,68,0,134,0,0,0,0,0,0,0,247,0,119,0,0,0,58,0,210,0,116,0,0,0,29,0,218,0,0,0,0,0,0,0,0,0,211,0,103,0,0,0,100,0,148,0,86,0,50,0,188,0,146,0,48,0,223,0,39,0,44,0,146,0,88,0,145,0,163,0,17,0,84,0,170,0,110,0,0,0,132,0,67,0,157,0,0,0,0,0,219,0,182,0,23,0,109,0,2,0,255,0,110,0,124,0,221,0,116,0,228,0,96,0,117,0,121,0,98,0,211,0,43,0,46,0,0,0,92,0,0,0,70,0,78,0,30,0,216,0,0,0,253,0,202,0,163,0,110,0,125,0,227,0,64,0,181,0,80,0,98,0,185,0,152,0,122,0,154,0,11,0,49,0,72,0,124,0,88,0,226,0,0,0,197,0,57,0,177,0,146,0,0,0,0,0,0,0,66,0,51,0,159,0,0,0,180,0,95,0,135,0,13,0,234,0,81,0,219,0,83,0,64,0,83,0,0,0,136,0,136,0,0,0,205,0,198,0,144,0,158,0,189,0,3,0,55,0,151,0,57,0,91,0,0,0,0,0,0,0,0,0,0,0,109,0,0,0,186,0,89,0,255,0,90,0,0,0,41,0,70,0,212,0,148,0,0,0,33,0,107,0,65,0,230,0,241,0,0,0,131,0,225,0,252,0,136,0,94,0,151,0,242,0,13,0,0,0,251,0,89,0,0,0,209,0,170,0,119,0,132,0,156,0,77,0,225,0,0,0,141,0,216,0,0,0,28,0,0,0,0,0,190,0,49,0,33,0,165,0,0,0,38,0,46,0,188,0,235,0,14,0,184,0,145,0,231,0,254,0,253,0,0,0,88,0,0,0,47,0,0,0,181,0,50,0,75,0,218,0,86,0,0,0,183,0,218,0,202,0,53,0,0,0,176,0,38,0,117,0,104,0,0,0,148,0,103,0,61,0,188,0,0,0,176,0,85,0,229,0,227,0,140,0,252,0,244,0,167,0,254,0,0,0,0,0,79,0,0,0,242,0,0,0,188,0,19,0,61,0,77,0,0,0,217,0,10,0,130,0,0,0,168,0,2,0,0,0,0,0,115,0,97,0,68,0,38,0,11,0,91,0,14,0,139,0,0,0,22,0,104,0,88,0,204,0,5,0,98,0,237,0,0,0,227,0,27,0,45,0,85,0,0,0,207,0,140,0,58,0,0,0,96,0,243,0,96,0,71,0,205,0,126,0,35,0,0,0,69,0,205,0,0,0,3,0,151,0,175,0,0,0,0,0,0,0,237,0,243,0,216,0,81,0,242,0,0,0,231,0,12,0,23,0,0,0,51,0,17,0,0,0,236,0,42,0,88,0,239,0,165,0,0,0,234,0,167,0,88,0,74,0,76,0,111,0,247,0,0,0,25,0,232,0,133,0,25,0,118,0,128,0,124,0,57,0,111,0,0,0,0,0,118,0,0,0,0,0,0,0,229,0,22,0,40,0,238,0,52,0,221,0,127,0,222,0,0,0,179,0,173,0,6,0,252,0,243,0,0,0,163,0,178,0,245,0,158,0,148,0,171,0,160,0,0,0,184,0,244,0,233,0,92,0,0,0,108,0,88,0,112,0,0,0,224,0,177,0,174,0,132,0,0,0,219,0,67,0,10,0,0,0,0,0,39,0,117,0,0,0,15,0,251,0,204,0,0,0,0,0,123,0,128,0,130,0,29,0,124,0,138,0,90,0,125,0,0,0,138,0,42,0,91,0,0,0,28,0,109,0,70,0,0,0,217,0,196,0,52,0,35,0,68,0,73,0,144,0,0,0,118,0,0,0,0,0,73,0,201,0,159,0,174,0,12,0,205,0,65,0,53,0,0,0,173,0,137,0,250,0,147,0,150,0,0,0,172,0,189,0,248,0,209,0,41,0,220,0,0,0,62,0,0,0,97,0,6,0,205,0,0,0,28,0,95,0,0,0,0,0,62,0,239,0,0,0);
signal scenario_full  : scenario_type := (88,31,88,31,242,31,220,31,168,31,168,30,32,31,15,31,244,31,244,30,201,31,201,30,213,31,156,31,157,31,10,31,223,31,223,30,22,31,22,30,166,31,38,31,140,31,152,31,36,31,93,31,194,31,12,31,168,31,168,31,130,31,145,31,80,31,190,31,164,31,8,31,192,31,109,31,227,31,11,31,240,31,60,31,19,31,19,30,172,31,172,30,100,31,31,31,210,31,112,31,103,31,156,31,156,30,27,31,115,31,201,31,235,31,230,31,166,31,175,31,120,31,63,31,63,30,147,31,34,31,43,31,197,31,16,31,153,31,251,31,51,31,51,30,197,31,84,31,196,31,196,30,185,31,80,31,74,31,74,30,191,31,165,31,165,30,22,31,237,31,214,31,32,31,32,30,95,31,90,31,90,30,90,29,205,31,205,30,205,29,35,31,52,31,248,31,51,31,16,31,154,31,43,31,59,31,59,30,219,31,227,31,65,31,30,31,209,31,113,31,213,31,7,31,241,31,189,31,41,31,229,31,124,31,98,31,206,31,244,31,235,31,225,31,101,31,217,31,217,30,218,31,106,31,95,31,95,30,229,31,132,31,73,31,73,30,191,31,134,31,129,31,135,31,135,30,99,31,171,31,249,31,199,31,199,30,199,29,200,31,125,31,246,31,2,31,159,31,159,30,156,31,217,31,71,31,229,31,229,30,215,31,215,30,198,31,201,31,201,30,75,31,56,31,170,31,170,31,43,31,60,31,36,31,36,30,153,31,64,31,89,31,163,31,163,30,140,31,32,31,155,31,55,31,238,31,115,31,137,31,106,31,75,31,75,30,187,31,8,31,159,31,112,31,52,31,181,31,181,30,216,31,188,31,227,31,110,31,154,31,189,31,189,30,189,29,189,28,189,27,189,26,115,31,244,31,61,31,48,31,90,31,223,31,223,30,144,31,150,31,113,31,43,31,171,31,171,30,190,31,190,30,5,31,5,30,159,31,8,31,223,31,154,31,36,31,196,31,153,31,78,31,218,31,25,31,25,31,25,30,185,31,169,31,179,31,179,30,172,31,26,31,235,31,183,31,151,31,225,31,65,31,252,31,77,31,250,31,61,31,61,30,44,31,164,31,231,31,136,31,35,31,64,31,64,30,56,31,46,31,57,31,108,31,108,30,139,31,226,31,185,31,40,31,134,31,133,31,133,30,133,29,52,31,82,31,42,31,178,31,215,31,230,31,63,31,185,31,1,31,1,30,189,31,20,31,235,31,235,30,163,31,163,30,163,29,163,28,195,31,7,31,47,31,12,31,1,31,44,31,124,31,138,31,124,31,124,30,221,31,215,31,215,30,210,31,207,31,207,30,207,29,207,28,187,31,245,31,155,31,123,31,114,31,115,31,124,31,197,31,126,31,94,31,122,31,136,31,136,31,161,31,50,31,253,31,253,30,172,31,196,31,196,30,92,31,113,31,193,31,193,30,244,31,86,31,196,31,10,31,101,31,101,30,225,31,225,30,150,31,91,31,91,30,132,31,132,31,210,31,193,31,239,31,245,31,78,31,28,31,189,31,78,31,144,31,122,31,145,31,76,31,226,31,36,31,36,30,105,31,201,31,155,31,212,31,250,31,234,31,183,31,163,31,199,31,43,31,242,31,151,31,56,31,245,31,103,31,60,31,188,31,188,30,188,29,49,31,121,31,145,31,145,30,145,29,145,28,140,31,140,30,2,31,34,31,157,31,125,31,53,31,228,31,235,31,155,31,189,31,189,30,149,31,142,31,183,31,153,31,33,31,48,31,48,30,38,31,8,31,175,31,25,31,39,31,233,31,215,31,189,31,189,30,189,29,135,31,18,31,44,31,197,31,197,30,128,31,128,30,64,31,47,31,246,31,58,31,58,30,213,31,54,31,103,31,174,31,173,31,177,31,177,30,212,31,183,31,196,31,114,31,78,31,78,30,232,31,209,31,49,31,87,31,212,31,26,31,229,31,12,31,12,30,14,31,162,31,16,31,175,31,198,31,198,30,79,31,70,31,216,31,249,31,249,30,21,31,201,31,255,31,94,31,94,30,194,31,57,31,57,30,5,31,66,31,2,31,210,31,5,31,20,31,20,30,67,31,27,31,90,31,182,31,197,31,149,31,249,31,178,31,191,31,191,30,191,29,190,31,190,30,190,29,190,28,147,31,147,30,48,31,67,31,147,31,223,31,69,31,148,31,107,31,227,31,30,31,45,31,26,31,146,31,138,31,108,31,29,31,198,31,198,30,157,31,228,31,124,31,16,31,238,31,8,31,31,31,157,31,164,31,104,31,104,30,93,31,16,31,16,30,225,31,180,31,180,30,137,31,21,31,227,31,22,31,78,31,126,31,126,30,126,29,100,31,245,31,184,31,200,31,60,31,167,31,56,31,186,31,23,31,23,30,223,31,105,31,197,31,120,31,116,31,75,31,157,31,47,31,47,30,149,31,189,31,189,30,106,31,234,31,165,31,78,31,78,30,30,31,117,31,16,31,70,31,72,31,193,31,36,31,251,31,251,30,227,31,227,30,227,29,159,31,66,31,184,31,76,31,18,31,85,31,103,31,37,31,68,31,134,31,134,30,134,29,134,28,247,31,119,31,119,30,58,31,210,31,116,31,116,30,29,31,218,31,218,30,218,29,218,28,218,27,211,31,103,31,103,30,100,31,148,31,86,31,50,31,188,31,146,31,48,31,223,31,39,31,44,31,146,31,88,31,145,31,163,31,17,31,84,31,170,31,110,31,110,30,132,31,67,31,157,31,157,30,157,29,219,31,182,31,23,31,109,31,2,31,255,31,110,31,124,31,221,31,116,31,228,31,96,31,117,31,121,31,98,31,211,31,43,31,46,31,46,30,92,31,92,30,70,31,78,31,30,31,216,31,216,30,253,31,202,31,163,31,110,31,125,31,227,31,64,31,181,31,80,31,98,31,185,31,152,31,122,31,154,31,11,31,49,31,72,31,124,31,88,31,226,31,226,30,197,31,57,31,177,31,146,31,146,30,146,29,146,28,66,31,51,31,159,31,159,30,180,31,95,31,135,31,13,31,234,31,81,31,219,31,83,31,64,31,83,31,83,30,136,31,136,31,136,30,205,31,198,31,144,31,158,31,189,31,3,31,55,31,151,31,57,31,91,31,91,30,91,29,91,28,91,27,91,26,109,31,109,30,186,31,89,31,255,31,90,31,90,30,41,31,70,31,212,31,148,31,148,30,33,31,107,31,65,31,230,31,241,31,241,30,131,31,225,31,252,31,136,31,94,31,151,31,242,31,13,31,13,30,251,31,89,31,89,30,209,31,170,31,119,31,132,31,156,31,77,31,225,31,225,30,141,31,216,31,216,30,28,31,28,30,28,29,190,31,49,31,33,31,165,31,165,30,38,31,46,31,188,31,235,31,14,31,184,31,145,31,231,31,254,31,253,31,253,30,88,31,88,30,47,31,47,30,181,31,50,31,75,31,218,31,86,31,86,30,183,31,218,31,202,31,53,31,53,30,176,31,38,31,117,31,104,31,104,30,148,31,103,31,61,31,188,31,188,30,176,31,85,31,229,31,227,31,140,31,252,31,244,31,167,31,254,31,254,30,254,29,79,31,79,30,242,31,242,30,188,31,19,31,61,31,77,31,77,30,217,31,10,31,130,31,130,30,168,31,2,31,2,30,2,29,115,31,97,31,68,31,38,31,11,31,91,31,14,31,139,31,139,30,22,31,104,31,88,31,204,31,5,31,98,31,237,31,237,30,227,31,27,31,45,31,85,31,85,30,207,31,140,31,58,31,58,30,96,31,243,31,96,31,71,31,205,31,126,31,35,31,35,30,69,31,205,31,205,30,3,31,151,31,175,31,175,30,175,29,175,28,237,31,243,31,216,31,81,31,242,31,242,30,231,31,12,31,23,31,23,30,51,31,17,31,17,30,236,31,42,31,88,31,239,31,165,31,165,30,234,31,167,31,88,31,74,31,76,31,111,31,247,31,247,30,25,31,232,31,133,31,25,31,118,31,128,31,124,31,57,31,111,31,111,30,111,29,118,31,118,30,118,29,118,28,229,31,22,31,40,31,238,31,52,31,221,31,127,31,222,31,222,30,179,31,173,31,6,31,252,31,243,31,243,30,163,31,178,31,245,31,158,31,148,31,171,31,160,31,160,30,184,31,244,31,233,31,92,31,92,30,108,31,88,31,112,31,112,30,224,31,177,31,174,31,132,31,132,30,219,31,67,31,10,31,10,30,10,29,39,31,117,31,117,30,15,31,251,31,204,31,204,30,204,29,123,31,128,31,130,31,29,31,124,31,138,31,90,31,125,31,125,30,138,31,42,31,91,31,91,30,28,31,109,31,70,31,70,30,217,31,196,31,52,31,35,31,68,31,73,31,144,31,144,30,118,31,118,30,118,29,73,31,201,31,159,31,174,31,12,31,205,31,65,31,53,31,53,30,173,31,137,31,250,31,147,31,150,31,150,30,172,31,189,31,248,31,209,31,41,31,220,31,220,30,62,31,62,30,97,31,6,31,205,31,205,30,28,31,95,31,95,30,95,29,62,31,239,31,239,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
