-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_236 is
end project_tb_236;

architecture project_tb_arch_236 of project_tb_236 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 912;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (232,0,197,0,79,0,0,0,0,0,10,0,140,0,164,0,86,0,194,0,243,0,158,0,0,0,144,0,120,0,185,0,231,0,23,0,195,0,22,0,224,0,0,0,73,0,90,0,123,0,1,0,0,0,5,0,208,0,0,0,183,0,142,0,142,0,95,0,255,0,171,0,37,0,47,0,71,0,53,0,155,0,38,0,226,0,167,0,155,0,203,0,252,0,231,0,4,0,151,0,229,0,0,0,0,0,68,0,0,0,126,0,211,0,27,0,236,0,209,0,77,0,96,0,0,0,254,0,215,0,127,0,51,0,103,0,209,0,0,0,82,0,35,0,48,0,4,0,71,0,141,0,249,0,194,0,28,0,0,0,57,0,169,0,62,0,215,0,178,0,0,0,187,0,117,0,213,0,153,0,9,0,94,0,61,0,0,0,5,0,113,0,16,0,255,0,45,0,109,0,175,0,76,0,220,0,127,0,233,0,5,0,161,0,0,0,34,0,188,0,135,0,136,0,48,0,61,0,113,0,245,0,197,0,243,0,221,0,178,0,151,0,130,0,238,0,240,0,211,0,235,0,197,0,0,0,68,0,0,0,192,0,148,0,191,0,109,0,0,0,172,0,125,0,0,0,189,0,80,0,129,0,150,0,132,0,144,0,33,0,36,0,232,0,0,0,91,0,151,0,128,0,245,0,89,0,172,0,254,0,0,0,7,0,30,0,35,0,185,0,100,0,0,0,29,0,226,0,76,0,151,0,211,0,2,0,120,0,0,0,50,0,243,0,191,0,62,0,81,0,0,0,125,0,240,0,186,0,118,0,0,0,59,0,133,0,184,0,32,0,0,0,0,0,249,0,0,0,224,0,62,0,0,0,0,0,28,0,86,0,63,0,74,0,178,0,33,0,196,0,121,0,14,0,9,0,228,0,134,0,193,0,116,0,196,0,204,0,0,0,58,0,0,0,123,0,79,0,36,0,0,0,114,0,0,0,118,0,213,0,158,0,0,0,0,0,71,0,187,0,23,0,118,0,120,0,241,0,6,0,247,0,126,0,0,0,50,0,53,0,229,0,158,0,0,0,0,0,0,0,0,0,205,0,150,0,178,0,95,0,87,0,0,0,84,0,0,0,173,0,36,0,175,0,49,0,139,0,124,0,128,0,65,0,171,0,175,0,191,0,219,0,188,0,73,0,27,0,0,0,0,0,60,0,231,0,175,0,0,0,109,0,195,0,70,0,17,0,0,0,109,0,194,0,86,0,167,0,120,0,227,0,102,0,178,0,20,0,81,0,56,0,239,0,194,0,233,0,167,0,217,0,110,0,68,0,13,0,0,0,77,0,140,0,52,0,2,0,82,0,81,0,133,0,10,0,231,0,91,0,0,0,119,0,221,0,225,0,84,0,40,0,64,0,206,0,241,0,156,0,172,0,0,0,130,0,235,0,194,0,217,0,47,0,197,0,160,0,0,0,65,0,0,0,107,0,94,0,0,0,38,0,191,0,74,0,200,0,70,0,228,0,96,0,189,0,61,0,10,0,195,0,5,0,221,0,157,0,0,0,191,0,164,0,0,0,17,0,246,0,0,0,195,0,85,0,162,0,0,0,103,0,0,0,253,0,222,0,0,0,225,0,151,0,0,0,168,0,229,0,210,0,0,0,163,0,221,0,174,0,106,0,127,0,71,0,49,0,70,0,0,0,0,0,248,0,136,0,183,0,148,0,138,0,83,0,100,0,20,0,207,0,108,0,155,0,208,0,13,0,156,0,78,0,17,0,110,0,164,0,0,0,0,0,2,0,0,0,109,0,84,0,166,0,60,0,132,0,80,0,0,0,156,0,222,0,33,0,37,0,173,0,211,0,106,0,223,0,214,0,233,0,194,0,57,0,224,0,133,0,73,0,83,0,105,0,251,0,115,0,253,0,32,0,76,0,179,0,222,0,247,0,170,0,123,0,209,0,132,0,164,0,204,0,84,0,50,0,0,0,180,0,95,0,44,0,0,0,71,0,42,0,0,0,85,0,147,0,242,0,18,0,0,0,0,0,0,0,241,0,172,0,0,0,36,0,157,0,222,0,223,0,0,0,103,0,0,0,0,0,0,0,112,0,252,0,223,0,28,0,205,0,216,0,168,0,23,0,122,0,196,0,0,0,195,0,22,0,120,0,157,0,0,0,236,0,0,0,0,0,211,0,0,0,0,0,183,0,177,0,24,0,0,0,57,0,61,0,5,0,0,0,11,0,167,0,62,0,131,0,244,0,78,0,56,0,49,0,180,0,97,0,203,0,128,0,0,0,160,0,162,0,167,0,90,0,0,0,193,0,245,0,171,0,0,0,105,0,244,0,57,0,172,0,227,0,239,0,184,0,77,0,225,0,0,0,38,0,248,0,158,0,49,0,70,0,254,0,86,0,195,0,179,0,215,0,68,0,185,0,129,0,145,0,0,0,0,0,99,0,162,0,71,0,0,0,240,0,90,0,195,0,161,0,0,0,107,0,49,0,0,0,185,0,21,0,153,0,43,0,151,0,10,0,154,0,99,0,195,0,170,0,69,0,10,0,237,0,176,0,0,0,176,0,121,0,0,0,0,0,37,0,97,0,99,0,35,0,0,0,103,0,0,0,209,0,192,0,149,0,115,0,38,0,32,0,34,0,0,0,115,0,169,0,225,0,48,0,148,0,218,0,52,0,21,0,0,0,48,0,252,0,128,0,44,0,126,0,64,0,14,0,230,0,87,0,13,0,129,0,202,0,113,0,0,0,0,0,223,0,160,0,115,0,217,0,157,0,34,0,214,0,101,0,94,0,8,0,82,0,68,0,116,0,0,0,223,0,67,0,83,0,149,0,40,0,153,0,70,0,210,0,58,0,0,0,136,0,158,0,0,0,182,0,0,0,27,0,36,0,234,0,195,0,229,0,41,0,243,0,83,0,93,0,0,0,4,0,166,0,194,0,171,0,88,0,143,0,0,0,227,0,143,0,8,0,245,0,109,0,0,0,29,0,0,0,218,0,80,0,52,0,65,0,46,0,70,0,0,0,98,0,186,0,157,0,184,0,48,0,112,0,218,0,35,0,45,0,3,0,109,0,117,0,0,0,101,0,0,0,57,0,40,0,237,0,153,0,59,0,133,0,45,0,0,0,0,0,82,0,27,0,209,0,28,0,0,0,97,0,0,0,98,0,11,0,0,0,207,0,247,0,120,0,54,0,6,0,0,0,120,0,37,0,40,0,35,0,189,0,132,0,17,0,125,0,90,0,48,0,166,0,233,0,202,0,159,0,32,0,136,0,176,0,90,0,209,0,74,0,168,0,137,0,32,0,0,0,251,0,74,0,0,0,151,0,69,0,0,0,0,0,161,0,83,0,146,0,123,0,0,0,0,0,0,0,52,0,0,0,75,0,205,0,170,0,118,0,110,0,14,0,31,0,0,0,0,0,99,0,70,0,0,0,0,0,46,0,115,0,176,0,55,0,0,0,215,0,235,0,199,0,99,0,45,0,205,0,109,0,32,0,56,0,246,0,61,0,0,0,102,0,253,0,227,0,242,0,88,0,0,0,0,0,27,0,170,0,226,0,201,0,156,0,163,0,104,0,0,0,58,0,48,0,228,0,2,0,168,0,31,0,43,0,45,0,170,0,8,0,253,0,57,0,255,0,69,0,0,0,37,0,230,0,0,0,175,0,20,0,0,0,166,0,114,0,34,0,189,0,185,0,14,0,170,0,95,0,199,0,1,0,138,0,116,0,8,0,30,0,232,0,46,0,0,0,28,0,147,0,217,0,199,0,26,0,214,0,0,0,78,0,109,0,225,0,92,0,148,0,0,0,112,0,247,0,42,0,51,0,171,0,115,0,1,0,0,0,0,0,0,0,0,0,131,0,111,0,42,0,79,0,45,0,36,0,65,0,83,0,111,0,81,0,27,0,43,0,100,0,18,0,50,0,253,0,253,0,168,0,33,0,74,0,188,0,161,0,97,0,169,0,162,0,70,0,249,0,161,0,155,0,140,0,211,0,14,0,253,0,252,0,201,0,202,0,242,0,96,0,10,0,145,0,81,0,208,0,0,0,0,0,219,0,0,0,144,0,138,0,132,0,0,0);
signal scenario_full  : scenario_type := (232,31,197,31,79,31,79,30,79,29,10,31,140,31,164,31,86,31,194,31,243,31,158,31,158,30,144,31,120,31,185,31,231,31,23,31,195,31,22,31,224,31,224,30,73,31,90,31,123,31,1,31,1,30,5,31,208,31,208,30,183,31,142,31,142,31,95,31,255,31,171,31,37,31,47,31,71,31,53,31,155,31,38,31,226,31,167,31,155,31,203,31,252,31,231,31,4,31,151,31,229,31,229,30,229,29,68,31,68,30,126,31,211,31,27,31,236,31,209,31,77,31,96,31,96,30,254,31,215,31,127,31,51,31,103,31,209,31,209,30,82,31,35,31,48,31,4,31,71,31,141,31,249,31,194,31,28,31,28,30,57,31,169,31,62,31,215,31,178,31,178,30,187,31,117,31,213,31,153,31,9,31,94,31,61,31,61,30,5,31,113,31,16,31,255,31,45,31,109,31,175,31,76,31,220,31,127,31,233,31,5,31,161,31,161,30,34,31,188,31,135,31,136,31,48,31,61,31,113,31,245,31,197,31,243,31,221,31,178,31,151,31,130,31,238,31,240,31,211,31,235,31,197,31,197,30,68,31,68,30,192,31,148,31,191,31,109,31,109,30,172,31,125,31,125,30,189,31,80,31,129,31,150,31,132,31,144,31,33,31,36,31,232,31,232,30,91,31,151,31,128,31,245,31,89,31,172,31,254,31,254,30,7,31,30,31,35,31,185,31,100,31,100,30,29,31,226,31,76,31,151,31,211,31,2,31,120,31,120,30,50,31,243,31,191,31,62,31,81,31,81,30,125,31,240,31,186,31,118,31,118,30,59,31,133,31,184,31,32,31,32,30,32,29,249,31,249,30,224,31,62,31,62,30,62,29,28,31,86,31,63,31,74,31,178,31,33,31,196,31,121,31,14,31,9,31,228,31,134,31,193,31,116,31,196,31,204,31,204,30,58,31,58,30,123,31,79,31,36,31,36,30,114,31,114,30,118,31,213,31,158,31,158,30,158,29,71,31,187,31,23,31,118,31,120,31,241,31,6,31,247,31,126,31,126,30,50,31,53,31,229,31,158,31,158,30,158,29,158,28,158,27,205,31,150,31,178,31,95,31,87,31,87,30,84,31,84,30,173,31,36,31,175,31,49,31,139,31,124,31,128,31,65,31,171,31,175,31,191,31,219,31,188,31,73,31,27,31,27,30,27,29,60,31,231,31,175,31,175,30,109,31,195,31,70,31,17,31,17,30,109,31,194,31,86,31,167,31,120,31,227,31,102,31,178,31,20,31,81,31,56,31,239,31,194,31,233,31,167,31,217,31,110,31,68,31,13,31,13,30,77,31,140,31,52,31,2,31,82,31,81,31,133,31,10,31,231,31,91,31,91,30,119,31,221,31,225,31,84,31,40,31,64,31,206,31,241,31,156,31,172,31,172,30,130,31,235,31,194,31,217,31,47,31,197,31,160,31,160,30,65,31,65,30,107,31,94,31,94,30,38,31,191,31,74,31,200,31,70,31,228,31,96,31,189,31,61,31,10,31,195,31,5,31,221,31,157,31,157,30,191,31,164,31,164,30,17,31,246,31,246,30,195,31,85,31,162,31,162,30,103,31,103,30,253,31,222,31,222,30,225,31,151,31,151,30,168,31,229,31,210,31,210,30,163,31,221,31,174,31,106,31,127,31,71,31,49,31,70,31,70,30,70,29,248,31,136,31,183,31,148,31,138,31,83,31,100,31,20,31,207,31,108,31,155,31,208,31,13,31,156,31,78,31,17,31,110,31,164,31,164,30,164,29,2,31,2,30,109,31,84,31,166,31,60,31,132,31,80,31,80,30,156,31,222,31,33,31,37,31,173,31,211,31,106,31,223,31,214,31,233,31,194,31,57,31,224,31,133,31,73,31,83,31,105,31,251,31,115,31,253,31,32,31,76,31,179,31,222,31,247,31,170,31,123,31,209,31,132,31,164,31,204,31,84,31,50,31,50,30,180,31,95,31,44,31,44,30,71,31,42,31,42,30,85,31,147,31,242,31,18,31,18,30,18,29,18,28,241,31,172,31,172,30,36,31,157,31,222,31,223,31,223,30,103,31,103,30,103,29,103,28,112,31,252,31,223,31,28,31,205,31,216,31,168,31,23,31,122,31,196,31,196,30,195,31,22,31,120,31,157,31,157,30,236,31,236,30,236,29,211,31,211,30,211,29,183,31,177,31,24,31,24,30,57,31,61,31,5,31,5,30,11,31,167,31,62,31,131,31,244,31,78,31,56,31,49,31,180,31,97,31,203,31,128,31,128,30,160,31,162,31,167,31,90,31,90,30,193,31,245,31,171,31,171,30,105,31,244,31,57,31,172,31,227,31,239,31,184,31,77,31,225,31,225,30,38,31,248,31,158,31,49,31,70,31,254,31,86,31,195,31,179,31,215,31,68,31,185,31,129,31,145,31,145,30,145,29,99,31,162,31,71,31,71,30,240,31,90,31,195,31,161,31,161,30,107,31,49,31,49,30,185,31,21,31,153,31,43,31,151,31,10,31,154,31,99,31,195,31,170,31,69,31,10,31,237,31,176,31,176,30,176,31,121,31,121,30,121,29,37,31,97,31,99,31,35,31,35,30,103,31,103,30,209,31,192,31,149,31,115,31,38,31,32,31,34,31,34,30,115,31,169,31,225,31,48,31,148,31,218,31,52,31,21,31,21,30,48,31,252,31,128,31,44,31,126,31,64,31,14,31,230,31,87,31,13,31,129,31,202,31,113,31,113,30,113,29,223,31,160,31,115,31,217,31,157,31,34,31,214,31,101,31,94,31,8,31,82,31,68,31,116,31,116,30,223,31,67,31,83,31,149,31,40,31,153,31,70,31,210,31,58,31,58,30,136,31,158,31,158,30,182,31,182,30,27,31,36,31,234,31,195,31,229,31,41,31,243,31,83,31,93,31,93,30,4,31,166,31,194,31,171,31,88,31,143,31,143,30,227,31,143,31,8,31,245,31,109,31,109,30,29,31,29,30,218,31,80,31,52,31,65,31,46,31,70,31,70,30,98,31,186,31,157,31,184,31,48,31,112,31,218,31,35,31,45,31,3,31,109,31,117,31,117,30,101,31,101,30,57,31,40,31,237,31,153,31,59,31,133,31,45,31,45,30,45,29,82,31,27,31,209,31,28,31,28,30,97,31,97,30,98,31,11,31,11,30,207,31,247,31,120,31,54,31,6,31,6,30,120,31,37,31,40,31,35,31,189,31,132,31,17,31,125,31,90,31,48,31,166,31,233,31,202,31,159,31,32,31,136,31,176,31,90,31,209,31,74,31,168,31,137,31,32,31,32,30,251,31,74,31,74,30,151,31,69,31,69,30,69,29,161,31,83,31,146,31,123,31,123,30,123,29,123,28,52,31,52,30,75,31,205,31,170,31,118,31,110,31,14,31,31,31,31,30,31,29,99,31,70,31,70,30,70,29,46,31,115,31,176,31,55,31,55,30,215,31,235,31,199,31,99,31,45,31,205,31,109,31,32,31,56,31,246,31,61,31,61,30,102,31,253,31,227,31,242,31,88,31,88,30,88,29,27,31,170,31,226,31,201,31,156,31,163,31,104,31,104,30,58,31,48,31,228,31,2,31,168,31,31,31,43,31,45,31,170,31,8,31,253,31,57,31,255,31,69,31,69,30,37,31,230,31,230,30,175,31,20,31,20,30,166,31,114,31,34,31,189,31,185,31,14,31,170,31,95,31,199,31,1,31,138,31,116,31,8,31,30,31,232,31,46,31,46,30,28,31,147,31,217,31,199,31,26,31,214,31,214,30,78,31,109,31,225,31,92,31,148,31,148,30,112,31,247,31,42,31,51,31,171,31,115,31,1,31,1,30,1,29,1,28,1,27,131,31,111,31,42,31,79,31,45,31,36,31,65,31,83,31,111,31,81,31,27,31,43,31,100,31,18,31,50,31,253,31,253,31,168,31,33,31,74,31,188,31,161,31,97,31,169,31,162,31,70,31,249,31,161,31,155,31,140,31,211,31,14,31,253,31,252,31,201,31,202,31,242,31,96,31,10,31,145,31,81,31,208,31,208,30,208,29,219,31,219,30,144,31,138,31,132,31,132,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
