-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 628;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,235,0,0,0,0,0,200,0,141,0,0,0,0,0,103,0,251,0,120,0,242,0,54,0,0,0,182,0,116,0,246,0,145,0,0,0,86,0,218,0,0,0,73,0,0,0,140,0,1,0,23,0,0,0,0,0,0,0,0,0,191,0,174,0,22,0,0,0,228,0,222,0,206,0,0,0,152,0,99,0,128,0,210,0,127,0,195,0,61,0,85,0,58,0,0,0,7,0,134,0,57,0,137,0,231,0,224,0,56,0,117,0,152,0,0,0,204,0,243,0,72,0,222,0,214,0,28,0,0,0,0,0,95,0,0,0,247,0,114,0,171,0,21,0,217,0,63,0,120,0,189,0,0,0,0,0,58,0,60,0,118,0,61,0,0,0,99,0,0,0,82,0,0,0,37,0,138,0,161,0,147,0,170,0,205,0,98,0,84,0,36,0,211,0,193,0,134,0,161,0,55,0,207,0,188,0,130,0,132,0,0,0,0,0,241,0,25,0,13,0,0,0,140,0,155,0,103,0,0,0,150,0,0,0,108,0,144,0,250,0,116,0,0,0,1,0,198,0,172,0,55,0,36,0,16,0,218,0,54,0,37,0,169,0,209,0,186,0,96,0,87,0,217,0,252,0,228,0,82,0,162,0,88,0,170,0,161,0,0,0,64,0,11,0,192,0,0,0,36,0,16,0,2,0,176,0,84,0,63,0,0,0,57,0,49,0,109,0,0,0,246,0,90,0,176,0,0,0,198,0,25,0,93,0,56,0,162,0,32,0,122,0,85,0,25,0,36,0,249,0,79,0,203,0,25,0,176,0,84,0,204,0,0,0,226,0,72,0,56,0,54,0,151,0,120,0,0,0,0,0,220,0,114,0,181,0,138,0,79,0,246,0,0,0,0,0,0,0,110,0,166,0,172,0,126,0,11,0,226,0,40,0,218,0,75,0,37,0,0,0,45,0,65,0,115,0,57,0,0,0,63,0,110,0,123,0,31,0,165,0,62,0,199,0,193,0,101,0,183,0,129,0,0,0,63,0,170,0,159,0,243,0,28,0,0,0,166,0,62,0,66,0,243,0,56,0,51,0,0,0,34,0,0,0,0,0,95,0,152,0,88,0,75,0,88,0,0,0,7,0,177,0,45,0,201,0,179,0,121,0,88,0,5,0,0,0,0,0,181,0,0,0,35,0,1,0,20,0,243,0,110,0,222,0,244,0,0,0,0,0,0,0,0,0,154,0,74,0,119,0,0,0,0,0,0,0,89,0,125,0,0,0,0,0,0,0,151,0,0,0,117,0,217,0,63,0,218,0,103,0,0,0,8,0,188,0,0,0,238,0,0,0,0,0,241,0,112,0,4,0,96,0,118,0,145,0,35,0,183,0,0,0,247,0,244,0,26,0,247,0,229,0,243,0,140,0,200,0,0,0,153,0,5,0,130,0,193,0,153,0,0,0,147,0,170,0,0,0,123,0,94,0,238,0,223,0,195,0,107,0,169,0,164,0,194,0,216,0,106,0,138,0,209,0,10,0,8,0,100,0,106,0,11,0,206,0,234,0,188,0,0,0,0,0,113,0,193,0,187,0,65,0,246,0,53,0,0,0,34,0,128,0,94,0,115,0,42,0,105,0,0,0,45,0,73,0,0,0,212,0,135,0,158,0,73,0,165,0,209,0,253,0,7,0,239,0,209,0,0,0,0,0,91,0,171,0,116,0,75,0,8,0,56,0,96,0,66,0,213,0,88,0,17,0,27,0,0,0,54,0,0,0,217,0,0,0,97,0,248,0,0,0,195,0,15,0,252,0,198,0,246,0,39,0,239,0,60,0,251,0,0,0,169,0,0,0,191,0,18,0,16,0,249,0,0,0,110,0,24,0,76,0,151,0,250,0,152,0,139,0,204,0,0,0,141,0,165,0,90,0,0,0,0,0,65,0,108,0,190,0,198,0,7,0,232,0,3,0,205,0,249,0,7,0,183,0,253,0,21,0,235,0,70,0,100,0,167,0,151,0,0,0,36,0,96,0,177,0,17,0,75,0,0,0,242,0,78,0,209,0,180,0,61,0,250,0,140,0,16,0,73,0,3,0,221,0,205,0,0,0,50,0,67,0,13,0,99,0,2,0,0,0,0,0,204,0,0,0,255,0,0,0,88,0,88,0,0,0,200,0,235,0,166,0,109,0,35,0,125,0,116,0,53,0,190,0,55,0,47,0,181,0,104,0,16,0,45,0,234,0,225,0,159,0,222,0,113,0,98,0,111,0,0,0,182,0,2,0,53,0,0,0,0,0,251,0,205,0,110,0,112,0,162,0,12,0,237,0,203,0,251,0,0,0,14,0,61,0,40,0,90,0,107,0,0,0,82,0,94,0,248,0,241,0,59,0,29,0,35,0,204,0,188,0,0,0,0,0,104,0,24,0,186,0,0,0,61,0,245,0,88,0,83,0,197,0,152,0,0,0,26,0,184,0,0,0,50,0,84,0,0,0,255,0,162,0,158,0,96,0,38,0,187,0,5,0,12,0,144,0,111,0,0,0,0,0,60,0,187,0,222,0,117,0,43,0,49,0,227,0,188,0,0,0,131,0,60,0,121,0,245,0,237,0,173,0,160,0,139,0,0,0,214,0,217,0,230,0,232,0,17,0,0,0,216,0,0,0,50,0,219,0,47,0,7,0,105,0,198,0,17,0,200,0,191,0,14,0,0,0,112,0,9,0,192,0,240,0,39,0,35,0,114,0,0,0,0,0,115,0,0,0,150,0,138,0,59,0,236,0,226,0,102,0,34,0,178,0,127,0,157,0,70,0,137,0,0,0,241,0,84,0,51,0);
signal scenario_full  : scenario_type := (0,0,235,31,235,30,235,29,200,31,141,31,141,30,141,29,103,31,251,31,120,31,242,31,54,31,54,30,182,31,116,31,246,31,145,31,145,30,86,31,218,31,218,30,73,31,73,30,140,31,1,31,23,31,23,30,23,29,23,28,23,27,191,31,174,31,22,31,22,30,228,31,222,31,206,31,206,30,152,31,99,31,128,31,210,31,127,31,195,31,61,31,85,31,58,31,58,30,7,31,134,31,57,31,137,31,231,31,224,31,56,31,117,31,152,31,152,30,204,31,243,31,72,31,222,31,214,31,28,31,28,30,28,29,95,31,95,30,247,31,114,31,171,31,21,31,217,31,63,31,120,31,189,31,189,30,189,29,58,31,60,31,118,31,61,31,61,30,99,31,99,30,82,31,82,30,37,31,138,31,161,31,147,31,170,31,205,31,98,31,84,31,36,31,211,31,193,31,134,31,161,31,55,31,207,31,188,31,130,31,132,31,132,30,132,29,241,31,25,31,13,31,13,30,140,31,155,31,103,31,103,30,150,31,150,30,108,31,144,31,250,31,116,31,116,30,1,31,198,31,172,31,55,31,36,31,16,31,218,31,54,31,37,31,169,31,209,31,186,31,96,31,87,31,217,31,252,31,228,31,82,31,162,31,88,31,170,31,161,31,161,30,64,31,11,31,192,31,192,30,36,31,16,31,2,31,176,31,84,31,63,31,63,30,57,31,49,31,109,31,109,30,246,31,90,31,176,31,176,30,198,31,25,31,93,31,56,31,162,31,32,31,122,31,85,31,25,31,36,31,249,31,79,31,203,31,25,31,176,31,84,31,204,31,204,30,226,31,72,31,56,31,54,31,151,31,120,31,120,30,120,29,220,31,114,31,181,31,138,31,79,31,246,31,246,30,246,29,246,28,110,31,166,31,172,31,126,31,11,31,226,31,40,31,218,31,75,31,37,31,37,30,45,31,65,31,115,31,57,31,57,30,63,31,110,31,123,31,31,31,165,31,62,31,199,31,193,31,101,31,183,31,129,31,129,30,63,31,170,31,159,31,243,31,28,31,28,30,166,31,62,31,66,31,243,31,56,31,51,31,51,30,34,31,34,30,34,29,95,31,152,31,88,31,75,31,88,31,88,30,7,31,177,31,45,31,201,31,179,31,121,31,88,31,5,31,5,30,5,29,181,31,181,30,35,31,1,31,20,31,243,31,110,31,222,31,244,31,244,30,244,29,244,28,244,27,154,31,74,31,119,31,119,30,119,29,119,28,89,31,125,31,125,30,125,29,125,28,151,31,151,30,117,31,217,31,63,31,218,31,103,31,103,30,8,31,188,31,188,30,238,31,238,30,238,29,241,31,112,31,4,31,96,31,118,31,145,31,35,31,183,31,183,30,247,31,244,31,26,31,247,31,229,31,243,31,140,31,200,31,200,30,153,31,5,31,130,31,193,31,153,31,153,30,147,31,170,31,170,30,123,31,94,31,238,31,223,31,195,31,107,31,169,31,164,31,194,31,216,31,106,31,138,31,209,31,10,31,8,31,100,31,106,31,11,31,206,31,234,31,188,31,188,30,188,29,113,31,193,31,187,31,65,31,246,31,53,31,53,30,34,31,128,31,94,31,115,31,42,31,105,31,105,30,45,31,73,31,73,30,212,31,135,31,158,31,73,31,165,31,209,31,253,31,7,31,239,31,209,31,209,30,209,29,91,31,171,31,116,31,75,31,8,31,56,31,96,31,66,31,213,31,88,31,17,31,27,31,27,30,54,31,54,30,217,31,217,30,97,31,248,31,248,30,195,31,15,31,252,31,198,31,246,31,39,31,239,31,60,31,251,31,251,30,169,31,169,30,191,31,18,31,16,31,249,31,249,30,110,31,24,31,76,31,151,31,250,31,152,31,139,31,204,31,204,30,141,31,165,31,90,31,90,30,90,29,65,31,108,31,190,31,198,31,7,31,232,31,3,31,205,31,249,31,7,31,183,31,253,31,21,31,235,31,70,31,100,31,167,31,151,31,151,30,36,31,96,31,177,31,17,31,75,31,75,30,242,31,78,31,209,31,180,31,61,31,250,31,140,31,16,31,73,31,3,31,221,31,205,31,205,30,50,31,67,31,13,31,99,31,2,31,2,30,2,29,204,31,204,30,255,31,255,30,88,31,88,31,88,30,200,31,235,31,166,31,109,31,35,31,125,31,116,31,53,31,190,31,55,31,47,31,181,31,104,31,16,31,45,31,234,31,225,31,159,31,222,31,113,31,98,31,111,31,111,30,182,31,2,31,53,31,53,30,53,29,251,31,205,31,110,31,112,31,162,31,12,31,237,31,203,31,251,31,251,30,14,31,61,31,40,31,90,31,107,31,107,30,82,31,94,31,248,31,241,31,59,31,29,31,35,31,204,31,188,31,188,30,188,29,104,31,24,31,186,31,186,30,61,31,245,31,88,31,83,31,197,31,152,31,152,30,26,31,184,31,184,30,50,31,84,31,84,30,255,31,162,31,158,31,96,31,38,31,187,31,5,31,12,31,144,31,111,31,111,30,111,29,60,31,187,31,222,31,117,31,43,31,49,31,227,31,188,31,188,30,131,31,60,31,121,31,245,31,237,31,173,31,160,31,139,31,139,30,214,31,217,31,230,31,232,31,17,31,17,30,216,31,216,30,50,31,219,31,47,31,7,31,105,31,198,31,17,31,200,31,191,31,14,31,14,30,112,31,9,31,192,31,240,31,39,31,35,31,114,31,114,30,114,29,115,31,115,30,150,31,138,31,59,31,236,31,226,31,102,31,34,31,178,31,127,31,157,31,70,31,137,31,137,30,241,31,84,31,51,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
