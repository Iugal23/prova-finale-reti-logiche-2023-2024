-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_384 is
end project_tb_384;

architecture project_tb_arch_384 of project_tb_384 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 861;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,212,0,236,0,19,0,67,0,152,0,0,0,240,0,98,0,19,0,88,0,60,0,0,0,0,0,0,0,159,0,248,0,187,0,175,0,150,0,102,0,112,0,216,0,102,0,208,0,193,0,24,0,132,0,0,0,54,0,187,0,0,0,101,0,248,0,0,0,31,0,237,0,101,0,0,0,0,0,66,0,184,0,35,0,64,0,0,0,0,0,0,0,189,0,251,0,0,0,167,0,0,0,36,0,96,0,172,0,71,0,144,0,32,0,0,0,111,0,143,0,0,0,100,0,53,0,138,0,154,0,125,0,177,0,223,0,0,0,77,0,74,0,0,0,153,0,0,0,44,0,0,0,236,0,26,0,0,0,163,0,78,0,0,0,112,0,129,0,154,0,84,0,149,0,17,0,15,0,88,0,230,0,76,0,88,0,83,0,48,0,83,0,0,0,6,0,173,0,55,0,251,0,217,0,190,0,155,0,206,0,227,0,180,0,0,0,0,0,95,0,8,0,184,0,165,0,134,0,197,0,0,0,54,0,145,0,134,0,42,0,86,0,229,0,135,0,232,0,0,0,0,0,0,0,46,0,0,0,248,0,3,0,168,0,166,0,151,0,47,0,2,0,147,0,0,0,100,0,103,0,0,0,0,0,205,0,102,0,117,0,109,0,27,0,158,0,0,0,1,0,146,0,0,0,98,0,59,0,39,0,0,0,138,0,117,0,215,0,0,0,105,0,201,0,99,0,222,0,169,0,204,0,16,0,0,0,0,0,123,0,189,0,54,0,104,0,184,0,196,0,158,0,250,0,92,0,119,0,0,0,126,0,189,0,235,0,245,0,3,0,0,0,51,0,185,0,160,0,0,0,103,0,75,0,214,0,64,0,131,0,235,0,0,0,142,0,161,0,90,0,134,0,216,0,245,0,178,0,16,0,0,0,13,0,209,0,8,0,212,0,114,0,182,0,155,0,155,0,154,0,142,0,241,0,0,0,186,0,0,0,94,0,174,0,128,0,240,0,53,0,45,0,60,0,0,0,141,0,206,0,203,0,173,0,103,0,35,0,82,0,236,0,0,0,0,0,0,0,0,0,0,0,228,0,205,0,178,0,155,0,110,0,0,0,0,0,204,0,0,0,169,0,168,0,68,0,237,0,183,0,249,0,30,0,0,0,0,0,165,0,181,0,128,0,0,0,18,0,126,0,208,0,191,0,67,0,0,0,0,0,184,0,208,0,31,0,0,0,0,0,166,0,168,0,35,0,210,0,80,0,236,0,81,0,222,0,190,0,45,0,196,0,0,0,108,0,80,0,45,0,35,0,152,0,111,0,0,0,43,0,189,0,44,0,137,0,0,0,156,0,28,0,67,0,0,0,158,0,0,0,14,0,126,0,0,0,194,0,0,0,219,0,0,0,22,0,0,0,0,0,220,0,58,0,131,0,25,0,0,0,6,0,61,0,0,0,188,0,208,0,127,0,112,0,172,0,104,0,79,0,0,0,205,0,0,0,99,0,232,0,65,0,0,0,27,0,65,0,133,0,202,0,182,0,0,0,54,0,91,0,84,0,106,0,0,0,0,0,246,0,6,0,202,0,134,0,0,0,97,0,198,0,0,0,0,0,139,0,231,0,126,0,0,0,246,0,93,0,98,0,0,0,0,0,238,0,220,0,92,0,120,0,0,0,183,0,0,0,0,0,179,0,237,0,0,0,186,0,114,0,63,0,0,0,22,0,131,0,39,0,220,0,0,0,20,0,233,0,5,0,169,0,36,0,212,0,96,0,59,0,5,0,189,0,200,0,0,0,212,0,247,0,0,0,11,0,71,0,125,0,79,0,126,0,123,0,201,0,0,0,85,0,93,0,219,0,0,0,66,0,0,0,210,0,155,0,0,0,40,0,125,0,217,0,255,0,230,0,0,0,0,0,0,0,55,0,113,0,38,0,115,0,192,0,33,0,0,0,81,0,11,0,216,0,75,0,53,0,0,0,44,0,57,0,0,0,137,0,0,0,199,0,236,0,78,0,42,0,8,0,76,0,155,0,0,0,64,0,38,0,0,0,219,0,139,0,110,0,236,0,11,0,29,0,235,0,0,0,17,0,54,0,196,0,187,0,133,0,80,0,62,0,206,0,33,0,202,0,248,0,69,0,0,0,0,0,0,0,51,0,228,0,59,0,71,0,166,0,139,0,98,0,68,0,246,0,181,0,96,0,0,0,122,0,56,0,26,0,192,0,149,0,134,0,123,0,66,0,58,0,1,0,0,0,134,0,21,0,0,0,251,0,187,0,244,0,126,0,21,0,61,0,0,0,0,0,154,0,217,0,0,0,253,0,68,0,214,0,55,0,32,0,0,0,0,0,215,0,185,0,165,0,0,0,0,0,0,0,0,0,0,0,21,0,207,0,29,0,70,0,0,0,162,0,57,0,52,0,0,0,233,0,0,0,75,0,173,0,65,0,10,0,0,0,0,0,25,0,108,0,73,0,0,0,44,0,92,0,246,0,0,0,0,0,53,0,157,0,0,0,39,0,24,0,103,0,241,0,0,0,0,0,0,0,0,0,0,0,42,0,29,0,139,0,7,0,0,0,53,0,0,0,82,0,171,0,11,0,53,0,0,0,75,0,173,0,0,0,24,0,164,0,10,0,35,0,239,0,37,0,39,0,0,0,174,0,245,0,79,0,150,0,119,0,28,0,222,0,169,0,23,0,0,0,0,0,43,0,164,0,212,0,53,0,222,0,141,0,9,0,121,0,107,0,129,0,35,0,50,0,153,0,0,0,242,0,99,0,0,0,46,0,0,0,141,0,0,0,129,0,60,0,238,0,94,0,104,0,89,0,244,0,59,0,175,0,56,0,61,0,0,0,78,0,14,0,240,0,18,0,0,0,0,0,0,0,58,0,135,0,206,0,0,0,189,0,151,0,228,0,0,0,0,0,27,0,239,0,44,0,7,0,48,0,201,0,181,0,116,0,192,0,255,0,187,0,110,0,177,0,0,0,0,0,14,0,98,0,222,0,0,0,105,0,1,0,0,0,216,0,127,0,225,0,0,0,48,0,104,0,231,0,0,0,34,0,0,0,238,0,64,0,93,0,99,0,221,0,0,0,132,0,130,0,66,0,135,0,0,0,65,0,252,0,231,0,54,0,201,0,80,0,166,0,166,0,56,0,31,0,128,0,151,0,12,0,25,0,110,0,138,0,0,0,70,0,137,0,0,0,93,0,150,0,75,0,241,0,25,0,198,0,211,0,140,0,178,0,175,0,24,0,90,0,0,0,69,0,0,0,254,0,22,0,148,0,0,0,106,0,6,0,53,0,2,0,0,0,153,0,134,0,47,0,253,0,0,0,250,0,60,0,0,0,161,0,140,0,0,0,83,0,77,0,0,0,98,0,179,0,183,0,0,0,50,0,6,0,0,0,0,0,0,0,250,0,151,0,66,0,226,0,0,0,229,0,236,0,75,0,22,0,0,0,0,0,57,0,0,0,145,0,221,0,28,0,0,0,219,0,26,0,58,0,239,0,70,0,141,0,37,0,0,0,0,0,0,0,0,0,0,0,100,0,44,0,47,0,172,0,178,0,154,0,0,0,83,0,244,0,112,0,146,0,61,0,80,0,34,0,127,0,0,0,158,0,135,0,55,0,0,0,6,0,0,0,75,0,0,0,107,0,185,0,7,0,152,0,195,0,0,0,47,0,164,0,233,0,37,0,125,0,106,0,0,0,0,0,61,0,225,0,168,0,33,0,133,0,186,0,224,0,48,0,26,0,128,0,0,0,0,0,223,0,107,0,61,0,194,0,30,0,0,0,196,0,148,0,0,0,7,0,176,0,128,0,48,0,0,0,17,0,228,0,254,0,181,0,158,0);
signal scenario_full  : scenario_type := (0,0,212,31,236,31,19,31,67,31,152,31,152,30,240,31,98,31,19,31,88,31,60,31,60,30,60,29,60,28,159,31,248,31,187,31,175,31,150,31,102,31,112,31,216,31,102,31,208,31,193,31,24,31,132,31,132,30,54,31,187,31,187,30,101,31,248,31,248,30,31,31,237,31,101,31,101,30,101,29,66,31,184,31,35,31,64,31,64,30,64,29,64,28,189,31,251,31,251,30,167,31,167,30,36,31,96,31,172,31,71,31,144,31,32,31,32,30,111,31,143,31,143,30,100,31,53,31,138,31,154,31,125,31,177,31,223,31,223,30,77,31,74,31,74,30,153,31,153,30,44,31,44,30,236,31,26,31,26,30,163,31,78,31,78,30,112,31,129,31,154,31,84,31,149,31,17,31,15,31,88,31,230,31,76,31,88,31,83,31,48,31,83,31,83,30,6,31,173,31,55,31,251,31,217,31,190,31,155,31,206,31,227,31,180,31,180,30,180,29,95,31,8,31,184,31,165,31,134,31,197,31,197,30,54,31,145,31,134,31,42,31,86,31,229,31,135,31,232,31,232,30,232,29,232,28,46,31,46,30,248,31,3,31,168,31,166,31,151,31,47,31,2,31,147,31,147,30,100,31,103,31,103,30,103,29,205,31,102,31,117,31,109,31,27,31,158,31,158,30,1,31,146,31,146,30,98,31,59,31,39,31,39,30,138,31,117,31,215,31,215,30,105,31,201,31,99,31,222,31,169,31,204,31,16,31,16,30,16,29,123,31,189,31,54,31,104,31,184,31,196,31,158,31,250,31,92,31,119,31,119,30,126,31,189,31,235,31,245,31,3,31,3,30,51,31,185,31,160,31,160,30,103,31,75,31,214,31,64,31,131,31,235,31,235,30,142,31,161,31,90,31,134,31,216,31,245,31,178,31,16,31,16,30,13,31,209,31,8,31,212,31,114,31,182,31,155,31,155,31,154,31,142,31,241,31,241,30,186,31,186,30,94,31,174,31,128,31,240,31,53,31,45,31,60,31,60,30,141,31,206,31,203,31,173,31,103,31,35,31,82,31,236,31,236,30,236,29,236,28,236,27,236,26,228,31,205,31,178,31,155,31,110,31,110,30,110,29,204,31,204,30,169,31,168,31,68,31,237,31,183,31,249,31,30,31,30,30,30,29,165,31,181,31,128,31,128,30,18,31,126,31,208,31,191,31,67,31,67,30,67,29,184,31,208,31,31,31,31,30,31,29,166,31,168,31,35,31,210,31,80,31,236,31,81,31,222,31,190,31,45,31,196,31,196,30,108,31,80,31,45,31,35,31,152,31,111,31,111,30,43,31,189,31,44,31,137,31,137,30,156,31,28,31,67,31,67,30,158,31,158,30,14,31,126,31,126,30,194,31,194,30,219,31,219,30,22,31,22,30,22,29,220,31,58,31,131,31,25,31,25,30,6,31,61,31,61,30,188,31,208,31,127,31,112,31,172,31,104,31,79,31,79,30,205,31,205,30,99,31,232,31,65,31,65,30,27,31,65,31,133,31,202,31,182,31,182,30,54,31,91,31,84,31,106,31,106,30,106,29,246,31,6,31,202,31,134,31,134,30,97,31,198,31,198,30,198,29,139,31,231,31,126,31,126,30,246,31,93,31,98,31,98,30,98,29,238,31,220,31,92,31,120,31,120,30,183,31,183,30,183,29,179,31,237,31,237,30,186,31,114,31,63,31,63,30,22,31,131,31,39,31,220,31,220,30,20,31,233,31,5,31,169,31,36,31,212,31,96,31,59,31,5,31,189,31,200,31,200,30,212,31,247,31,247,30,11,31,71,31,125,31,79,31,126,31,123,31,201,31,201,30,85,31,93,31,219,31,219,30,66,31,66,30,210,31,155,31,155,30,40,31,125,31,217,31,255,31,230,31,230,30,230,29,230,28,55,31,113,31,38,31,115,31,192,31,33,31,33,30,81,31,11,31,216,31,75,31,53,31,53,30,44,31,57,31,57,30,137,31,137,30,199,31,236,31,78,31,42,31,8,31,76,31,155,31,155,30,64,31,38,31,38,30,219,31,139,31,110,31,236,31,11,31,29,31,235,31,235,30,17,31,54,31,196,31,187,31,133,31,80,31,62,31,206,31,33,31,202,31,248,31,69,31,69,30,69,29,69,28,51,31,228,31,59,31,71,31,166,31,139,31,98,31,68,31,246,31,181,31,96,31,96,30,122,31,56,31,26,31,192,31,149,31,134,31,123,31,66,31,58,31,1,31,1,30,134,31,21,31,21,30,251,31,187,31,244,31,126,31,21,31,61,31,61,30,61,29,154,31,217,31,217,30,253,31,68,31,214,31,55,31,32,31,32,30,32,29,215,31,185,31,165,31,165,30,165,29,165,28,165,27,165,26,21,31,207,31,29,31,70,31,70,30,162,31,57,31,52,31,52,30,233,31,233,30,75,31,173,31,65,31,10,31,10,30,10,29,25,31,108,31,73,31,73,30,44,31,92,31,246,31,246,30,246,29,53,31,157,31,157,30,39,31,24,31,103,31,241,31,241,30,241,29,241,28,241,27,241,26,42,31,29,31,139,31,7,31,7,30,53,31,53,30,82,31,171,31,11,31,53,31,53,30,75,31,173,31,173,30,24,31,164,31,10,31,35,31,239,31,37,31,39,31,39,30,174,31,245,31,79,31,150,31,119,31,28,31,222,31,169,31,23,31,23,30,23,29,43,31,164,31,212,31,53,31,222,31,141,31,9,31,121,31,107,31,129,31,35,31,50,31,153,31,153,30,242,31,99,31,99,30,46,31,46,30,141,31,141,30,129,31,60,31,238,31,94,31,104,31,89,31,244,31,59,31,175,31,56,31,61,31,61,30,78,31,14,31,240,31,18,31,18,30,18,29,18,28,58,31,135,31,206,31,206,30,189,31,151,31,228,31,228,30,228,29,27,31,239,31,44,31,7,31,48,31,201,31,181,31,116,31,192,31,255,31,187,31,110,31,177,31,177,30,177,29,14,31,98,31,222,31,222,30,105,31,1,31,1,30,216,31,127,31,225,31,225,30,48,31,104,31,231,31,231,30,34,31,34,30,238,31,64,31,93,31,99,31,221,31,221,30,132,31,130,31,66,31,135,31,135,30,65,31,252,31,231,31,54,31,201,31,80,31,166,31,166,31,56,31,31,31,128,31,151,31,12,31,25,31,110,31,138,31,138,30,70,31,137,31,137,30,93,31,150,31,75,31,241,31,25,31,198,31,211,31,140,31,178,31,175,31,24,31,90,31,90,30,69,31,69,30,254,31,22,31,148,31,148,30,106,31,6,31,53,31,2,31,2,30,153,31,134,31,47,31,253,31,253,30,250,31,60,31,60,30,161,31,140,31,140,30,83,31,77,31,77,30,98,31,179,31,183,31,183,30,50,31,6,31,6,30,6,29,6,28,250,31,151,31,66,31,226,31,226,30,229,31,236,31,75,31,22,31,22,30,22,29,57,31,57,30,145,31,221,31,28,31,28,30,219,31,26,31,58,31,239,31,70,31,141,31,37,31,37,30,37,29,37,28,37,27,37,26,100,31,44,31,47,31,172,31,178,31,154,31,154,30,83,31,244,31,112,31,146,31,61,31,80,31,34,31,127,31,127,30,158,31,135,31,55,31,55,30,6,31,6,30,75,31,75,30,107,31,185,31,7,31,152,31,195,31,195,30,47,31,164,31,233,31,37,31,125,31,106,31,106,30,106,29,61,31,225,31,168,31,33,31,133,31,186,31,224,31,48,31,26,31,128,31,128,30,128,29,223,31,107,31,61,31,194,31,30,31,30,30,196,31,148,31,148,30,7,31,176,31,128,31,48,31,48,30,17,31,228,31,254,31,181,31,158,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
