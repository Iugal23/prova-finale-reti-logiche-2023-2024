-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_495 is
end project_tb_495;

architecture project_tb_arch_495 of project_tb_495 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 432;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (12,0,53,0,208,0,11,0,0,0,0,0,24,0,16,0,154,0,96,0,197,0,85,0,5,0,237,0,97,0,0,0,56,0,0,0,0,0,43,0,55,0,228,0,212,0,82,0,0,0,6,0,0,0,163,0,12,0,3,0,166,0,149,0,111,0,129,0,0,0,199,0,0,0,201,0,181,0,230,0,187,0,197,0,234,0,149,0,222,0,221,0,0,0,58,0,0,0,113,0,170,0,122,0,166,0,174,0,0,0,145,0,139,0,47,0,0,0,253,0,234,0,229,0,167,0,0,0,107,0,140,0,0,0,0,0,105,0,5,0,145,0,123,0,55,0,0,0,69,0,96,0,217,0,0,0,141,0,171,0,224,0,94,0,247,0,145,0,15,0,48,0,50,0,196,0,76,0,0,0,222,0,213,0,189,0,0,0,207,0,51,0,27,0,27,0,155,0,10,0,221,0,207,0,227,0,149,0,26,0,25,0,251,0,81,0,143,0,0,0,79,0,208,0,0,0,81,0,31,0,19,0,110,0,0,0,0,0,119,0,127,0,246,0,213,0,115,0,0,0,185,0,157,0,51,0,165,0,225,0,223,0,3,0,0,0,106,0,193,0,182,0,210,0,130,0,253,0,182,0,0,0,29,0,97,0,163,0,106,0,98,0,0,0,176,0,94,0,52,0,135,0,156,0,38,0,5,0,163,0,34,0,151,0,115,0,185,0,185,0,5,0,23,0,153,0,215,0,181,0,52,0,105,0,138,0,201,0,0,0,115,0,0,0,45,0,0,0,0,0,70,0,52,0,0,0,253,0,36,0,128,0,43,0,38,0,240,0,0,0,31,0,0,0,182,0,252,0,0,0,64,0,112,0,169,0,0,0,20,0,214,0,237,0,239,0,0,0,198,0,0,0,237,0,86,0,67,0,62,0,131,0,151,0,127,0,0,0,212,0,232,0,0,0,212,0,0,0,215,0,171,0,229,0,0,0,43,0,220,0,3,0,172,0,0,0,158,0,185,0,216,0,26,0,0,0,7,0,156,0,127,0,85,0,227,0,0,0,66,0,45,0,255,0,0,0,240,0,0,0,178,0,12,0,33,0,124,0,2,0,189,0,193,0,238,0,214,0,57,0,0,0,23,0,45,0,169,0,235,0,0,0,8,0,161,0,156,0,208,0,157,0,17,0,24,0,196,0,197,0,186,0,151,0,184,0,127,0,228,0,251,0,89,0,207,0,12,0,0,0,197,0,63,0,39,0,142,0,0,0,0,0,32,0,49,0,0,0,76,0,5,0,1,0,0,0,27,0,175,0,78,0,0,0,86,0,6,0,207,0,36,0,0,0,60,0,18,0,0,0,195,0,73,0,1,0,139,0,86,0,129,0,0,0,101,0,17,0,0,0,0,0,143,0,216,0,5,0,54,0,209,0,106,0,123,0,151,0,240,0,147,0,4,0,86,0,211,0,70,0,210,0,118,0,7,0,78,0,0,0,178,0,239,0,143,0,60,0,115,0,80,0,193,0,113,0,0,0,126,0,0,0,0,0,156,0,152,0,172,0,59,0,98,0,155,0,139,0,65,0,66,0,40,0,94,0,240,0,0,0,56,0,0,0,63,0,224,0,254,0,44,0,241,0,0,0,227,0,0,0,106,0,98,0,243,0,36,0,26,0,0,0,18,0,49,0,142,0,230,0,36,0,26,0,84,0,57,0,233,0,51,0,18,0,0,0,38,0,150,0,27,0,177,0,111,0,176,0,0,0,158,0,56,0,102,0,47,0,249,0,0,0,24,0,141,0,0,0,89,0,0,0,34,0,170,0,156,0,249,0,112,0,185,0,34,0,69,0,23,0,0,0,103,0,0,0,151,0,186,0,38,0,200,0,195,0,115,0,0,0,194,0,19,0,0,0,64,0,99,0,247,0,0,0,1,0,249,0,76,0,152,0,221,0);
signal scenario_full  : scenario_type := (12,31,53,31,208,31,11,31,11,30,11,29,24,31,16,31,154,31,96,31,197,31,85,31,5,31,237,31,97,31,97,30,56,31,56,30,56,29,43,31,55,31,228,31,212,31,82,31,82,30,6,31,6,30,163,31,12,31,3,31,166,31,149,31,111,31,129,31,129,30,199,31,199,30,201,31,181,31,230,31,187,31,197,31,234,31,149,31,222,31,221,31,221,30,58,31,58,30,113,31,170,31,122,31,166,31,174,31,174,30,145,31,139,31,47,31,47,30,253,31,234,31,229,31,167,31,167,30,107,31,140,31,140,30,140,29,105,31,5,31,145,31,123,31,55,31,55,30,69,31,96,31,217,31,217,30,141,31,171,31,224,31,94,31,247,31,145,31,15,31,48,31,50,31,196,31,76,31,76,30,222,31,213,31,189,31,189,30,207,31,51,31,27,31,27,31,155,31,10,31,221,31,207,31,227,31,149,31,26,31,25,31,251,31,81,31,143,31,143,30,79,31,208,31,208,30,81,31,31,31,19,31,110,31,110,30,110,29,119,31,127,31,246,31,213,31,115,31,115,30,185,31,157,31,51,31,165,31,225,31,223,31,3,31,3,30,106,31,193,31,182,31,210,31,130,31,253,31,182,31,182,30,29,31,97,31,163,31,106,31,98,31,98,30,176,31,94,31,52,31,135,31,156,31,38,31,5,31,163,31,34,31,151,31,115,31,185,31,185,31,5,31,23,31,153,31,215,31,181,31,52,31,105,31,138,31,201,31,201,30,115,31,115,30,45,31,45,30,45,29,70,31,52,31,52,30,253,31,36,31,128,31,43,31,38,31,240,31,240,30,31,31,31,30,182,31,252,31,252,30,64,31,112,31,169,31,169,30,20,31,214,31,237,31,239,31,239,30,198,31,198,30,237,31,86,31,67,31,62,31,131,31,151,31,127,31,127,30,212,31,232,31,232,30,212,31,212,30,215,31,171,31,229,31,229,30,43,31,220,31,3,31,172,31,172,30,158,31,185,31,216,31,26,31,26,30,7,31,156,31,127,31,85,31,227,31,227,30,66,31,45,31,255,31,255,30,240,31,240,30,178,31,12,31,33,31,124,31,2,31,189,31,193,31,238,31,214,31,57,31,57,30,23,31,45,31,169,31,235,31,235,30,8,31,161,31,156,31,208,31,157,31,17,31,24,31,196,31,197,31,186,31,151,31,184,31,127,31,228,31,251,31,89,31,207,31,12,31,12,30,197,31,63,31,39,31,142,31,142,30,142,29,32,31,49,31,49,30,76,31,5,31,1,31,1,30,27,31,175,31,78,31,78,30,86,31,6,31,207,31,36,31,36,30,60,31,18,31,18,30,195,31,73,31,1,31,139,31,86,31,129,31,129,30,101,31,17,31,17,30,17,29,143,31,216,31,5,31,54,31,209,31,106,31,123,31,151,31,240,31,147,31,4,31,86,31,211,31,70,31,210,31,118,31,7,31,78,31,78,30,178,31,239,31,143,31,60,31,115,31,80,31,193,31,113,31,113,30,126,31,126,30,126,29,156,31,152,31,172,31,59,31,98,31,155,31,139,31,65,31,66,31,40,31,94,31,240,31,240,30,56,31,56,30,63,31,224,31,254,31,44,31,241,31,241,30,227,31,227,30,106,31,98,31,243,31,36,31,26,31,26,30,18,31,49,31,142,31,230,31,36,31,26,31,84,31,57,31,233,31,51,31,18,31,18,30,38,31,150,31,27,31,177,31,111,31,176,31,176,30,158,31,56,31,102,31,47,31,249,31,249,30,24,31,141,31,141,30,89,31,89,30,34,31,170,31,156,31,249,31,112,31,185,31,34,31,69,31,23,31,23,30,103,31,103,30,151,31,186,31,38,31,200,31,195,31,115,31,115,30,194,31,19,31,19,30,64,31,99,31,247,31,247,30,1,31,249,31,76,31,152,31,221,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
