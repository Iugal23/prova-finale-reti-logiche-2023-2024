-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1006;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (53,0,0,0,0,0,0,0,102,0,187,0,27,0,68,0,159,0,93,0,200,0,177,0,0,0,62,0,34,0,198,0,94,0,107,0,63,0,81,0,30,0,31,0,9,0,0,0,166,0,193,0,31,0,134,0,132,0,0,0,65,0,240,0,78,0,188,0,0,0,242,0,39,0,114,0,19,0,15,0,136,0,5,0,220,0,0,0,43,0,159,0,128,0,0,0,113,0,0,0,136,0,0,0,184,0,5,0,166,0,225,0,131,0,99,0,144,0,215,0,39,0,11,0,62,0,222,0,196,0,64,0,131,0,219,0,0,0,0,0,207,0,105,0,15,0,219,0,186,0,205,0,87,0,152,0,14,0,17,0,40,0,5,0,211,0,68,0,0,0,133,0,183,0,0,0,192,0,219,0,130,0,80,0,165,0,150,0,85,0,159,0,0,0,0,0,77,0,1,0,79,0,214,0,244,0,69,0,56,0,163,0,0,0,190,0,11,0,0,0,0,0,172,0,50,0,244,0,183,0,0,0,122,0,232,0,0,0,240,0,0,0,117,0,0,0,141,0,218,0,148,0,85,0,137,0,168,0,233,0,43,0,43,0,170,0,142,0,123,0,229,0,122,0,0,0,153,0,211,0,134,0,0,0,179,0,0,0,0,0,0,0,96,0,0,0,130,0,142,0,136,0,149,0,25,0,93,0,239,0,111,0,232,0,145,0,75,0,86,0,236,0,172,0,150,0,169,0,11,0,0,0,80,0,254,0,132,0,241,0,32,0,147,0,154,0,0,0,0,0,26,0,83,0,39,0,0,0,238,0,40,0,0,0,0,0,78,0,187,0,133,0,89,0,92,0,144,0,195,0,57,0,189,0,0,0,0,0,209,0,44,0,0,0,139,0,103,0,0,0,215,0,0,0,0,0,68,0,210,0,117,0,122,0,0,0,227,0,53,0,150,0,0,0,159,0,0,0,231,0,194,0,109,0,69,0,223,0,50,0,103,0,163,0,216,0,106,0,203,0,0,0,21,0,243,0,214,0,38,0,63,0,131,0,0,0,0,0,56,0,1,0,0,0,200,0,18,0,152,0,132,0,0,0,0,0,0,0,33,0,0,0,169,0,233,0,188,0,19,0,123,0,0,0,25,0,0,0,247,0,106,0,138,0,0,0,0,0,168,0,41,0,0,0,0,0,149,0,128,0,57,0,156,0,55,0,15,0,249,0,150,0,0,0,187,0,224,0,209,0,191,0,192,0,0,0,178,0,86,0,123,0,0,0,109,0,211,0,70,0,216,0,27,0,235,0,254,0,163,0,6,0,213,0,0,0,150,0,74,0,111,0,245,0,97,0,114,0,66,0,187,0,171,0,230,0,74,0,85,0,0,0,219,0,142,0,62,0,178,0,9,0,94,0,157,0,178,0,108,0,202,0,53,0,245,0,197,0,49,0,0,0,180,0,69,0,70,0,228,0,222,0,88,0,11,0,101,0,1,0,85,0,68,0,0,0,214,0,44,0,0,0,19,0,119,0,0,0,213,0,133,0,121,0,214,0,33,0,244,0,226,0,191,0,190,0,40,0,168,0,0,0,221,0,178,0,98,0,253,0,21,0,99,0,77,0,0,0,0,0,133,0,126,0,0,0,0,0,0,0,203,0,177,0,0,0,216,0,172,0,210,0,0,0,170,0,207,0,77,0,171,0,242,0,169,0,163,0,166,0,0,0,249,0,86,0,145,0,0,0,150,0,253,0,103,0,180,0,52,0,0,0,0,0,0,0,219,0,0,0,191,0,0,0,92,0,206,0,101,0,105,0,155,0,37,0,106,0,159,0,208,0,36,0,125,0,184,0,230,0,116,0,216,0,154,0,0,0,255,0,127,0,18,0,0,0,44,0,219,0,0,0,221,0,13,0,235,0,254,0,13,0,142,0,224,0,18,0,141,0,226,0,194,0,109,0,59,0,96,0,126,0,227,0,209,0,240,0,157,0,0,0,215,0,146,0,88,0,97,0,135,0,63,0,0,0,177,0,225,0,0,0,0,0,0,0,152,0,134,0,143,0,0,0,135,0,245,0,242,0,108,0,154,0,53,0,0,0,169,0,241,0,0,0,7,0,0,0,8,0,232,0,0,0,10,0,0,0,215,0,0,0,126,0,24,0,57,0,211,0,32,0,0,0,0,0,79,0,228,0,128,0,245,0,158,0,137,0,61,0,74,0,0,0,2,0,72,0,251,0,108,0,114,0,0,0,205,0,0,0,0,0,87,0,209,0,186,0,0,0,14,0,17,0,72,0,45,0,63,0,63,0,244,0,228,0,0,0,113,0,166,0,225,0,149,0,0,0,14,0,188,0,187,0,118,0,49,0,0,0,216,0,68,0,85,0,0,0,97,0,222,0,31,0,47,0,251,0,137,0,0,0,0,0,115,0,0,0,158,0,53,0,133,0,162,0,86,0,119,0,158,0,20,0,252,0,184,0,0,0,156,0,101,0,12,0,69,0,152,0,210,0,23,0,0,0,28,0,182,0,0,0,33,0,130,0,74,0,44,0,228,0,243,0,200,0,74,0,32,0,0,0,74,0,106,0,106,0,220,0,0,0,145,0,105,0,52,0,172,0,0,0,124,0,83,0,166,0,188,0,157,0,75,0,0,0,0,0,71,0,22,0,87,0,38,0,58,0,124,0,0,0,82,0,195,0,64,0,18,0,0,0,197,0,83,0,104,0,193,0,118,0,68,0,3,0,158,0,0,0,242,0,134,0,150,0,135,0,0,0,206,0,0,0,243,0,253,0,3,0,11,0,119,0,9,0,204,0,255,0,197,0,139,0,0,0,207,0,218,0,0,0,246,0,0,0,249,0,255,0,105,0,0,0,46,0,172,0,0,0,0,0,41,0,184,0,0,0,166,0,203,0,101,0,238,0,117,0,216,0,0,0,0,0,52,0,58,0,65,0,32,0,200,0,72,0,50,0,244,0,145,0,202,0,0,0,69,0,67,0,242,0,186,0,118,0,0,0,138,0,27,0,199,0,144,0,180,0,0,0,5,0,7,0,0,0,7,0,0,0,225,0,0,0,0,0,167,0,139,0,0,0,113,0,91,0,0,0,152,0,77,0,144,0,51,0,76,0,0,0,84,0,151,0,14,0,0,0,135,0,136,0,211,0,82,0,243,0,183,0,127,0,62,0,36,0,70,0,197,0,140,0,137,0,149,0,235,0,173,0,0,0,43,0,30,0,57,0,20,0,0,0,18,0,0,0,209,0,31,0,0,0,36,0,20,0,127,0,0,0,107,0,31,0,158,0,0,0,182,0,6,0,92,0,152,0,138,0,0,0,10,0,59,0,155,0,0,0,0,0,132,0,119,0,79,0,244,0,144,0,3,0,0,0,244,0,99,0,0,0,77,0,136,0,253,0,161,0,162,0,0,0,53,0,150,0,255,0,0,0,0,0,55,0,4,0,12,0,0,0,160,0,125,0,150,0,0,0,251,0,0,0,27,0,64,0,252,0,87,0,134,0,113,0,215,0,47,0,127,0,118,0,0,0,225,0,75,0,184,0,95,0,146,0,195,0,193,0,135,0,28,0,168,0,143,0,15,0,42,0,49,0,80,0,136,0,38,0,116,0,0,0,0,0,193,0,0,0,85,0,0,0,0,0,70,0,0,0,0,0,132,0,95,0,0,0,27,0,101,0,206,0,197,0,0,0,99,0,184,0,168,0,210,0,214,0,131,0,0,0,93,0,6,0,130,0,100,0,227,0,0,0,189,0,255,0,8,0,0,0,236,0,191,0,75,0,15,0,153,0,0,0,0,0,0,0,167,0,174,0,182,0,48,0,113,0,158,0,34,0,78,0,78,0,174,0,0,0,191,0,86,0,0,0,238,0,122,0,57,0,133,0,49,0,121,0,1,0,0,0,92,0,137,0,50,0,4,0,98,0,22,0,0,0,0,0,0,0,117,0,236,0,155,0,0,0,99,0,136,0,0,0,15,0,17,0,88,0,0,0,50,0,0,0,149,0,100,0,165,0,0,0,204,0,89,0,0,0,128,0,158,0,246,0,191,0,226,0,148,0,77,0,227,0,17,0,0,0,19,0,162,0,119,0,128,0,2,0,102,0,151,0,222,0,21,0,60,0,170,0,0,0,94,0,84,0,248,0,94,0,0,0,199,0,133,0,0,0,218,0,129,0,0,0,0,0,80,0,39,0,160,0,116,0,8,0,32,0,30,0,20,0,30,0,159,0,30,0,0,0,195,0,225,0,222,0,250,0,179,0,28,0,222,0,22,0,241,0,0,0,151,0,57,0,0,0,83,0,132,0,213,0,6,0,231,0,131,0,16,0,123,0,15,0,185,0,213,0,0,0,128,0,0,0,156,0,148,0,174,0,172,0,145,0,247,0,12,0,169,0,207,0,0,0,58,0,0,0,108,0,2,0,235,0,154,0,78,0,0,0,113,0,1,0,0,0,108,0,244,0,210,0,242,0,0,0,0,0,31,0,238,0,208,0,244,0,185,0,53,0,183,0);
signal scenario_full  : scenario_type := (53,31,53,30,53,29,53,28,102,31,187,31,27,31,68,31,159,31,93,31,200,31,177,31,177,30,62,31,34,31,198,31,94,31,107,31,63,31,81,31,30,31,31,31,9,31,9,30,166,31,193,31,31,31,134,31,132,31,132,30,65,31,240,31,78,31,188,31,188,30,242,31,39,31,114,31,19,31,15,31,136,31,5,31,220,31,220,30,43,31,159,31,128,31,128,30,113,31,113,30,136,31,136,30,184,31,5,31,166,31,225,31,131,31,99,31,144,31,215,31,39,31,11,31,62,31,222,31,196,31,64,31,131,31,219,31,219,30,219,29,207,31,105,31,15,31,219,31,186,31,205,31,87,31,152,31,14,31,17,31,40,31,5,31,211,31,68,31,68,30,133,31,183,31,183,30,192,31,219,31,130,31,80,31,165,31,150,31,85,31,159,31,159,30,159,29,77,31,1,31,79,31,214,31,244,31,69,31,56,31,163,31,163,30,190,31,11,31,11,30,11,29,172,31,50,31,244,31,183,31,183,30,122,31,232,31,232,30,240,31,240,30,117,31,117,30,141,31,218,31,148,31,85,31,137,31,168,31,233,31,43,31,43,31,170,31,142,31,123,31,229,31,122,31,122,30,153,31,211,31,134,31,134,30,179,31,179,30,179,29,179,28,96,31,96,30,130,31,142,31,136,31,149,31,25,31,93,31,239,31,111,31,232,31,145,31,75,31,86,31,236,31,172,31,150,31,169,31,11,31,11,30,80,31,254,31,132,31,241,31,32,31,147,31,154,31,154,30,154,29,26,31,83,31,39,31,39,30,238,31,40,31,40,30,40,29,78,31,187,31,133,31,89,31,92,31,144,31,195,31,57,31,189,31,189,30,189,29,209,31,44,31,44,30,139,31,103,31,103,30,215,31,215,30,215,29,68,31,210,31,117,31,122,31,122,30,227,31,53,31,150,31,150,30,159,31,159,30,231,31,194,31,109,31,69,31,223,31,50,31,103,31,163,31,216,31,106,31,203,31,203,30,21,31,243,31,214,31,38,31,63,31,131,31,131,30,131,29,56,31,1,31,1,30,200,31,18,31,152,31,132,31,132,30,132,29,132,28,33,31,33,30,169,31,233,31,188,31,19,31,123,31,123,30,25,31,25,30,247,31,106,31,138,31,138,30,138,29,168,31,41,31,41,30,41,29,149,31,128,31,57,31,156,31,55,31,15,31,249,31,150,31,150,30,187,31,224,31,209,31,191,31,192,31,192,30,178,31,86,31,123,31,123,30,109,31,211,31,70,31,216,31,27,31,235,31,254,31,163,31,6,31,213,31,213,30,150,31,74,31,111,31,245,31,97,31,114,31,66,31,187,31,171,31,230,31,74,31,85,31,85,30,219,31,142,31,62,31,178,31,9,31,94,31,157,31,178,31,108,31,202,31,53,31,245,31,197,31,49,31,49,30,180,31,69,31,70,31,228,31,222,31,88,31,11,31,101,31,1,31,85,31,68,31,68,30,214,31,44,31,44,30,19,31,119,31,119,30,213,31,133,31,121,31,214,31,33,31,244,31,226,31,191,31,190,31,40,31,168,31,168,30,221,31,178,31,98,31,253,31,21,31,99,31,77,31,77,30,77,29,133,31,126,31,126,30,126,29,126,28,203,31,177,31,177,30,216,31,172,31,210,31,210,30,170,31,207,31,77,31,171,31,242,31,169,31,163,31,166,31,166,30,249,31,86,31,145,31,145,30,150,31,253,31,103,31,180,31,52,31,52,30,52,29,52,28,219,31,219,30,191,31,191,30,92,31,206,31,101,31,105,31,155,31,37,31,106,31,159,31,208,31,36,31,125,31,184,31,230,31,116,31,216,31,154,31,154,30,255,31,127,31,18,31,18,30,44,31,219,31,219,30,221,31,13,31,235,31,254,31,13,31,142,31,224,31,18,31,141,31,226,31,194,31,109,31,59,31,96,31,126,31,227,31,209,31,240,31,157,31,157,30,215,31,146,31,88,31,97,31,135,31,63,31,63,30,177,31,225,31,225,30,225,29,225,28,152,31,134,31,143,31,143,30,135,31,245,31,242,31,108,31,154,31,53,31,53,30,169,31,241,31,241,30,7,31,7,30,8,31,232,31,232,30,10,31,10,30,215,31,215,30,126,31,24,31,57,31,211,31,32,31,32,30,32,29,79,31,228,31,128,31,245,31,158,31,137,31,61,31,74,31,74,30,2,31,72,31,251,31,108,31,114,31,114,30,205,31,205,30,205,29,87,31,209,31,186,31,186,30,14,31,17,31,72,31,45,31,63,31,63,31,244,31,228,31,228,30,113,31,166,31,225,31,149,31,149,30,14,31,188,31,187,31,118,31,49,31,49,30,216,31,68,31,85,31,85,30,97,31,222,31,31,31,47,31,251,31,137,31,137,30,137,29,115,31,115,30,158,31,53,31,133,31,162,31,86,31,119,31,158,31,20,31,252,31,184,31,184,30,156,31,101,31,12,31,69,31,152,31,210,31,23,31,23,30,28,31,182,31,182,30,33,31,130,31,74,31,44,31,228,31,243,31,200,31,74,31,32,31,32,30,74,31,106,31,106,31,220,31,220,30,145,31,105,31,52,31,172,31,172,30,124,31,83,31,166,31,188,31,157,31,75,31,75,30,75,29,71,31,22,31,87,31,38,31,58,31,124,31,124,30,82,31,195,31,64,31,18,31,18,30,197,31,83,31,104,31,193,31,118,31,68,31,3,31,158,31,158,30,242,31,134,31,150,31,135,31,135,30,206,31,206,30,243,31,253,31,3,31,11,31,119,31,9,31,204,31,255,31,197,31,139,31,139,30,207,31,218,31,218,30,246,31,246,30,249,31,255,31,105,31,105,30,46,31,172,31,172,30,172,29,41,31,184,31,184,30,166,31,203,31,101,31,238,31,117,31,216,31,216,30,216,29,52,31,58,31,65,31,32,31,200,31,72,31,50,31,244,31,145,31,202,31,202,30,69,31,67,31,242,31,186,31,118,31,118,30,138,31,27,31,199,31,144,31,180,31,180,30,5,31,7,31,7,30,7,31,7,30,225,31,225,30,225,29,167,31,139,31,139,30,113,31,91,31,91,30,152,31,77,31,144,31,51,31,76,31,76,30,84,31,151,31,14,31,14,30,135,31,136,31,211,31,82,31,243,31,183,31,127,31,62,31,36,31,70,31,197,31,140,31,137,31,149,31,235,31,173,31,173,30,43,31,30,31,57,31,20,31,20,30,18,31,18,30,209,31,31,31,31,30,36,31,20,31,127,31,127,30,107,31,31,31,158,31,158,30,182,31,6,31,92,31,152,31,138,31,138,30,10,31,59,31,155,31,155,30,155,29,132,31,119,31,79,31,244,31,144,31,3,31,3,30,244,31,99,31,99,30,77,31,136,31,253,31,161,31,162,31,162,30,53,31,150,31,255,31,255,30,255,29,55,31,4,31,12,31,12,30,160,31,125,31,150,31,150,30,251,31,251,30,27,31,64,31,252,31,87,31,134,31,113,31,215,31,47,31,127,31,118,31,118,30,225,31,75,31,184,31,95,31,146,31,195,31,193,31,135,31,28,31,168,31,143,31,15,31,42,31,49,31,80,31,136,31,38,31,116,31,116,30,116,29,193,31,193,30,85,31,85,30,85,29,70,31,70,30,70,29,132,31,95,31,95,30,27,31,101,31,206,31,197,31,197,30,99,31,184,31,168,31,210,31,214,31,131,31,131,30,93,31,6,31,130,31,100,31,227,31,227,30,189,31,255,31,8,31,8,30,236,31,191,31,75,31,15,31,153,31,153,30,153,29,153,28,167,31,174,31,182,31,48,31,113,31,158,31,34,31,78,31,78,31,174,31,174,30,191,31,86,31,86,30,238,31,122,31,57,31,133,31,49,31,121,31,1,31,1,30,92,31,137,31,50,31,4,31,98,31,22,31,22,30,22,29,22,28,117,31,236,31,155,31,155,30,99,31,136,31,136,30,15,31,17,31,88,31,88,30,50,31,50,30,149,31,100,31,165,31,165,30,204,31,89,31,89,30,128,31,158,31,246,31,191,31,226,31,148,31,77,31,227,31,17,31,17,30,19,31,162,31,119,31,128,31,2,31,102,31,151,31,222,31,21,31,60,31,170,31,170,30,94,31,84,31,248,31,94,31,94,30,199,31,133,31,133,30,218,31,129,31,129,30,129,29,80,31,39,31,160,31,116,31,8,31,32,31,30,31,20,31,30,31,159,31,30,31,30,30,195,31,225,31,222,31,250,31,179,31,28,31,222,31,22,31,241,31,241,30,151,31,57,31,57,30,83,31,132,31,213,31,6,31,231,31,131,31,16,31,123,31,15,31,185,31,213,31,213,30,128,31,128,30,156,31,148,31,174,31,172,31,145,31,247,31,12,31,169,31,207,31,207,30,58,31,58,30,108,31,2,31,235,31,154,31,78,31,78,30,113,31,1,31,1,30,108,31,244,31,210,31,242,31,242,30,242,29,31,31,238,31,208,31,244,31,185,31,53,31,183,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
