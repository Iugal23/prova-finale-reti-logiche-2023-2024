-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_543 is
end project_tb_543;

architecture project_tb_arch_543 of project_tb_543 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 951;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (140,0,11,0,47,0,31,0,33,0,194,0,180,0,114,0,115,0,33,0,11,0,63,0,42,0,0,0,253,0,180,0,182,0,43,0,241,0,248,0,87,0,49,0,29,0,33,0,171,0,79,0,107,0,34,0,32,0,0,0,245,0,192,0,216,0,51,0,51,0,16,0,72,0,64,0,0,0,178,0,237,0,26,0,127,0,207,0,14,0,160,0,0,0,137,0,152,0,13,0,125,0,243,0,0,0,206,0,34,0,137,0,107,0,0,0,196,0,212,0,137,0,227,0,213,0,0,0,19,0,113,0,204,0,117,0,80,0,229,0,9,0,76,0,23,0,0,0,7,0,0,0,75,0,128,0,0,0,162,0,39,0,200,0,163,0,0,0,0,0,0,0,107,0,30,0,75,0,224,0,89,0,118,0,220,0,102,0,248,0,157,0,88,0,115,0,167,0,96,0,194,0,177,0,23,0,137,0,72,0,20,0,89,0,83,0,221,0,11,0,0,0,48,0,55,0,45,0,235,0,246,0,0,0,23,0,228,0,64,0,0,0,45,0,125,0,186,0,58,0,68,0,213,0,0,0,187,0,126,0,94,0,135,0,74,0,140,0,0,0,99,0,4,0,180,0,50,0,72,0,13,0,214,0,243,0,0,0,0,0,227,0,57,0,86,0,61,0,36,0,3,0,29,0,236,0,93,0,54,0,0,0,238,0,72,0,252,0,240,0,252,0,60,0,0,0,141,0,247,0,107,0,67,0,28,0,157,0,46,0,86,0,78,0,175,0,51,0,194,0,0,0,76,0,78,0,44,0,94,0,198,0,165,0,0,0,218,0,0,0,0,0,73,0,182,0,0,0,83,0,0,0,56,0,0,0,0,0,0,0,34,0,61,0,175,0,189,0,180,0,27,0,23,0,35,0,83,0,9,0,134,0,231,0,219,0,19,0,83,0,116,0,59,0,202,0,0,0,71,0,57,0,3,0,44,0,185,0,142,0,192,0,8,0,0,0,30,0,12,0,156,0,69,0,140,0,11,0,0,0,39,0,121,0,250,0,0,0,84,0,41,0,94,0,65,0,144,0,49,0,152,0,113,0,42,0,49,0,8,0,198,0,149,0,7,0,119,0,0,0,0,0,254,0,38,0,34,0,1,0,156,0,216,0,0,0,65,0,0,0,67,0,103,0,195,0,138,0,157,0,48,0,81,0,0,0,154,0,251,0,214,0,150,0,119,0,231,0,12,0,151,0,34,0,185,0,0,0,0,0,60,0,0,0,70,0,86,0,155,0,71,0,226,0,218,0,13,0,0,0,88,0,8,0,196,0,58,0,0,0,131,0,87,0,0,0,107,0,0,0,201,0,125,0,169,0,210,0,194,0,204,0,105,0,46,0,241,0,219,0,187,0,117,0,23,0,0,0,0,0,46,0,168,0,50,0,142,0,0,0,88,0,149,0,46,0,39,0,83,0,34,0,176,0,243,0,230,0,56,0,0,0,31,0,178,0,138,0,38,0,0,0,103,0,0,0,159,0,243,0,242,0,206,0,183,0,42,0,19,0,0,0,199,0,37,0,100,0,58,0,137,0,0,0,164,0,193,0,199,0,10,0,168,0,147,0,47,0,192,0,96,0,0,0,110,0,142,0,103,0,195,0,0,0,248,0,40,0,196,0,0,0,0,0,0,0,0,0,108,0,179,0,87,0,199,0,220,0,161,0,89,0,82,0,193,0,213,0,49,0,127,0,127,0,59,0,113,0,18,0,247,0,0,0,126,0,16,0,179,0,12,0,159,0,13,0,249,0,231,0,53,0,252,0,180,0,173,0,0,0,63,0,50,0,96,0,77,0,59,0,13,0,202,0,251,0,0,0,0,0,16,0,236,0,43,0,10,0,185,0,65,0,80,0,217,0,195,0,0,0,20,0,210,0,0,0,194,0,0,0,221,0,0,0,43,0,173,0,152,0,179,0,42,0,39,0,78,0,136,0,0,0,227,0,134,0,123,0,196,0,56,0,188,0,188,0,153,0,0,0,138,0,0,0,0,0,72,0,147,0,28,0,14,0,166,0,164,0,214,0,7,0,231,0,117,0,0,0,59,0,27,0,32,0,217,0,91,0,189,0,0,0,3,0,59,0,0,0,0,0,54,0,134,0,0,0,12,0,18,0,98,0,0,0,0,0,0,0,125,0,197,0,93,0,196,0,109,0,135,0,38,0,91,0,55,0,175,0,236,0,204,0,136,0,11,0,251,0,165,0,203,0,218,0,161,0,230,0,139,0,122,0,150,0,0,0,46,0,121,0,12,0,176,0,0,0,139,0,188,0,210,0,236,0,13,0,0,0,177,0,248,0,4,0,128,0,0,0,101,0,0,0,75,0,0,0,233,0,135,0,210,0,31,0,246,0,164,0,92,0,0,0,0,0,57,0,78,0,34,0,0,0,151,0,0,0,0,0,126,0,69,0,92,0,154,0,224,0,89,0,94,0,169,0,0,0,143,0,0,0,139,0,138,0,212,0,38,0,142,0,175,0,0,0,0,0,72,0,112,0,160,0,0,0,12,0,123,0,193,0,189,0,0,0,202,0,115,0,38,0,13,0,216,0,166,0,18,0,43,0,0,0,1,0,0,0,46,0,208,0,209,0,181,0,0,0,237,0,236,0,233,0,0,0,0,0,78,0,0,0,38,0,0,0,169,0,154,0,0,0,210,0,60,0,109,0,111,0,58,0,0,0,249,0,12,0,214,0,214,0,113,0,0,0,99,0,243,0,50,0,47,0,47,0,0,0,187,0,253,0,213,0,174,0,17,0,143,0,0,0,142,0,0,0,144,0,81,0,26,0,78,0,0,0,0,0,30,0,45,0,140,0,215,0,55,0,11,0,58,0,49,0,28,0,80,0,0,0,134,0,189,0,188,0,52,0,96,0,57,0,103,0,35,0,243,0,60,0,1,0,178,0,85,0,20,0,0,0,198,0,139,0,0,0,51,0,233,0,53,0,108,0,129,0,0,0,91,0,201,0,145,0,131,0,0,0,169,0,171,0,209,0,7,0,141,0,230,0,0,0,0,0,125,0,249,0,190,0,121,0,52,0,156,0,176,0,0,0,5,0,0,0,33,0,0,0,82,0,231,0,203,0,58,0,86,0,250,0,241,0,42,0,60,0,0,0,0,0,55,0,172,0,162,0,62,0,195,0,163,0,0,0,95,0,161,0,251,0,238,0,200,0,102,0,0,0,251,0,115,0,254,0,102,0,22,0,53,0,109,0,165,0,189,0,151,0,8,0,235,0,0,0,144,0,0,0,145,0,246,0,40,0,69,0,47,0,88,0,117,0,0,0,214,0,0,0,0,0,189,0,87,0,0,0,61,0,200,0,0,0,237,0,65,0,145,0,205,0,87,0,134,0,0,0,8,0,0,0,78,0,73,0,17,0,106,0,41,0,0,0,94,0,131,0,0,0,69,0,114,0,146,0,42,0,0,0,114,0,43,0,0,0,134,0,252,0,212,0,32,0,69,0,146,0,0,0,0,0,145,0,200,0,204,0,188,0,0,0,0,0,103,0,0,0,94,0,0,0,235,0,98,0,155,0,172,0,15,0,210,0,192,0,90,0,0,0,201,0,0,0,174,0,20,0,35,0,0,0,119,0,213,0,191,0,0,0,182,0,254,0,38,0,227,0,21,0,0,0,0,0,166,0,0,0,54,0,82,0,122,0,88,0,165,0,0,0,161,0,11,0,42,0,102,0,112,0,123,0,191,0,116,0,204,0,13,0,55,0,100,0,223,0,39,0,0,0,86,0,200,0,154,0,97,0,40,0,6,0,158,0,0,0,52,0,177,0,121,0,77,0,90,0,17,0,101,0,145,0,112,0,99,0,255,0,111,0,0,0,102,0,26,0,201,0,164,0,174,0,9,0,226,0,0,0,163,0,0,0,227,0,251,0,161,0,177,0,0,0,66,0,200,0,215,0,70,0,131,0,128,0,0,0,201,0,65,0,198,0,114,0,0,0,245,0,14,0,226,0,18,0,140,0,147,0,110,0,246,0,181,0,19,0,19,0,8,0,66,0,115,0,0,0,0,0,13,0,237,0,84,0,135,0,25,0,17,0,194,0,96,0,45,0,60,0,164,0,219,0,2,0,90,0,82,0,114,0,43,0,0,0,218,0,225,0,179,0,87,0,247,0,22,0,114,0,0,0,0,0,220,0,125,0,170,0,240,0,0,0,83,0,0,0,148,0,223,0,97,0,98,0,195,0,131,0,197,0,14,0,0,0,130,0);
signal scenario_full  : scenario_type := (140,31,11,31,47,31,31,31,33,31,194,31,180,31,114,31,115,31,33,31,11,31,63,31,42,31,42,30,253,31,180,31,182,31,43,31,241,31,248,31,87,31,49,31,29,31,33,31,171,31,79,31,107,31,34,31,32,31,32,30,245,31,192,31,216,31,51,31,51,31,16,31,72,31,64,31,64,30,178,31,237,31,26,31,127,31,207,31,14,31,160,31,160,30,137,31,152,31,13,31,125,31,243,31,243,30,206,31,34,31,137,31,107,31,107,30,196,31,212,31,137,31,227,31,213,31,213,30,19,31,113,31,204,31,117,31,80,31,229,31,9,31,76,31,23,31,23,30,7,31,7,30,75,31,128,31,128,30,162,31,39,31,200,31,163,31,163,30,163,29,163,28,107,31,30,31,75,31,224,31,89,31,118,31,220,31,102,31,248,31,157,31,88,31,115,31,167,31,96,31,194,31,177,31,23,31,137,31,72,31,20,31,89,31,83,31,221,31,11,31,11,30,48,31,55,31,45,31,235,31,246,31,246,30,23,31,228,31,64,31,64,30,45,31,125,31,186,31,58,31,68,31,213,31,213,30,187,31,126,31,94,31,135,31,74,31,140,31,140,30,99,31,4,31,180,31,50,31,72,31,13,31,214,31,243,31,243,30,243,29,227,31,57,31,86,31,61,31,36,31,3,31,29,31,236,31,93,31,54,31,54,30,238,31,72,31,252,31,240,31,252,31,60,31,60,30,141,31,247,31,107,31,67,31,28,31,157,31,46,31,86,31,78,31,175,31,51,31,194,31,194,30,76,31,78,31,44,31,94,31,198,31,165,31,165,30,218,31,218,30,218,29,73,31,182,31,182,30,83,31,83,30,56,31,56,30,56,29,56,28,34,31,61,31,175,31,189,31,180,31,27,31,23,31,35,31,83,31,9,31,134,31,231,31,219,31,19,31,83,31,116,31,59,31,202,31,202,30,71,31,57,31,3,31,44,31,185,31,142,31,192,31,8,31,8,30,30,31,12,31,156,31,69,31,140,31,11,31,11,30,39,31,121,31,250,31,250,30,84,31,41,31,94,31,65,31,144,31,49,31,152,31,113,31,42,31,49,31,8,31,198,31,149,31,7,31,119,31,119,30,119,29,254,31,38,31,34,31,1,31,156,31,216,31,216,30,65,31,65,30,67,31,103,31,195,31,138,31,157,31,48,31,81,31,81,30,154,31,251,31,214,31,150,31,119,31,231,31,12,31,151,31,34,31,185,31,185,30,185,29,60,31,60,30,70,31,86,31,155,31,71,31,226,31,218,31,13,31,13,30,88,31,8,31,196,31,58,31,58,30,131,31,87,31,87,30,107,31,107,30,201,31,125,31,169,31,210,31,194,31,204,31,105,31,46,31,241,31,219,31,187,31,117,31,23,31,23,30,23,29,46,31,168,31,50,31,142,31,142,30,88,31,149,31,46,31,39,31,83,31,34,31,176,31,243,31,230,31,56,31,56,30,31,31,178,31,138,31,38,31,38,30,103,31,103,30,159,31,243,31,242,31,206,31,183,31,42,31,19,31,19,30,199,31,37,31,100,31,58,31,137,31,137,30,164,31,193,31,199,31,10,31,168,31,147,31,47,31,192,31,96,31,96,30,110,31,142,31,103,31,195,31,195,30,248,31,40,31,196,31,196,30,196,29,196,28,196,27,108,31,179,31,87,31,199,31,220,31,161,31,89,31,82,31,193,31,213,31,49,31,127,31,127,31,59,31,113,31,18,31,247,31,247,30,126,31,16,31,179,31,12,31,159,31,13,31,249,31,231,31,53,31,252,31,180,31,173,31,173,30,63,31,50,31,96,31,77,31,59,31,13,31,202,31,251,31,251,30,251,29,16,31,236,31,43,31,10,31,185,31,65,31,80,31,217,31,195,31,195,30,20,31,210,31,210,30,194,31,194,30,221,31,221,30,43,31,173,31,152,31,179,31,42,31,39,31,78,31,136,31,136,30,227,31,134,31,123,31,196,31,56,31,188,31,188,31,153,31,153,30,138,31,138,30,138,29,72,31,147,31,28,31,14,31,166,31,164,31,214,31,7,31,231,31,117,31,117,30,59,31,27,31,32,31,217,31,91,31,189,31,189,30,3,31,59,31,59,30,59,29,54,31,134,31,134,30,12,31,18,31,98,31,98,30,98,29,98,28,125,31,197,31,93,31,196,31,109,31,135,31,38,31,91,31,55,31,175,31,236,31,204,31,136,31,11,31,251,31,165,31,203,31,218,31,161,31,230,31,139,31,122,31,150,31,150,30,46,31,121,31,12,31,176,31,176,30,139,31,188,31,210,31,236,31,13,31,13,30,177,31,248,31,4,31,128,31,128,30,101,31,101,30,75,31,75,30,233,31,135,31,210,31,31,31,246,31,164,31,92,31,92,30,92,29,57,31,78,31,34,31,34,30,151,31,151,30,151,29,126,31,69,31,92,31,154,31,224,31,89,31,94,31,169,31,169,30,143,31,143,30,139,31,138,31,212,31,38,31,142,31,175,31,175,30,175,29,72,31,112,31,160,31,160,30,12,31,123,31,193,31,189,31,189,30,202,31,115,31,38,31,13,31,216,31,166,31,18,31,43,31,43,30,1,31,1,30,46,31,208,31,209,31,181,31,181,30,237,31,236,31,233,31,233,30,233,29,78,31,78,30,38,31,38,30,169,31,154,31,154,30,210,31,60,31,109,31,111,31,58,31,58,30,249,31,12,31,214,31,214,31,113,31,113,30,99,31,243,31,50,31,47,31,47,31,47,30,187,31,253,31,213,31,174,31,17,31,143,31,143,30,142,31,142,30,144,31,81,31,26,31,78,31,78,30,78,29,30,31,45,31,140,31,215,31,55,31,11,31,58,31,49,31,28,31,80,31,80,30,134,31,189,31,188,31,52,31,96,31,57,31,103,31,35,31,243,31,60,31,1,31,178,31,85,31,20,31,20,30,198,31,139,31,139,30,51,31,233,31,53,31,108,31,129,31,129,30,91,31,201,31,145,31,131,31,131,30,169,31,171,31,209,31,7,31,141,31,230,31,230,30,230,29,125,31,249,31,190,31,121,31,52,31,156,31,176,31,176,30,5,31,5,30,33,31,33,30,82,31,231,31,203,31,58,31,86,31,250,31,241,31,42,31,60,31,60,30,60,29,55,31,172,31,162,31,62,31,195,31,163,31,163,30,95,31,161,31,251,31,238,31,200,31,102,31,102,30,251,31,115,31,254,31,102,31,22,31,53,31,109,31,165,31,189,31,151,31,8,31,235,31,235,30,144,31,144,30,145,31,246,31,40,31,69,31,47,31,88,31,117,31,117,30,214,31,214,30,214,29,189,31,87,31,87,30,61,31,200,31,200,30,237,31,65,31,145,31,205,31,87,31,134,31,134,30,8,31,8,30,78,31,73,31,17,31,106,31,41,31,41,30,94,31,131,31,131,30,69,31,114,31,146,31,42,31,42,30,114,31,43,31,43,30,134,31,252,31,212,31,32,31,69,31,146,31,146,30,146,29,145,31,200,31,204,31,188,31,188,30,188,29,103,31,103,30,94,31,94,30,235,31,98,31,155,31,172,31,15,31,210,31,192,31,90,31,90,30,201,31,201,30,174,31,20,31,35,31,35,30,119,31,213,31,191,31,191,30,182,31,254,31,38,31,227,31,21,31,21,30,21,29,166,31,166,30,54,31,82,31,122,31,88,31,165,31,165,30,161,31,11,31,42,31,102,31,112,31,123,31,191,31,116,31,204,31,13,31,55,31,100,31,223,31,39,31,39,30,86,31,200,31,154,31,97,31,40,31,6,31,158,31,158,30,52,31,177,31,121,31,77,31,90,31,17,31,101,31,145,31,112,31,99,31,255,31,111,31,111,30,102,31,26,31,201,31,164,31,174,31,9,31,226,31,226,30,163,31,163,30,227,31,251,31,161,31,177,31,177,30,66,31,200,31,215,31,70,31,131,31,128,31,128,30,201,31,65,31,198,31,114,31,114,30,245,31,14,31,226,31,18,31,140,31,147,31,110,31,246,31,181,31,19,31,19,31,8,31,66,31,115,31,115,30,115,29,13,31,237,31,84,31,135,31,25,31,17,31,194,31,96,31,45,31,60,31,164,31,219,31,2,31,90,31,82,31,114,31,43,31,43,30,218,31,225,31,179,31,87,31,247,31,22,31,114,31,114,30,114,29,220,31,125,31,170,31,240,31,240,30,83,31,83,30,148,31,223,31,97,31,98,31,195,31,131,31,197,31,14,31,14,30,130,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
