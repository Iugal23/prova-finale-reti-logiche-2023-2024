-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 665;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,0,0,150,0,189,0,196,0,94,0,67,0,0,0,216,0,189,0,91,0,232,0,215,0,78,0,29,0,185,0,39,0,66,0,0,0,52,0,222,0,231,0,252,0,80,0,242,0,146,0,0,0,38,0,36,0,0,0,203,0,229,0,154,0,230,0,55,0,133,0,162,0,3,0,0,0,36,0,0,0,16,0,111,0,135,0,0,0,39,0,189,0,85,0,175,0,134,0,181,0,223,0,206,0,0,0,0,0,102,0,161,0,110,0,255,0,0,0,238,0,90,0,254,0,197,0,67,0,251,0,0,0,67,0,169,0,249,0,91,0,216,0,171,0,9,0,223,0,135,0,224,0,140,0,236,0,0,0,0,0,104,0,32,0,182,0,132,0,0,0,0,0,21,0,76,0,58,0,196,0,99,0,36,0,235,0,0,0,94,0,9,0,94,0,237,0,94,0,221,0,229,0,0,0,0,0,153,0,147,0,0,0,122,0,183,0,231,0,167,0,0,0,98,0,157,0,0,0,97,0,67,0,239,0,18,0,236,0,135,0,0,0,5,0,0,0,0,0,82,0,148,0,225,0,91,0,31,0,182,0,0,0,0,0,0,0,73,0,0,0,0,0,197,0,144,0,19,0,0,0,183,0,119,0,4,0,141,0,201,0,202,0,0,0,0,0,73,0,120,0,123,0,0,0,125,0,236,0,14,0,112,0,228,0,63,0,157,0,138,0,18,0,104,0,98,0,201,0,40,0,0,0,0,0,98,0,70,0,239,0,87,0,8,0,100,0,160,0,133,0,123,0,117,0,252,0,157,0,39,0,110,0,48,0,96,0,57,0,199,0,234,0,196,0,105,0,6,0,187,0,241,0,14,0,232,0,146,0,35,0,144,0,184,0,27,0,0,0,44,0,177,0,151,0,83,0,0,0,56,0,19,0,66,0,18,0,186,0,0,0,46,0,160,0,59,0,45,0,0,0,134,0,0,0,0,0,200,0,160,0,5,0,108,0,25,0,0,0,244,0,183,0,129,0,136,0,162,0,66,0,63,0,129,0,0,0,0,0,0,0,251,0,0,0,143,0,214,0,239,0,0,0,0,0,0,0,64,0,4,0,35,0,194,0,248,0,0,0,0,0,249,0,158,0,82,0,0,0,56,0,183,0,0,0,208,0,207,0,130,0,213,0,54,0,0,0,80,0,229,0,241,0,0,0,90,0,0,0,133,0,118,0,0,0,7,0,169,0,92,0,10,0,0,0,34,0,219,0,235,0,32,0,221,0,214,0,0,0,0,0,253,0,16,0,60,0,145,0,160,0,0,0,51,0,93,0,131,0,84,0,215,0,106,0,179,0,195,0,26,0,32,0,173,0,0,0,15,0,134,0,92,0,225,0,100,0,240,0,0,0,31,0,123,0,191,0,205,0,134,0,122,0,238,0,183,0,45,0,132,0,33,0,0,0,40,0,236,0,46,0,26,0,0,0,34,0,0,0,0,0,75,0,62,0,11,0,83,0,0,0,120,0,152,0,148,0,157,0,186,0,132,0,227,0,53,0,0,0,164,0,94,0,182,0,226,0,51,0,49,0,84,0,34,0,144,0,0,0,216,0,232,0,174,0,31,0,19,0,0,0,96,0,75,0,74,0,158,0,52,0,0,0,0,0,170,0,93,0,0,0,90,0,67,0,238,0,19,0,72,0,5,0,147,0,74,0,4,0,79,0,241,0,0,0,154,0,244,0,48,0,15,0,0,0,0,0,126,0,189,0,196,0,0,0,11,0,0,0,224,0,233,0,0,0,77,0,222,0,243,0,165,0,0,0,199,0,168,0,212,0,197,0,34,0,193,0,0,0,42,0,225,0,0,0,25,0,110,0,55,0,0,0,107,0,69,0,39,0,147,0,0,0,68,0,32,0,212,0,239,0,253,0,53,0,152,0,89,0,205,0,117,0,127,0,144,0,109,0,0,0,195,0,170,0,68,0,176,0,248,0,149,0,148,0,235,0,61,0,0,0,76,0,124,0,88,0,231,0,0,0,145,0,85,0,9,0,242,0,45,0,14,0,161,0,240,0,53,0,163,0,138,0,144,0,21,0,120,0,211,0,26,0,236,0,94,0,47,0,101,0,0,0,6,0,202,0,235,0,188,0,0,0,0,0,22,0,201,0,162,0,98,0,164,0,0,0,162,0,107,0,72,0,0,0,59,0,0,0,253,0,231,0,60,0,61,0,245,0,188,0,0,0,30,0,98,0,125,0,0,0,114,0,114,0,251,0,150,0,171,0,168,0,161,0,20,0,0,0,215,0,157,0,215,0,194,0,158,0,107,0,38,0,0,0,14,0,247,0,242,0,48,0,0,0,0,0,224,0,7,0,180,0,2,0,0,0,2,0,67,0,102,0,253,0,240,0,0,0,81,0,184,0,22,0,78,0,142,0,0,0,107,0,147,0,0,0,0,0,107,0,89,0,58,0,137,0,160,0,0,0,166,0,177,0,0,0,163,0,125,0,99,0,155,0,186,0,212,0,0,0,0,0,19,0,212,0,242,0,65,0,213,0,229,0,0,0,0,0,166,0,0,0,215,0,40,0,35,0,250,0,137,0,141,0,143,0,0,0,0,0,237,0,39,0,203,0,194,0,189,0,108,0,0,0,83,0,14,0,0,0,227,0,214,0,221,0,0,0,97,0,0,0,0,0,213,0,0,0,0,0,206,0,72,0,9,0,1,0,240,0,180,0,246,0,121,0,122,0,247,0,238,0,67,0,52,0,138,0,198,0,6,0,180,0,103,0,0,0,185,0,183,0,5,0,153,0,0,0,224,0,131,0,247,0,108,0,228,0,188,0,152,0,209,0,164,0,0,0,0,0,0,0,158,0,250,0,248,0,132,0,30,0,147,0,129,0,118,0,198,0,34,0,197,0,120,0,0,0,19,0,238,0,146,0,17,0,224,0,154,0,0,0,1,0,0,0,0,0,128,0,157,0,58,0,132,0);
signal scenario_full  : scenario_type := (0,0,0,0,0,0,150,31,189,31,196,31,94,31,67,31,67,30,216,31,189,31,91,31,232,31,215,31,78,31,29,31,185,31,39,31,66,31,66,30,52,31,222,31,231,31,252,31,80,31,242,31,146,31,146,30,38,31,36,31,36,30,203,31,229,31,154,31,230,31,55,31,133,31,162,31,3,31,3,30,36,31,36,30,16,31,111,31,135,31,135,30,39,31,189,31,85,31,175,31,134,31,181,31,223,31,206,31,206,30,206,29,102,31,161,31,110,31,255,31,255,30,238,31,90,31,254,31,197,31,67,31,251,31,251,30,67,31,169,31,249,31,91,31,216,31,171,31,9,31,223,31,135,31,224,31,140,31,236,31,236,30,236,29,104,31,32,31,182,31,132,31,132,30,132,29,21,31,76,31,58,31,196,31,99,31,36,31,235,31,235,30,94,31,9,31,94,31,237,31,94,31,221,31,229,31,229,30,229,29,153,31,147,31,147,30,122,31,183,31,231,31,167,31,167,30,98,31,157,31,157,30,97,31,67,31,239,31,18,31,236,31,135,31,135,30,5,31,5,30,5,29,82,31,148,31,225,31,91,31,31,31,182,31,182,30,182,29,182,28,73,31,73,30,73,29,197,31,144,31,19,31,19,30,183,31,119,31,4,31,141,31,201,31,202,31,202,30,202,29,73,31,120,31,123,31,123,30,125,31,236,31,14,31,112,31,228,31,63,31,157,31,138,31,18,31,104,31,98,31,201,31,40,31,40,30,40,29,98,31,70,31,239,31,87,31,8,31,100,31,160,31,133,31,123,31,117,31,252,31,157,31,39,31,110,31,48,31,96,31,57,31,199,31,234,31,196,31,105,31,6,31,187,31,241,31,14,31,232,31,146,31,35,31,144,31,184,31,27,31,27,30,44,31,177,31,151,31,83,31,83,30,56,31,19,31,66,31,18,31,186,31,186,30,46,31,160,31,59,31,45,31,45,30,134,31,134,30,134,29,200,31,160,31,5,31,108,31,25,31,25,30,244,31,183,31,129,31,136,31,162,31,66,31,63,31,129,31,129,30,129,29,129,28,251,31,251,30,143,31,214,31,239,31,239,30,239,29,239,28,64,31,4,31,35,31,194,31,248,31,248,30,248,29,249,31,158,31,82,31,82,30,56,31,183,31,183,30,208,31,207,31,130,31,213,31,54,31,54,30,80,31,229,31,241,31,241,30,90,31,90,30,133,31,118,31,118,30,7,31,169,31,92,31,10,31,10,30,34,31,219,31,235,31,32,31,221,31,214,31,214,30,214,29,253,31,16,31,60,31,145,31,160,31,160,30,51,31,93,31,131,31,84,31,215,31,106,31,179,31,195,31,26,31,32,31,173,31,173,30,15,31,134,31,92,31,225,31,100,31,240,31,240,30,31,31,123,31,191,31,205,31,134,31,122,31,238,31,183,31,45,31,132,31,33,31,33,30,40,31,236,31,46,31,26,31,26,30,34,31,34,30,34,29,75,31,62,31,11,31,83,31,83,30,120,31,152,31,148,31,157,31,186,31,132,31,227,31,53,31,53,30,164,31,94,31,182,31,226,31,51,31,49,31,84,31,34,31,144,31,144,30,216,31,232,31,174,31,31,31,19,31,19,30,96,31,75,31,74,31,158,31,52,31,52,30,52,29,170,31,93,31,93,30,90,31,67,31,238,31,19,31,72,31,5,31,147,31,74,31,4,31,79,31,241,31,241,30,154,31,244,31,48,31,15,31,15,30,15,29,126,31,189,31,196,31,196,30,11,31,11,30,224,31,233,31,233,30,77,31,222,31,243,31,165,31,165,30,199,31,168,31,212,31,197,31,34,31,193,31,193,30,42,31,225,31,225,30,25,31,110,31,55,31,55,30,107,31,69,31,39,31,147,31,147,30,68,31,32,31,212,31,239,31,253,31,53,31,152,31,89,31,205,31,117,31,127,31,144,31,109,31,109,30,195,31,170,31,68,31,176,31,248,31,149,31,148,31,235,31,61,31,61,30,76,31,124,31,88,31,231,31,231,30,145,31,85,31,9,31,242,31,45,31,14,31,161,31,240,31,53,31,163,31,138,31,144,31,21,31,120,31,211,31,26,31,236,31,94,31,47,31,101,31,101,30,6,31,202,31,235,31,188,31,188,30,188,29,22,31,201,31,162,31,98,31,164,31,164,30,162,31,107,31,72,31,72,30,59,31,59,30,253,31,231,31,60,31,61,31,245,31,188,31,188,30,30,31,98,31,125,31,125,30,114,31,114,31,251,31,150,31,171,31,168,31,161,31,20,31,20,30,215,31,157,31,215,31,194,31,158,31,107,31,38,31,38,30,14,31,247,31,242,31,48,31,48,30,48,29,224,31,7,31,180,31,2,31,2,30,2,31,67,31,102,31,253,31,240,31,240,30,81,31,184,31,22,31,78,31,142,31,142,30,107,31,147,31,147,30,147,29,107,31,89,31,58,31,137,31,160,31,160,30,166,31,177,31,177,30,163,31,125,31,99,31,155,31,186,31,212,31,212,30,212,29,19,31,212,31,242,31,65,31,213,31,229,31,229,30,229,29,166,31,166,30,215,31,40,31,35,31,250,31,137,31,141,31,143,31,143,30,143,29,237,31,39,31,203,31,194,31,189,31,108,31,108,30,83,31,14,31,14,30,227,31,214,31,221,31,221,30,97,31,97,30,97,29,213,31,213,30,213,29,206,31,72,31,9,31,1,31,240,31,180,31,246,31,121,31,122,31,247,31,238,31,67,31,52,31,138,31,198,31,6,31,180,31,103,31,103,30,185,31,183,31,5,31,153,31,153,30,224,31,131,31,247,31,108,31,228,31,188,31,152,31,209,31,164,31,164,30,164,29,164,28,158,31,250,31,248,31,132,31,30,31,147,31,129,31,118,31,198,31,34,31,197,31,120,31,120,30,19,31,238,31,146,31,17,31,224,31,154,31,154,30,1,31,1,30,1,29,128,31,157,31,58,31,132,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
