-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 464;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (186,0,0,0,158,0,110,0,66,0,224,0,0,0,128,0,228,0,71,0,9,0,53,0,22,0,29,0,164,0,82,0,134,0,206,0,53,0,68,0,0,0,5,0,184,0,190,0,0,0,156,0,168,0,93,0,105,0,32,0,0,0,255,0,215,0,159,0,79,0,144,0,17,0,0,0,0,0,95,0,0,0,96,0,166,0,121,0,0,0,151,0,154,0,0,0,204,0,201,0,0,0,188,0,71,0,0,0,32,0,34,0,62,0,8,0,191,0,189,0,0,0,0,0,163,0,176,0,0,0,0,0,171,0,189,0,0,0,225,0,14,0,167,0,0,0,211,0,210,0,0,0,207,0,56,0,254,0,156,0,164,0,132,0,88,0,25,0,113,0,249,0,245,0,0,0,166,0,133,0,21,0,0,0,241,0,220,0,83,0,0,0,37,0,135,0,0,0,15,0,178,0,90,0,132,0,205,0,90,0,26,0,83,0,217,0,0,0,0,0,161,0,185,0,74,0,205,0,67,0,0,0,237,0,36,0,3,0,186,0,231,0,0,0,0,0,0,0,124,0,222,0,209,0,98,0,139,0,155,0,214,0,25,0,0,0,240,0,25,0,0,0,6,0,20,0,202,0,207,0,113,0,147,0,190,0,0,0,37,0,7,0,0,0,213,0,0,0,214,0,222,0,94,0,0,0,134,0,228,0,165,0,0,0,8,0,81,0,131,0,197,0,0,0,37,0,204,0,211,0,148,0,210,0,74,0,173,0,16,0,233,0,190,0,218,0,107,0,0,0,103,0,125,0,37,0,36,0,214,0,211,0,167,0,174,0,77,0,132,0,0,0,20,0,158,0,62,0,38,0,83,0,0,0,0,0,34,0,5,0,24,0,0,0,249,0,163,0,117,0,198,0,158,0,39,0,0,0,85,0,62,0,55,0,0,0,188,0,106,0,223,0,238,0,31,0,8,0,103,0,0,0,0,0,185,0,0,0,125,0,44,0,130,0,0,0,233,0,222,0,208,0,197,0,0,0,90,0,117,0,106,0,92,0,0,0,89,0,0,0,117,0,240,0,14,0,0,0,80,0,117,0,95,0,242,0,0,0,13,0,74,0,41,0,0,0,32,0,197,0,13,0,0,0,0,0,0,0,140,0,39,0,79,0,0,0,180,0,119,0,252,0,173,0,219,0,174,0,215,0,245,0,0,0,127,0,218,0,0,0,233,0,14,0,115,0,62,0,244,0,55,0,202,0,0,0,82,0,140,0,92,0,132,0,79,0,11,0,157,0,8,0,19,0,213,0,124,0,129,0,144,0,13,0,6,0,0,0,15,0,83,0,122,0,47,0,8,0,217,0,132,0,9,0,149,0,193,0,0,0,0,0,209,0,87,0,0,0,23,0,227,0,202,0,180,0,226,0,188,0,0,0,142,0,69,0,0,0,49,0,139,0,0,0,0,0,147,0,0,0,103,0,185,0,84,0,192,0,27,0,230,0,0,0,20,0,46,0,0,0,0,0,86,0,185,0,238,0,167,0,41,0,71,0,30,0,246,0,105,0,0,0,72,0,28,0,134,0,101,0,233,0,86,0,143,0,229,0,101,0,231,0,14,0,20,0,47,0,146,0,255,0,66,0,3,0,217,0,112,0,118,0,0,0,127,0,7,0,28,0,18,0,54,0,21,0,167,0,123,0,0,0,20,0,0,0,19,0,176,0,0,0,201,0,33,0,0,0,0,0,59,0,222,0,61,0,142,0,38,0,11,0,58,0,20,0,30,0,113,0,97,0,109,0,225,0,36,0,106,0,254,0,4,0,0,0,249,0,56,0,0,0,198,0,143,0,183,0,0,0,81,0,123,0,94,0,100,0,143,0,17,0,176,0,209,0,90,0,236,0,16,0,67,0,192,0,191,0,0,0,159,0,226,0,0,0,0,0,0,0,117,0,227,0,246,0,158,0,65,0,0,0,223,0,0,0,171,0,73,0,107,0,242,0,0,0,0,0,215,0,225,0,159,0,192,0,218,0,254,0,71,0,61,0,9,0,97,0,104,0,60,0,106,0,63,0,88,0,45,0,244,0,117,0,85,0,208,0);
signal scenario_full  : scenario_type := (186,31,186,30,158,31,110,31,66,31,224,31,224,30,128,31,228,31,71,31,9,31,53,31,22,31,29,31,164,31,82,31,134,31,206,31,53,31,68,31,68,30,5,31,184,31,190,31,190,30,156,31,168,31,93,31,105,31,32,31,32,30,255,31,215,31,159,31,79,31,144,31,17,31,17,30,17,29,95,31,95,30,96,31,166,31,121,31,121,30,151,31,154,31,154,30,204,31,201,31,201,30,188,31,71,31,71,30,32,31,34,31,62,31,8,31,191,31,189,31,189,30,189,29,163,31,176,31,176,30,176,29,171,31,189,31,189,30,225,31,14,31,167,31,167,30,211,31,210,31,210,30,207,31,56,31,254,31,156,31,164,31,132,31,88,31,25,31,113,31,249,31,245,31,245,30,166,31,133,31,21,31,21,30,241,31,220,31,83,31,83,30,37,31,135,31,135,30,15,31,178,31,90,31,132,31,205,31,90,31,26,31,83,31,217,31,217,30,217,29,161,31,185,31,74,31,205,31,67,31,67,30,237,31,36,31,3,31,186,31,231,31,231,30,231,29,231,28,124,31,222,31,209,31,98,31,139,31,155,31,214,31,25,31,25,30,240,31,25,31,25,30,6,31,20,31,202,31,207,31,113,31,147,31,190,31,190,30,37,31,7,31,7,30,213,31,213,30,214,31,222,31,94,31,94,30,134,31,228,31,165,31,165,30,8,31,81,31,131,31,197,31,197,30,37,31,204,31,211,31,148,31,210,31,74,31,173,31,16,31,233,31,190,31,218,31,107,31,107,30,103,31,125,31,37,31,36,31,214,31,211,31,167,31,174,31,77,31,132,31,132,30,20,31,158,31,62,31,38,31,83,31,83,30,83,29,34,31,5,31,24,31,24,30,249,31,163,31,117,31,198,31,158,31,39,31,39,30,85,31,62,31,55,31,55,30,188,31,106,31,223,31,238,31,31,31,8,31,103,31,103,30,103,29,185,31,185,30,125,31,44,31,130,31,130,30,233,31,222,31,208,31,197,31,197,30,90,31,117,31,106,31,92,31,92,30,89,31,89,30,117,31,240,31,14,31,14,30,80,31,117,31,95,31,242,31,242,30,13,31,74,31,41,31,41,30,32,31,197,31,13,31,13,30,13,29,13,28,140,31,39,31,79,31,79,30,180,31,119,31,252,31,173,31,219,31,174,31,215,31,245,31,245,30,127,31,218,31,218,30,233,31,14,31,115,31,62,31,244,31,55,31,202,31,202,30,82,31,140,31,92,31,132,31,79,31,11,31,157,31,8,31,19,31,213,31,124,31,129,31,144,31,13,31,6,31,6,30,15,31,83,31,122,31,47,31,8,31,217,31,132,31,9,31,149,31,193,31,193,30,193,29,209,31,87,31,87,30,23,31,227,31,202,31,180,31,226,31,188,31,188,30,142,31,69,31,69,30,49,31,139,31,139,30,139,29,147,31,147,30,103,31,185,31,84,31,192,31,27,31,230,31,230,30,20,31,46,31,46,30,46,29,86,31,185,31,238,31,167,31,41,31,71,31,30,31,246,31,105,31,105,30,72,31,28,31,134,31,101,31,233,31,86,31,143,31,229,31,101,31,231,31,14,31,20,31,47,31,146,31,255,31,66,31,3,31,217,31,112,31,118,31,118,30,127,31,7,31,28,31,18,31,54,31,21,31,167,31,123,31,123,30,20,31,20,30,19,31,176,31,176,30,201,31,33,31,33,30,33,29,59,31,222,31,61,31,142,31,38,31,11,31,58,31,20,31,30,31,113,31,97,31,109,31,225,31,36,31,106,31,254,31,4,31,4,30,249,31,56,31,56,30,198,31,143,31,183,31,183,30,81,31,123,31,94,31,100,31,143,31,17,31,176,31,209,31,90,31,236,31,16,31,67,31,192,31,191,31,191,30,159,31,226,31,226,30,226,29,226,28,117,31,227,31,246,31,158,31,65,31,65,30,223,31,223,30,171,31,73,31,107,31,242,31,242,30,242,29,215,31,225,31,159,31,192,31,218,31,254,31,71,31,61,31,9,31,97,31,104,31,60,31,106,31,63,31,88,31,45,31,244,31,117,31,85,31,208,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
