-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 993;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (197,0,118,0,0,0,55,0,96,0,201,0,177,0,0,0,0,0,0,0,0,0,0,0,206,0,216,0,38,0,219,0,187,0,0,0,21,0,181,0,186,0,135,0,195,0,152,0,137,0,184,0,43,0,81,0,151,0,154,0,0,0,120,0,107,0,165,0,198,0,17,0,12,0,56,0,187,0,33,0,0,0,128,0,118,0,168,0,92,0,229,0,143,0,228,0,207,0,44,0,144,0,108,0,57,0,45,0,156,0,0,0,78,0,206,0,134,0,126,0,200,0,0,0,0,0,235,0,0,0,220,0,254,0,241,0,73,0,222,0,0,0,26,0,112,0,0,0,208,0,137,0,0,0,143,0,94,0,0,0,0,0,0,0,191,0,0,0,95,0,41,0,0,0,0,0,0,0,112,0,0,0,80,0,190,0,236,0,110,0,70,0,156,0,91,0,49,0,7,0,0,0,0,0,196,0,108,0,0,0,102,0,0,0,55,0,0,0,0,0,0,0,77,0,158,0,247,0,85,0,0,0,109,0,74,0,214,0,143,0,128,0,174,0,75,0,19,0,183,0,204,0,2,0,0,0,225,0,8,0,8,0,103,0,129,0,25,0,0,0,193,0,229,0,0,0,7,0,0,0,21,0,18,0,14,0,130,0,68,0,17,0,125,0,141,0,112,0,248,0,130,0,168,0,10,0,0,0,162,0,184,0,142,0,0,0,210,0,136,0,113,0,0,0,0,0,189,0,0,0,2,0,191,0,58,0,235,0,22,0,82,0,250,0,0,0,0,0,139,0,140,0,34,0,0,0,157,0,87,0,253,0,144,0,0,0,46,0,0,0,0,0,108,0,92,0,0,0,243,0,146,0,110,0,1,0,18,0,0,0,229,0,255,0,218,0,144,0,0,0,125,0,105,0,218,0,35,0,22,0,72,0,191,0,102,0,146,0,90,0,208,0,0,0,29,0,125,0,0,0,166,0,77,0,58,0,51,0,77,0,194,0,0,0,232,0,209,0,12,0,103,0,249,0,0,0,137,0,157,0,40,0,0,0,0,0,141,0,62,0,133,0,122,0,142,0,208,0,141,0,240,0,0,0,0,0,119,0,81,0,122,0,255,0,0,0,31,0,211,0,0,0,225,0,69,0,92,0,214,0,48,0,0,0,245,0,27,0,8,0,102,0,78,0,235,0,64,0,106,0,50,0,154,0,177,0,62,0,0,0,116,0,46,0,122,0,0,0,236,0,228,0,223,0,128,0,142,0,62,0,198,0,73,0,113,0,215,0,181,0,54,0,154,0,85,0,163,0,169,0,126,0,80,0,8,0,100,0,155,0,19,0,0,0,0,0,0,0,86,0,0,0,31,0,111,0,211,0,243,0,213,0,0,0,0,0,126,0,195,0,0,0,219,0,71,0,0,0,12,0,0,0,223,0,219,0,165,0,0,0,61,0,224,0,107,0,209,0,119,0,10,0,0,0,233,0,56,0,0,0,0,0,0,0,18,0,16,0,0,0,240,0,44,0,0,0,216,0,172,0,201,0,0,0,144,0,42,0,188,0,15,0,57,0,36,0,116,0,118,0,82,0,10,0,113,0,18,0,71,0,204,0,162,0,40,0,0,0,155,0,138,0,235,0,0,0,236,0,135,0,228,0,226,0,43,0,186,0,140,0,248,0,99,0,228,0,149,0,209,0,0,0,0,0,131,0,252,0,199,0,96,0,0,0,16,0,133,0,129,0,0,0,23,0,7,0,1,0,147,0,202,0,134,0,72,0,226,0,0,0,76,0,96,0,0,0,245,0,0,0,27,0,0,0,55,0,70,0,74,0,58,0,86,0,174,0,232,0,0,0,0,0,68,0,172,0,0,0,159,0,202,0,90,0,87,0,33,0,5,0,50,0,123,0,231,0,26,0,64,0,90,0,0,0,141,0,0,0,176,0,0,0,8,0,213,0,195,0,0,0,0,0,152,0,204,0,3,0,125,0,214,0,90,0,78,0,141,0,111,0,160,0,207,0,66,0,249,0,181,0,39,0,137,0,120,0,38,0,0,0,127,0,21,0,9,0,116,0,243,0,178,0,89,0,242,0,58,0,117,0,235,0,104,0,41,0,142,0,81,0,139,0,0,0,204,0,14,0,61,0,4,0,0,0,223,0,172,0,39,0,216,0,90,0,0,0,0,0,67,0,102,0,207,0,239,0,213,0,48,0,0,0,50,0,0,0,18,0,80,0,148,0,106,0,34,0,226,0,55,0,0,0,0,0,219,0,0,0,175,0,41,0,44,0,128,0,0,0,0,0,179,0,167,0,66,0,65,0,64,0,215,0,0,0,208,0,23,0,13,0,133,0,226,0,0,0,131,0,15,0,244,0,191,0,144,0,0,0,102,0,0,0,238,0,227,0,186,0,174,0,215,0,50,0,11,0,238,0,47,0,161,0,0,0,214,0,182,0,10,0,29,0,98,0,209,0,182,0,49,0,213,0,172,0,251,0,0,0,114,0,37,0,162,0,255,0,212,0,107,0,254,0,184,0,0,0,0,0,0,0,217,0,0,0,92,0,155,0,223,0,250,0,173,0,48,0,193,0,37,0,68,0,239,0,8,0,120,0,195,0,0,0,3,0,89,0,37,0,169,0,0,0,36,0,216,0,131,0,110,0,135,0,50,0,213,0,228,0,192,0,14,0,71,0,0,0,63,0,252,0,0,0,16,0,1,0,169,0,0,0,251,0,182,0,95,0,64,0,2,0,246,0,206,0,149,0,27,0,27,0,66,0,163,0,89,0,148,0,0,0,220,0,135,0,6,0,157,0,127,0,247,0,0,0,0,0,122,0,156,0,116,0,0,0,144,0,73,0,160,0,188,0,159,0,153,0,0,0,104,0,0,0,28,0,0,0,113,0,0,0,0,0,230,0,170,0,170,0,161,0,138,0,157,0,61,0,122,0,163,0,190,0,87,0,128,0,160,0,150,0,65,0,187,0,203,0,93,0,39,0,127,0,130,0,141,0,30,0,65,0,31,0,39,0,162,0,161,0,2,0,226,0,0,0,102,0,0,0,57,0,108,0,71,0,0,0,185,0,66,0,22,0,16,0,147,0,229,0,0,0,122,0,0,0,146,0,220,0,0,0,205,0,88,0,94,0,149,0,0,0,45,0,0,0,157,0,227,0,139,0,48,0,0,0,0,0,210,0,0,0,101,0,225,0,249,0,0,0,207,0,91,0,0,0,6,0,200,0,0,0,41,0,121,0,0,0,172,0,97,0,0,0,167,0,22,0,139,0,139,0,119,0,26,0,47,0,79,0,63,0,94,0,55,0,120,0,0,0,22,0,61,0,144,0,161,0,84,0,10,0,0,0,0,0,210,0,251,0,184,0,0,0,136,0,82,0,215,0,250,0,118,0,52,0,0,0,220,0,30,0,225,0,76,0,28,0,0,0,117,0,0,0,242,0,119,0,249,0,101,0,104,0,127,0,79,0,214,0,41,0,128,0,162,0,225,0,27,0,240,0,0,0,131,0,162,0,244,0,108,0,161,0,113,0,192,0,9,0,131,0,172,0,32,0,172,0,100,0,70,0,0,0,251,0,0,0,119,0,41,0,115,0,169,0,20,0,61,0,0,0,88,0,58,0,187,0,185,0,21,0,100,0,0,0,225,0,224,0,0,0,131,0,239,0,0,0,34,0,81,0,86,0,150,0,0,0,182,0,218,0,0,0,87,0,155,0,48,0,14,0,100,0,165,0,0,0,107,0,172,0,94,0,0,0,124,0,41,0,182,0,10,0,0,0,221,0,0,0,42,0,0,0,84,0,188,0,183,0,216,0,60,0,0,0,132,0,186,0,198,0,141,0,10,0,147,0,52,0,0,0,104,0,78,0,0,0,14,0,103,0,149,0,214,0,172,0,209,0,69,0,76,0,0,0,244,0,210,0,99,0,179,0,207,0,0,0,143,0,2,0,0,0,0,0,5,0,0,0,0,0,18,0,198,0,225,0,137,0,35,0,0,0,153,0,120,0,222,0,71,0,82,0,43,0,16,0,114,0,0,0,248,0,14,0,23,0,207,0,19,0,190,0,114,0,24,0,34,0,173,0,168,0,179,0,12,0,105,0,0,0,0,0,0,0,217,0,225,0,54,0,163,0,254,0,245,0,37,0,4,0,168,0,14,0,161,0,236,0,0,0,250,0,209,0,192,0,0,0,251,0,127,0,0,0,190,0,188,0,0,0,51,0,66,0,0,0,194,0,148,0,208,0,0,0,23,0,15,0,129,0,252,0,75,0,196,0,207,0,120,0,51,0,0,0,0,0,28,0,226,0,227,0,0,0,0,0,193,0,241,0,0,0,94,0,123,0,119,0,0,0,250,0,194,0,0,0,0,0,241,0,0,0,0,0,59,0,127,0,156,0,20,0,18,0,43,0,96,0,0,0,26,0,193,0,128,0,79,0,103,0,0,0,188,0,127,0);
signal scenario_full  : scenario_type := (197,31,118,31,118,30,55,31,96,31,201,31,177,31,177,30,177,29,177,28,177,27,177,26,206,31,216,31,38,31,219,31,187,31,187,30,21,31,181,31,186,31,135,31,195,31,152,31,137,31,184,31,43,31,81,31,151,31,154,31,154,30,120,31,107,31,165,31,198,31,17,31,12,31,56,31,187,31,33,31,33,30,128,31,118,31,168,31,92,31,229,31,143,31,228,31,207,31,44,31,144,31,108,31,57,31,45,31,156,31,156,30,78,31,206,31,134,31,126,31,200,31,200,30,200,29,235,31,235,30,220,31,254,31,241,31,73,31,222,31,222,30,26,31,112,31,112,30,208,31,137,31,137,30,143,31,94,31,94,30,94,29,94,28,191,31,191,30,95,31,41,31,41,30,41,29,41,28,112,31,112,30,80,31,190,31,236,31,110,31,70,31,156,31,91,31,49,31,7,31,7,30,7,29,196,31,108,31,108,30,102,31,102,30,55,31,55,30,55,29,55,28,77,31,158,31,247,31,85,31,85,30,109,31,74,31,214,31,143,31,128,31,174,31,75,31,19,31,183,31,204,31,2,31,2,30,225,31,8,31,8,31,103,31,129,31,25,31,25,30,193,31,229,31,229,30,7,31,7,30,21,31,18,31,14,31,130,31,68,31,17,31,125,31,141,31,112,31,248,31,130,31,168,31,10,31,10,30,162,31,184,31,142,31,142,30,210,31,136,31,113,31,113,30,113,29,189,31,189,30,2,31,191,31,58,31,235,31,22,31,82,31,250,31,250,30,250,29,139,31,140,31,34,31,34,30,157,31,87,31,253,31,144,31,144,30,46,31,46,30,46,29,108,31,92,31,92,30,243,31,146,31,110,31,1,31,18,31,18,30,229,31,255,31,218,31,144,31,144,30,125,31,105,31,218,31,35,31,22,31,72,31,191,31,102,31,146,31,90,31,208,31,208,30,29,31,125,31,125,30,166,31,77,31,58,31,51,31,77,31,194,31,194,30,232,31,209,31,12,31,103,31,249,31,249,30,137,31,157,31,40,31,40,30,40,29,141,31,62,31,133,31,122,31,142,31,208,31,141,31,240,31,240,30,240,29,119,31,81,31,122,31,255,31,255,30,31,31,211,31,211,30,225,31,69,31,92,31,214,31,48,31,48,30,245,31,27,31,8,31,102,31,78,31,235,31,64,31,106,31,50,31,154,31,177,31,62,31,62,30,116,31,46,31,122,31,122,30,236,31,228,31,223,31,128,31,142,31,62,31,198,31,73,31,113,31,215,31,181,31,54,31,154,31,85,31,163,31,169,31,126,31,80,31,8,31,100,31,155,31,19,31,19,30,19,29,19,28,86,31,86,30,31,31,111,31,211,31,243,31,213,31,213,30,213,29,126,31,195,31,195,30,219,31,71,31,71,30,12,31,12,30,223,31,219,31,165,31,165,30,61,31,224,31,107,31,209,31,119,31,10,31,10,30,233,31,56,31,56,30,56,29,56,28,18,31,16,31,16,30,240,31,44,31,44,30,216,31,172,31,201,31,201,30,144,31,42,31,188,31,15,31,57,31,36,31,116,31,118,31,82,31,10,31,113,31,18,31,71,31,204,31,162,31,40,31,40,30,155,31,138,31,235,31,235,30,236,31,135,31,228,31,226,31,43,31,186,31,140,31,248,31,99,31,228,31,149,31,209,31,209,30,209,29,131,31,252,31,199,31,96,31,96,30,16,31,133,31,129,31,129,30,23,31,7,31,1,31,147,31,202,31,134,31,72,31,226,31,226,30,76,31,96,31,96,30,245,31,245,30,27,31,27,30,55,31,70,31,74,31,58,31,86,31,174,31,232,31,232,30,232,29,68,31,172,31,172,30,159,31,202,31,90,31,87,31,33,31,5,31,50,31,123,31,231,31,26,31,64,31,90,31,90,30,141,31,141,30,176,31,176,30,8,31,213,31,195,31,195,30,195,29,152,31,204,31,3,31,125,31,214,31,90,31,78,31,141,31,111,31,160,31,207,31,66,31,249,31,181,31,39,31,137,31,120,31,38,31,38,30,127,31,21,31,9,31,116,31,243,31,178,31,89,31,242,31,58,31,117,31,235,31,104,31,41,31,142,31,81,31,139,31,139,30,204,31,14,31,61,31,4,31,4,30,223,31,172,31,39,31,216,31,90,31,90,30,90,29,67,31,102,31,207,31,239,31,213,31,48,31,48,30,50,31,50,30,18,31,80,31,148,31,106,31,34,31,226,31,55,31,55,30,55,29,219,31,219,30,175,31,41,31,44,31,128,31,128,30,128,29,179,31,167,31,66,31,65,31,64,31,215,31,215,30,208,31,23,31,13,31,133,31,226,31,226,30,131,31,15,31,244,31,191,31,144,31,144,30,102,31,102,30,238,31,227,31,186,31,174,31,215,31,50,31,11,31,238,31,47,31,161,31,161,30,214,31,182,31,10,31,29,31,98,31,209,31,182,31,49,31,213,31,172,31,251,31,251,30,114,31,37,31,162,31,255,31,212,31,107,31,254,31,184,31,184,30,184,29,184,28,217,31,217,30,92,31,155,31,223,31,250,31,173,31,48,31,193,31,37,31,68,31,239,31,8,31,120,31,195,31,195,30,3,31,89,31,37,31,169,31,169,30,36,31,216,31,131,31,110,31,135,31,50,31,213,31,228,31,192,31,14,31,71,31,71,30,63,31,252,31,252,30,16,31,1,31,169,31,169,30,251,31,182,31,95,31,64,31,2,31,246,31,206,31,149,31,27,31,27,31,66,31,163,31,89,31,148,31,148,30,220,31,135,31,6,31,157,31,127,31,247,31,247,30,247,29,122,31,156,31,116,31,116,30,144,31,73,31,160,31,188,31,159,31,153,31,153,30,104,31,104,30,28,31,28,30,113,31,113,30,113,29,230,31,170,31,170,31,161,31,138,31,157,31,61,31,122,31,163,31,190,31,87,31,128,31,160,31,150,31,65,31,187,31,203,31,93,31,39,31,127,31,130,31,141,31,30,31,65,31,31,31,39,31,162,31,161,31,2,31,226,31,226,30,102,31,102,30,57,31,108,31,71,31,71,30,185,31,66,31,22,31,16,31,147,31,229,31,229,30,122,31,122,30,146,31,220,31,220,30,205,31,88,31,94,31,149,31,149,30,45,31,45,30,157,31,227,31,139,31,48,31,48,30,48,29,210,31,210,30,101,31,225,31,249,31,249,30,207,31,91,31,91,30,6,31,200,31,200,30,41,31,121,31,121,30,172,31,97,31,97,30,167,31,22,31,139,31,139,31,119,31,26,31,47,31,79,31,63,31,94,31,55,31,120,31,120,30,22,31,61,31,144,31,161,31,84,31,10,31,10,30,10,29,210,31,251,31,184,31,184,30,136,31,82,31,215,31,250,31,118,31,52,31,52,30,220,31,30,31,225,31,76,31,28,31,28,30,117,31,117,30,242,31,119,31,249,31,101,31,104,31,127,31,79,31,214,31,41,31,128,31,162,31,225,31,27,31,240,31,240,30,131,31,162,31,244,31,108,31,161,31,113,31,192,31,9,31,131,31,172,31,32,31,172,31,100,31,70,31,70,30,251,31,251,30,119,31,41,31,115,31,169,31,20,31,61,31,61,30,88,31,58,31,187,31,185,31,21,31,100,31,100,30,225,31,224,31,224,30,131,31,239,31,239,30,34,31,81,31,86,31,150,31,150,30,182,31,218,31,218,30,87,31,155,31,48,31,14,31,100,31,165,31,165,30,107,31,172,31,94,31,94,30,124,31,41,31,182,31,10,31,10,30,221,31,221,30,42,31,42,30,84,31,188,31,183,31,216,31,60,31,60,30,132,31,186,31,198,31,141,31,10,31,147,31,52,31,52,30,104,31,78,31,78,30,14,31,103,31,149,31,214,31,172,31,209,31,69,31,76,31,76,30,244,31,210,31,99,31,179,31,207,31,207,30,143,31,2,31,2,30,2,29,5,31,5,30,5,29,18,31,198,31,225,31,137,31,35,31,35,30,153,31,120,31,222,31,71,31,82,31,43,31,16,31,114,31,114,30,248,31,14,31,23,31,207,31,19,31,190,31,114,31,24,31,34,31,173,31,168,31,179,31,12,31,105,31,105,30,105,29,105,28,217,31,225,31,54,31,163,31,254,31,245,31,37,31,4,31,168,31,14,31,161,31,236,31,236,30,250,31,209,31,192,31,192,30,251,31,127,31,127,30,190,31,188,31,188,30,51,31,66,31,66,30,194,31,148,31,208,31,208,30,23,31,15,31,129,31,252,31,75,31,196,31,207,31,120,31,51,31,51,30,51,29,28,31,226,31,227,31,227,30,227,29,193,31,241,31,241,30,94,31,123,31,119,31,119,30,250,31,194,31,194,30,194,29,241,31,241,30,241,29,59,31,127,31,156,31,20,31,18,31,43,31,96,31,96,30,26,31,193,31,128,31,79,31,103,31,103,30,188,31,127,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
