-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 311;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (139,0,22,0,34,0,110,0,167,0,210,0,38,0,238,0,95,0,0,0,0,0,178,0,26,0,144,0,0,0,0,0,135,0,250,0,0,0,228,0,0,0,88,0,136,0,238,0,93,0,94,0,146,0,135,0,13,0,0,0,152,0,236,0,0,0,0,0,187,0,0,0,55,0,9,0,163,0,168,0,47,0,0,0,142,0,150,0,224,0,94,0,75,0,90,0,58,0,108,0,190,0,0,0,0,0,56,0,0,0,27,0,26,0,211,0,112,0,189,0,144,0,65,0,207,0,252,0,110,0,102,0,10,0,218,0,0,0,126,0,255,0,88,0,181,0,75,0,30,0,0,0,248,0,185,0,92,0,0,0,0,0,212,0,0,0,0,0,28,0,226,0,253,0,35,0,140,0,15,0,163,0,54,0,141,0,183,0,46,0,207,0,24,0,0,0,230,0,246,0,72,0,71,0,102,0,69,0,125,0,0,0,129,0,226,0,147,0,248,0,203,0,0,0,150,0,144,0,0,0,217,0,160,0,178,0,111,0,0,0,0,0,32,0,198,0,0,0,122,0,163,0,0,0,123,0,0,0,0,0,232,0,0,0,0,0,0,0,18,0,89,0,190,0,72,0,73,0,0,0,248,0,211,0,173,0,154,0,159,0,121,0,162,0,0,0,149,0,127,0,0,0,17,0,131,0,227,0,0,0,164,0,29,0,15,0,48,0,0,0,0,0,255,0,208,0,219,0,216,0,0,0,65,0,124,0,0,0,230,0,124,0,245,0,103,0,131,0,252,0,22,0,27,0,132,0,88,0,0,0,0,0,0,0,0,0,64,0,0,0,130,0,34,0,98,0,197,0,25,0,81,0,142,0,201,0,168,0,246,0,0,0,213,0,0,0,0,0,15,0,0,0,155,0,175,0,0,0,83,0,68,0,33,0,69,0,191,0,42,0,192,0,0,0,45,0,38,0,0,0,146,0,253,0,29,0,90,0,233,0,224,0,44,0,209,0,75,0,25,0,141,0,122,0,45,0,142,0,0,0,27,0,154,0,135,0,0,0,101,0,230,0,0,0,242,0,6,0,172,0,0,0,0,0,50,0,243,0,214,0,119,0,27,0,62,0,3,0,114,0,144,0,98,0,126,0,197,0,81,0,95,0,45,0,245,0,176,0,129,0,30,0,178,0,241,0,0,0,128,0,23,0,0,0,0,0,141,0,220,0,0,0,23,0,137,0,152,0,139,0,78,0,213,0,40,0,181,0,190,0,10,0,130,0,246,0,0,0,102,0,0,0,205,0,205,0,148,0,4,0,228,0,23,0,37,0,19,0,110,0,178,0,255,0,134,0,46,0,141,0,155,0,60,0,0,0,103,0,237,0,105,0,80,0,106,0,252,0,12,0,31,0);
signal scenario_full  : scenario_type := (139,31,22,31,34,31,110,31,167,31,210,31,38,31,238,31,95,31,95,30,95,29,178,31,26,31,144,31,144,30,144,29,135,31,250,31,250,30,228,31,228,30,88,31,136,31,238,31,93,31,94,31,146,31,135,31,13,31,13,30,152,31,236,31,236,30,236,29,187,31,187,30,55,31,9,31,163,31,168,31,47,31,47,30,142,31,150,31,224,31,94,31,75,31,90,31,58,31,108,31,190,31,190,30,190,29,56,31,56,30,27,31,26,31,211,31,112,31,189,31,144,31,65,31,207,31,252,31,110,31,102,31,10,31,218,31,218,30,126,31,255,31,88,31,181,31,75,31,30,31,30,30,248,31,185,31,92,31,92,30,92,29,212,31,212,30,212,29,28,31,226,31,253,31,35,31,140,31,15,31,163,31,54,31,141,31,183,31,46,31,207,31,24,31,24,30,230,31,246,31,72,31,71,31,102,31,69,31,125,31,125,30,129,31,226,31,147,31,248,31,203,31,203,30,150,31,144,31,144,30,217,31,160,31,178,31,111,31,111,30,111,29,32,31,198,31,198,30,122,31,163,31,163,30,123,31,123,30,123,29,232,31,232,30,232,29,232,28,18,31,89,31,190,31,72,31,73,31,73,30,248,31,211,31,173,31,154,31,159,31,121,31,162,31,162,30,149,31,127,31,127,30,17,31,131,31,227,31,227,30,164,31,29,31,15,31,48,31,48,30,48,29,255,31,208,31,219,31,216,31,216,30,65,31,124,31,124,30,230,31,124,31,245,31,103,31,131,31,252,31,22,31,27,31,132,31,88,31,88,30,88,29,88,28,88,27,64,31,64,30,130,31,34,31,98,31,197,31,25,31,81,31,142,31,201,31,168,31,246,31,246,30,213,31,213,30,213,29,15,31,15,30,155,31,175,31,175,30,83,31,68,31,33,31,69,31,191,31,42,31,192,31,192,30,45,31,38,31,38,30,146,31,253,31,29,31,90,31,233,31,224,31,44,31,209,31,75,31,25,31,141,31,122,31,45,31,142,31,142,30,27,31,154,31,135,31,135,30,101,31,230,31,230,30,242,31,6,31,172,31,172,30,172,29,50,31,243,31,214,31,119,31,27,31,62,31,3,31,114,31,144,31,98,31,126,31,197,31,81,31,95,31,45,31,245,31,176,31,129,31,30,31,178,31,241,31,241,30,128,31,23,31,23,30,23,29,141,31,220,31,220,30,23,31,137,31,152,31,139,31,78,31,213,31,40,31,181,31,190,31,10,31,130,31,246,31,246,30,102,31,102,30,205,31,205,31,148,31,4,31,228,31,23,31,37,31,19,31,110,31,178,31,255,31,134,31,46,31,141,31,155,31,60,31,60,30,103,31,237,31,105,31,80,31,106,31,252,31,12,31,31,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
