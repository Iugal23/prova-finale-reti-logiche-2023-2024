-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_453 is
end project_tb_453;

architecture project_tb_arch_453 of project_tb_453 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 930;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (68,0,211,0,0,0,0,0,0,0,0,0,141,0,0,0,0,0,0,0,0,0,61,0,92,0,83,0,212,0,0,0,88,0,0,0,0,0,108,0,68,0,65,0,0,0,210,0,227,0,54,0,50,0,241,0,53,0,57,0,90,0,61,0,50,0,0,0,0,0,179,0,0,0,0,0,159,0,20,0,167,0,137,0,68,0,0,0,87,0,51,0,60,0,0,0,150,0,59,0,141,0,59,0,149,0,0,0,111,0,201,0,0,0,0,0,37,0,229,0,51,0,107,0,36,0,244,0,32,0,0,0,28,0,38,0,0,0,167,0,5,0,39,0,215,0,198,0,184,0,0,0,0,0,24,0,255,0,39,0,108,0,42,0,110,0,119,0,105,0,119,0,253,0,190,0,32,0,0,0,0,0,219,0,43,0,199,0,167,0,78,0,73,0,0,0,59,0,0,0,0,0,48,0,226,0,130,0,5,0,167,0,251,0,142,0,202,0,0,0,148,0,188,0,155,0,37,0,215,0,43,0,0,0,3,0,176,0,113,0,7,0,83,0,0,0,54,0,0,0,243,0,0,0,1,0,62,0,148,0,165,0,175,0,0,0,190,0,7,0,215,0,32,0,30,0,205,0,148,0,83,0,53,0,167,0,8,0,51,0,82,0,131,0,243,0,43,0,24,0,210,0,244,0,24,0,165,0,0,0,0,0,0,0,0,0,208,0,130,0,70,0,22,0,112,0,137,0,174,0,235,0,106,0,0,0,189,0,161,0,185,0,202,0,25,0,104,0,100,0,91,0,217,0,101,0,0,0,219,0,97,0,99,0,227,0,79,0,65,0,98,0,160,0,131,0,21,0,0,0,0,0,145,0,162,0,0,0,0,0,20,0,232,0,201,0,118,0,0,0,199,0,30,0,219,0,110,0,213,0,158,0,122,0,163,0,114,0,41,0,0,0,230,0,0,0,0,0,208,0,0,0,221,0,29,0,235,0,3,0,238,0,125,0,0,0,0,0,0,0,161,0,27,0,63,0,248,0,150,0,74,0,139,0,108,0,0,0,54,0,50,0,104,0,0,0,55,0,158,0,221,0,48,0,217,0,218,0,28,0,249,0,205,0,90,0,239,0,59,0,193,0,0,0,79,0,0,0,0,0,249,0,70,0,0,0,177,0,69,0,161,0,83,0,0,0,117,0,0,0,82,0,247,0,96,0,75,0,203,0,55,0,50,0,0,0,0,0,253,0,117,0,209,0,105,0,115,0,176,0,164,0,0,0,0,0,244,0,110,0,34,0,0,0,86,0,132,0,84,0,0,0,48,0,149,0,1,0,132,0,151,0,0,0,204,0,0,0,0,0,194,0,242,0,200,0,113,0,153,0,0,0,0,0,0,0,11,0,134,0,101,0,221,0,0,0,99,0,0,0,143,0,38,0,0,0,0,0,94,0,88,0,0,0,0,0,218,0,138,0,231,0,60,0,87,0,230,0,0,0,145,0,166,0,0,0,0,0,229,0,154,0,153,0,210,0,87,0,231,0,110,0,180,0,210,0,149,0,17,0,147,0,0,0,63,0,197,0,145,0,0,0,129,0,1,0,51,0,67,0,0,0,196,0,164,0,43,0,19,0,16,0,30,0,222,0,254,0,245,0,146,0,177,0,147,0,82,0,80,0,51,0,0,0,34,0,221,0,106,0,220,0,42,0,162,0,1,0,41,0,202,0,144,0,77,0,85,0,83,0,0,0,138,0,219,0,0,0,0,0,254,0,140,0,159,0,224,0,0,0,229,0,47,0,0,0,31,0,34,0,141,0,114,0,0,0,63,0,130,0,83,0,54,0,48,0,132,0,214,0,164,0,0,0,118,0,0,0,27,0,250,0,0,0,139,0,109,0,0,0,18,0,16,0,0,0,0,0,24,0,214,0,0,0,13,0,0,0,163,0,145,0,44,0,0,0,40,0,191,0,58,0,153,0,147,0,107,0,0,0,0,0,0,0,162,0,207,0,129,0,50,0,196,0,59,0,37,0,2,0,88,0,10,0,253,0,0,0,121,0,5,0,20,0,31,0,150,0,36,0,124,0,0,0,238,0,103,0,136,0,0,0,140,0,0,0,0,0,0,0,151,0,0,0,26,0,226,0,255,0,0,0,94,0,119,0,236,0,0,0,0,0,221,0,63,0,18,0,35,0,0,0,159,0,94,0,176,0,0,0,193,0,96,0,16,0,56,0,129,0,0,0,0,0,23,0,145,0,0,0,0,0,135,0,0,0,231,0,93,0,68,0,0,0,113,0,156,0,0,0,62,0,46,0,0,0,248,0,92,0,0,0,41,0,253,0,64,0,13,0,56,0,163,0,135,0,0,0,165,0,204,0,193,0,0,0,14,0,48,0,129,0,212,0,172,0,25,0,0,0,51,0,237,0,25,0,208,0,211,0,107,0,241,0,57,0,83,0,45,0,8,0,24,0,0,0,28,0,64,0,0,0,24,0,253,0,0,0,200,0,82,0,0,0,142,0,36,0,0,0,139,0,130,0,0,0,198,0,209,0,52,0,140,0,49,0,246,0,0,0,229,0,29,0,133,0,31,0,137,0,99,0,87,0,233,0,11,0,250,0,241,0,11,0,195,0,26,0,90,0,195,0,173,0,44,0,0,0,0,0,155,0,20,0,224,0,128,0,72,0,187,0,214,0,198,0,103,0,0,0,77,0,69,0,159,0,140,0,0,0,83,0,18,0,49,0,156,0,189,0,173,0,31,0,21,0,0,0,0,0,241,0,156,0,0,0,57,0,162,0,97,0,0,0,255,0,73,0,0,0,54,0,147,0,152,0,221,0,243,0,115,0,37,0,40,0,213,0,69,0,156,0,0,0,61,0,99,0,116,0,0,0,0,0,56,0,251,0,68,0,8,0,84,0,73,0,0,0,212,0,111,0,70,0,189,0,0,0,111,0,148,0,202,0,62,0,0,0,49,0,135,0,0,0,0,0,228,0,217,0,0,0,173,0,39,0,78,0,0,0,0,0,12,0,148,0,0,0,45,0,145,0,232,0,0,0,39,0,238,0,255,0,62,0,170,0,170,0,48,0,67,0,60,0,224,0,198,0,251,0,7,0,0,0,0,0,102,0,0,0,113,0,52,0,240,0,137,0,252,0,192,0,92,0,198,0,167,0,13,0,132,0,0,0,110,0,234,0,68,0,19,0,93,0,233,0,194,0,87,0,225,0,0,0,155,0,0,0,205,0,0,0,168,0,135,0,56,0,117,0,0,0,207,0,145,0,81,0,50,0,0,0,149,0,215,0,243,0,232,0,24,0,14,0,0,0,0,0,175,0,54,0,197,0,0,0,214,0,19,0,147,0,0,0,99,0,2,0,22,0,0,0,235,0,149,0,16,0,0,0,93,0,49,0,161,0,230,0,0,0,60,0,0,0,184,0,168,0,0,0,0,0,17,0,187,0,0,0,0,0,117,0,108,0,0,0,151,0,160,0,147,0,185,0,0,0,206,0,31,0,46,0,0,0,221,0,0,0,149,0,143,0,0,0,1,0,83,0,0,0,232,0,204,0,0,0,218,0,202,0,39,0,0,0,242,0,120,0,195,0,63,0,232,0,27,0,0,0,238,0,199,0,131,0,246,0,0,0,131,0,190,0,157,0,61,0,10,0,57,0,223,0,225,0,226,0,67,0,0,0,0,0,203,0,200,0,107,0,64,0,137,0,21,0,71,0,114,0,175,0,194,0,0,0,127,0,211,0,113,0,80,0,105,0,0,0,22,0,185,0,67,0,180,0,0,0,9,0,28,0,10,0,90,0,233,0,48,0,31,0,215,0,175,0,251,0,135,0,180,0,102,0,48,0,226,0,74,0,83,0,42,0,6,0,0,0,152,0,80,0,17,0,244,0,187,0,82,0,5,0,218,0,215,0,219,0,38,0,0,0,1,0,48,0,241,0,168,0,0,0,33,0,0,0,3,0,219,0,236,0,136,0,39,0,170,0,81,0,0,0,163,0,1,0,88,0,23,0,101,0,89,0,57,0,176,0,226,0,9,0,0,0,240,0,38,0,14,0,181,0,94,0,22,0,236,0,155,0,0,0,0,0,192,0,252,0,47,0,172,0,197,0,230,0,17,0,0,0,60,0,41,0,46,0,149,0,0,0,8,0,44,0,191,0,81,0,0,0,0,0);
signal scenario_full  : scenario_type := (68,31,211,31,211,30,211,29,211,28,211,27,141,31,141,30,141,29,141,28,141,27,61,31,92,31,83,31,212,31,212,30,88,31,88,30,88,29,108,31,68,31,65,31,65,30,210,31,227,31,54,31,50,31,241,31,53,31,57,31,90,31,61,31,50,31,50,30,50,29,179,31,179,30,179,29,159,31,20,31,167,31,137,31,68,31,68,30,87,31,51,31,60,31,60,30,150,31,59,31,141,31,59,31,149,31,149,30,111,31,201,31,201,30,201,29,37,31,229,31,51,31,107,31,36,31,244,31,32,31,32,30,28,31,38,31,38,30,167,31,5,31,39,31,215,31,198,31,184,31,184,30,184,29,24,31,255,31,39,31,108,31,42,31,110,31,119,31,105,31,119,31,253,31,190,31,32,31,32,30,32,29,219,31,43,31,199,31,167,31,78,31,73,31,73,30,59,31,59,30,59,29,48,31,226,31,130,31,5,31,167,31,251,31,142,31,202,31,202,30,148,31,188,31,155,31,37,31,215,31,43,31,43,30,3,31,176,31,113,31,7,31,83,31,83,30,54,31,54,30,243,31,243,30,1,31,62,31,148,31,165,31,175,31,175,30,190,31,7,31,215,31,32,31,30,31,205,31,148,31,83,31,53,31,167,31,8,31,51,31,82,31,131,31,243,31,43,31,24,31,210,31,244,31,24,31,165,31,165,30,165,29,165,28,165,27,208,31,130,31,70,31,22,31,112,31,137,31,174,31,235,31,106,31,106,30,189,31,161,31,185,31,202,31,25,31,104,31,100,31,91,31,217,31,101,31,101,30,219,31,97,31,99,31,227,31,79,31,65,31,98,31,160,31,131,31,21,31,21,30,21,29,145,31,162,31,162,30,162,29,20,31,232,31,201,31,118,31,118,30,199,31,30,31,219,31,110,31,213,31,158,31,122,31,163,31,114,31,41,31,41,30,230,31,230,30,230,29,208,31,208,30,221,31,29,31,235,31,3,31,238,31,125,31,125,30,125,29,125,28,161,31,27,31,63,31,248,31,150,31,74,31,139,31,108,31,108,30,54,31,50,31,104,31,104,30,55,31,158,31,221,31,48,31,217,31,218,31,28,31,249,31,205,31,90,31,239,31,59,31,193,31,193,30,79,31,79,30,79,29,249,31,70,31,70,30,177,31,69,31,161,31,83,31,83,30,117,31,117,30,82,31,247,31,96,31,75,31,203,31,55,31,50,31,50,30,50,29,253,31,117,31,209,31,105,31,115,31,176,31,164,31,164,30,164,29,244,31,110,31,34,31,34,30,86,31,132,31,84,31,84,30,48,31,149,31,1,31,132,31,151,31,151,30,204,31,204,30,204,29,194,31,242,31,200,31,113,31,153,31,153,30,153,29,153,28,11,31,134,31,101,31,221,31,221,30,99,31,99,30,143,31,38,31,38,30,38,29,94,31,88,31,88,30,88,29,218,31,138,31,231,31,60,31,87,31,230,31,230,30,145,31,166,31,166,30,166,29,229,31,154,31,153,31,210,31,87,31,231,31,110,31,180,31,210,31,149,31,17,31,147,31,147,30,63,31,197,31,145,31,145,30,129,31,1,31,51,31,67,31,67,30,196,31,164,31,43,31,19,31,16,31,30,31,222,31,254,31,245,31,146,31,177,31,147,31,82,31,80,31,51,31,51,30,34,31,221,31,106,31,220,31,42,31,162,31,1,31,41,31,202,31,144,31,77,31,85,31,83,31,83,30,138,31,219,31,219,30,219,29,254,31,140,31,159,31,224,31,224,30,229,31,47,31,47,30,31,31,34,31,141,31,114,31,114,30,63,31,130,31,83,31,54,31,48,31,132,31,214,31,164,31,164,30,118,31,118,30,27,31,250,31,250,30,139,31,109,31,109,30,18,31,16,31,16,30,16,29,24,31,214,31,214,30,13,31,13,30,163,31,145,31,44,31,44,30,40,31,191,31,58,31,153,31,147,31,107,31,107,30,107,29,107,28,162,31,207,31,129,31,50,31,196,31,59,31,37,31,2,31,88,31,10,31,253,31,253,30,121,31,5,31,20,31,31,31,150,31,36,31,124,31,124,30,238,31,103,31,136,31,136,30,140,31,140,30,140,29,140,28,151,31,151,30,26,31,226,31,255,31,255,30,94,31,119,31,236,31,236,30,236,29,221,31,63,31,18,31,35,31,35,30,159,31,94,31,176,31,176,30,193,31,96,31,16,31,56,31,129,31,129,30,129,29,23,31,145,31,145,30,145,29,135,31,135,30,231,31,93,31,68,31,68,30,113,31,156,31,156,30,62,31,46,31,46,30,248,31,92,31,92,30,41,31,253,31,64,31,13,31,56,31,163,31,135,31,135,30,165,31,204,31,193,31,193,30,14,31,48,31,129,31,212,31,172,31,25,31,25,30,51,31,237,31,25,31,208,31,211,31,107,31,241,31,57,31,83,31,45,31,8,31,24,31,24,30,28,31,64,31,64,30,24,31,253,31,253,30,200,31,82,31,82,30,142,31,36,31,36,30,139,31,130,31,130,30,198,31,209,31,52,31,140,31,49,31,246,31,246,30,229,31,29,31,133,31,31,31,137,31,99,31,87,31,233,31,11,31,250,31,241,31,11,31,195,31,26,31,90,31,195,31,173,31,44,31,44,30,44,29,155,31,20,31,224,31,128,31,72,31,187,31,214,31,198,31,103,31,103,30,77,31,69,31,159,31,140,31,140,30,83,31,18,31,49,31,156,31,189,31,173,31,31,31,21,31,21,30,21,29,241,31,156,31,156,30,57,31,162,31,97,31,97,30,255,31,73,31,73,30,54,31,147,31,152,31,221,31,243,31,115,31,37,31,40,31,213,31,69,31,156,31,156,30,61,31,99,31,116,31,116,30,116,29,56,31,251,31,68,31,8,31,84,31,73,31,73,30,212,31,111,31,70,31,189,31,189,30,111,31,148,31,202,31,62,31,62,30,49,31,135,31,135,30,135,29,228,31,217,31,217,30,173,31,39,31,78,31,78,30,78,29,12,31,148,31,148,30,45,31,145,31,232,31,232,30,39,31,238,31,255,31,62,31,170,31,170,31,48,31,67,31,60,31,224,31,198,31,251,31,7,31,7,30,7,29,102,31,102,30,113,31,52,31,240,31,137,31,252,31,192,31,92,31,198,31,167,31,13,31,132,31,132,30,110,31,234,31,68,31,19,31,93,31,233,31,194,31,87,31,225,31,225,30,155,31,155,30,205,31,205,30,168,31,135,31,56,31,117,31,117,30,207,31,145,31,81,31,50,31,50,30,149,31,215,31,243,31,232,31,24,31,14,31,14,30,14,29,175,31,54,31,197,31,197,30,214,31,19,31,147,31,147,30,99,31,2,31,22,31,22,30,235,31,149,31,16,31,16,30,93,31,49,31,161,31,230,31,230,30,60,31,60,30,184,31,168,31,168,30,168,29,17,31,187,31,187,30,187,29,117,31,108,31,108,30,151,31,160,31,147,31,185,31,185,30,206,31,31,31,46,31,46,30,221,31,221,30,149,31,143,31,143,30,1,31,83,31,83,30,232,31,204,31,204,30,218,31,202,31,39,31,39,30,242,31,120,31,195,31,63,31,232,31,27,31,27,30,238,31,199,31,131,31,246,31,246,30,131,31,190,31,157,31,61,31,10,31,57,31,223,31,225,31,226,31,67,31,67,30,67,29,203,31,200,31,107,31,64,31,137,31,21,31,71,31,114,31,175,31,194,31,194,30,127,31,211,31,113,31,80,31,105,31,105,30,22,31,185,31,67,31,180,31,180,30,9,31,28,31,10,31,90,31,233,31,48,31,31,31,215,31,175,31,251,31,135,31,180,31,102,31,48,31,226,31,74,31,83,31,42,31,6,31,6,30,152,31,80,31,17,31,244,31,187,31,82,31,5,31,218,31,215,31,219,31,38,31,38,30,1,31,48,31,241,31,168,31,168,30,33,31,33,30,3,31,219,31,236,31,136,31,39,31,170,31,81,31,81,30,163,31,1,31,88,31,23,31,101,31,89,31,57,31,176,31,226,31,9,31,9,30,240,31,38,31,14,31,181,31,94,31,22,31,236,31,155,31,155,30,155,29,192,31,252,31,47,31,172,31,197,31,230,31,17,31,17,30,60,31,41,31,46,31,149,31,149,30,8,31,44,31,191,31,81,31,81,30,81,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
