-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 853;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (237,0,0,0,48,0,35,0,25,0,190,0,244,0,0,0,105,0,53,0,0,0,50,0,121,0,207,0,165,0,189,0,240,0,62,0,242,0,71,0,244,0,69,0,96,0,74,0,252,0,130,0,70,0,19,0,65,0,0,0,47,0,125,0,0,0,85,0,202,0,0,0,190,0,26,0,43,0,118,0,78,0,35,0,160,0,212,0,89,0,12,0,0,0,2,0,66,0,252,0,0,0,172,0,202,0,208,0,60,0,191,0,240,0,22,0,38,0,0,0,176,0,22,0,235,0,86,0,69,0,119,0,0,0,0,0,0,0,194,0,241,0,173,0,210,0,0,0,0,0,72,0,213,0,209,0,125,0,5,0,0,0,152,0,0,0,106,0,239,0,186,0,154,0,56,0,117,0,186,0,38,0,145,0,0,0,171,0,251,0,198,0,188,0,20,0,147,0,128,0,63,0,0,0,14,0,0,0,0,0,186,0,100,0,161,0,224,0,135,0,157,0,107,0,40,0,162,0,144,0,41,0,187,0,101,0,216,0,0,0,28,0,20,0,165,0,101,0,75,0,44,0,0,0,180,0,250,0,22,0,157,0,175,0,99,0,79,0,238,0,197,0,105,0,0,0,160,0,159,0,12,0,63,0,207,0,0,0,0,0,0,0,174,0,65,0,79,0,24,0,179,0,48,0,50,0,219,0,41,0,131,0,141,0,242,0,105,0,0,0,90,0,0,0,0,0,0,0,0,0,245,0,0,0,0,0,213,0,250,0,199,0,89,0,6,0,180,0,48,0,162,0,21,0,246,0,9,0,178,0,165,0,223,0,0,0,41,0,0,0,140,0,0,0,117,0,0,0,0,0,177,0,15,0,159,0,168,0,210,0,165,0,174,0,37,0,158,0,0,0,209,0,0,0,0,0,23,0,102,0,8,0,86,0,15,0,0,0,147,0,12,0,183,0,0,0,127,0,15,0,0,0,173,0,217,0,0,0,24,0,0,0,119,0,169,0,73,0,129,0,138,0,0,0,178,0,16,0,176,0,141,0,35,0,233,0,0,0,58,0,0,0,147,0,86,0,84,0,98,0,0,0,40,0,254,0,149,0,0,0,78,0,117,0,129,0,105,0,79,0,114,0,0,0,234,0,29,0,36,0,177,0,0,0,8,0,38,0,110,0,188,0,0,0,64,0,23,0,242,0,154,0,39,0,181,0,227,0,0,0,28,0,0,0,49,0,119,0,102,0,28,0,255,0,69,0,64,0,197,0,181,0,169,0,102,0,0,0,54,0,0,0,249,0,184,0,79,0,160,0,0,0,163,0,0,0,28,0,106,0,86,0,108,0,0,0,7,0,68,0,36,0,226,0,61,0,0,0,167,0,110,0,136,0,109,0,146,0,91,0,221,0,115,0,113,0,127,0,22,0,121,0,0,0,0,0,244,0,0,0,28,0,0,0,100,0,0,0,0,0,32,0,216,0,0,0,0,0,0,0,0,0,107,0,21,0,81,0,0,0,37,0,0,0,245,0,173,0,67,0,25,0,0,0,122,0,26,0,171,0,29,0,17,0,79,0,181,0,0,0,32,0,0,0,167,0,90,0,210,0,91,0,0,0,0,0,218,0,195,0,224,0,26,0,57,0,99,0,70,0,0,0,41,0,128,0,15,0,213,0,138,0,214,0,152,0,200,0,54,0,100,0,19,0,5,0,167,0,169,0,147,0,142,0,243,0,131,0,0,0,103,0,0,0,121,0,156,0,50,0,96,0,217,0,36,0,0,0,231,0,109,0,246,0,58,0,0,0,147,0,162,0,230,0,188,0,0,0,91,0,242,0,39,0,6,0,77,0,242,0,79,0,0,0,19,0,106,0,108,0,0,0,135,0,213,0,45,0,193,0,28,0,195,0,37,0,0,0,22,0,0,0,254,0,59,0,185,0,0,0,82,0,213,0,5,0,28,0,212,0,82,0,17,0,0,0,0,0,107,0,53,0,158,0,17,0,231,0,203,0,171,0,29,0,251,0,205,0,146,0,0,0,254,0,127,0,0,0,231,0,42,0,16,0,0,0,144,0,181,0,0,0,55,0,122,0,179,0,102,0,171,0,0,0,82,0,121,0,2,0,0,0,69,0,0,0,15,0,219,0,141,0,127,0,0,0,142,0,24,0,63,0,81,0,0,0,224,0,220,0,51,0,110,0,95,0,231,0,33,0,79,0,203,0,67,0,102,0,9,0,178,0,0,0,192,0,138,0,179,0,213,0,58,0,98,0,178,0,183,0,21,0,105,0,0,0,5,0,5,0,161,0,8,0,0,0,178,0,173,0,86,0,73,0,249,0,194,0,219,0,86,0,36,0,35,0,40,0,0,0,82,0,160,0,229,0,78,0,154,0,69,0,150,0,131,0,28,0,167,0,75,0,174,0,200,0,54,0,112,0,247,0,0,0,76,0,9,0,27,0,12,0,22,0,0,0,128,0,32,0,44,0,212,0,156,0,126,0,104,0,0,0,0,0,52,0,0,0,59,0,93,0,223,0,34,0,105,0,62,0,114,0,6,0,45,0,0,0,158,0,168,0,92,0,0,0,170,0,212,0,134,0,241,0,0,0,23,0,87,0,132,0,0,0,51,0,28,0,29,0,252,0,93,0,202,0,0,0,69,0,0,0,15,0,0,0,0,0,0,0,22,0,209,0,46,0,156,0,0,0,205,0,0,0,63,0,38,0,44,0,238,0,150,0,0,0,83,0,0,0,121,0,131,0,0,0,57,0,85,0,213,0,233,0,0,0,97,0,141,0,186,0,5,0,0,0,0,0,236,0,0,0,234,0,0,0,83,0,0,0,251,0,235,0,33,0,56,0,168,0,248,0,104,0,0,0,50,0,0,0,28,0,200,0,154,0,0,0,131,0,218,0,53,0,0,0,172,0,74,0,0,0,187,0,0,0,110,0,0,0,93,0,109,0,131,0,7,0,197,0,234,0,140,0,123,0,112,0,128,0,166,0,0,0,219,0,123,0,49,0,0,0,0,0,242,0,178,0,110,0,0,0,83,0,45,0,208,0,131,0,57,0,241,0,53,0,47,0,28,0,205,0,0,0,144,0,116,0,113,0,191,0,29,0,77,0,2,0,218,0,144,0,103,0,56,0,38,0,167,0,16,0,174,0,194,0,0,0,250,0,96,0,63,0,108,0,2,0,138,0,221,0,204,0,0,0,0,0,234,0,81,0,209,0,174,0,18,0,236,0,224,0,0,0,204,0,64,0,156,0,0,0,95,0,24,0,0,0,139,0,0,0,43,0,0,0,149,0,81,0,226,0,12,0,0,0,173,0,77,0,246,0,152,0,0,0,239,0,125,0,0,0,44,0,0,0,159,0,0,0,36,0,65,0,22,0,96,0,0,0,155,0,0,0,115,0,34,0,56,0,45,0,26,0,159,0,147,0,101,0,199,0,0,0,46,0,207,0,138,0,211,0,82,0,92,0,156,0,166,0,0,0,113,0,176,0,8,0,30,0,0,0,212,0,0,0,191,0,138,0,195,0,145,0,105,0,82,0,0,0,132,0,222,0,12,0,109,0,38,0,0,0,14,0,96,0,224,0,26,0,0,0,0,0,89,0,136,0,159,0,31,0,98,0,46,0,19,0,236,0,152,0,90,0,114,0,0,0,142,0,0,0,96,0,237,0,229,0,175,0,173,0,30,0,0,0,0,0,202,0,57,0,232,0,139,0,213,0,202,0,224,0,198,0,68,0,28,0,0,0,105,0,0,0,225,0,129,0,9,0,168,0,147,0,0,0,95,0,0,0,252,0,63,0,52,0,0,0,162,0,202,0,199,0,7,0);
signal scenario_full  : scenario_type := (237,31,237,30,48,31,35,31,25,31,190,31,244,31,244,30,105,31,53,31,53,30,50,31,121,31,207,31,165,31,189,31,240,31,62,31,242,31,71,31,244,31,69,31,96,31,74,31,252,31,130,31,70,31,19,31,65,31,65,30,47,31,125,31,125,30,85,31,202,31,202,30,190,31,26,31,43,31,118,31,78,31,35,31,160,31,212,31,89,31,12,31,12,30,2,31,66,31,252,31,252,30,172,31,202,31,208,31,60,31,191,31,240,31,22,31,38,31,38,30,176,31,22,31,235,31,86,31,69,31,119,31,119,30,119,29,119,28,194,31,241,31,173,31,210,31,210,30,210,29,72,31,213,31,209,31,125,31,5,31,5,30,152,31,152,30,106,31,239,31,186,31,154,31,56,31,117,31,186,31,38,31,145,31,145,30,171,31,251,31,198,31,188,31,20,31,147,31,128,31,63,31,63,30,14,31,14,30,14,29,186,31,100,31,161,31,224,31,135,31,157,31,107,31,40,31,162,31,144,31,41,31,187,31,101,31,216,31,216,30,28,31,20,31,165,31,101,31,75,31,44,31,44,30,180,31,250,31,22,31,157,31,175,31,99,31,79,31,238,31,197,31,105,31,105,30,160,31,159,31,12,31,63,31,207,31,207,30,207,29,207,28,174,31,65,31,79,31,24,31,179,31,48,31,50,31,219,31,41,31,131,31,141,31,242,31,105,31,105,30,90,31,90,30,90,29,90,28,90,27,245,31,245,30,245,29,213,31,250,31,199,31,89,31,6,31,180,31,48,31,162,31,21,31,246,31,9,31,178,31,165,31,223,31,223,30,41,31,41,30,140,31,140,30,117,31,117,30,117,29,177,31,15,31,159,31,168,31,210,31,165,31,174,31,37,31,158,31,158,30,209,31,209,30,209,29,23,31,102,31,8,31,86,31,15,31,15,30,147,31,12,31,183,31,183,30,127,31,15,31,15,30,173,31,217,31,217,30,24,31,24,30,119,31,169,31,73,31,129,31,138,31,138,30,178,31,16,31,176,31,141,31,35,31,233,31,233,30,58,31,58,30,147,31,86,31,84,31,98,31,98,30,40,31,254,31,149,31,149,30,78,31,117,31,129,31,105,31,79,31,114,31,114,30,234,31,29,31,36,31,177,31,177,30,8,31,38,31,110,31,188,31,188,30,64,31,23,31,242,31,154,31,39,31,181,31,227,31,227,30,28,31,28,30,49,31,119,31,102,31,28,31,255,31,69,31,64,31,197,31,181,31,169,31,102,31,102,30,54,31,54,30,249,31,184,31,79,31,160,31,160,30,163,31,163,30,28,31,106,31,86,31,108,31,108,30,7,31,68,31,36,31,226,31,61,31,61,30,167,31,110,31,136,31,109,31,146,31,91,31,221,31,115,31,113,31,127,31,22,31,121,31,121,30,121,29,244,31,244,30,28,31,28,30,100,31,100,30,100,29,32,31,216,31,216,30,216,29,216,28,216,27,107,31,21,31,81,31,81,30,37,31,37,30,245,31,173,31,67,31,25,31,25,30,122,31,26,31,171,31,29,31,17,31,79,31,181,31,181,30,32,31,32,30,167,31,90,31,210,31,91,31,91,30,91,29,218,31,195,31,224,31,26,31,57,31,99,31,70,31,70,30,41,31,128,31,15,31,213,31,138,31,214,31,152,31,200,31,54,31,100,31,19,31,5,31,167,31,169,31,147,31,142,31,243,31,131,31,131,30,103,31,103,30,121,31,156,31,50,31,96,31,217,31,36,31,36,30,231,31,109,31,246,31,58,31,58,30,147,31,162,31,230,31,188,31,188,30,91,31,242,31,39,31,6,31,77,31,242,31,79,31,79,30,19,31,106,31,108,31,108,30,135,31,213,31,45,31,193,31,28,31,195,31,37,31,37,30,22,31,22,30,254,31,59,31,185,31,185,30,82,31,213,31,5,31,28,31,212,31,82,31,17,31,17,30,17,29,107,31,53,31,158,31,17,31,231,31,203,31,171,31,29,31,251,31,205,31,146,31,146,30,254,31,127,31,127,30,231,31,42,31,16,31,16,30,144,31,181,31,181,30,55,31,122,31,179,31,102,31,171,31,171,30,82,31,121,31,2,31,2,30,69,31,69,30,15,31,219,31,141,31,127,31,127,30,142,31,24,31,63,31,81,31,81,30,224,31,220,31,51,31,110,31,95,31,231,31,33,31,79,31,203,31,67,31,102,31,9,31,178,31,178,30,192,31,138,31,179,31,213,31,58,31,98,31,178,31,183,31,21,31,105,31,105,30,5,31,5,31,161,31,8,31,8,30,178,31,173,31,86,31,73,31,249,31,194,31,219,31,86,31,36,31,35,31,40,31,40,30,82,31,160,31,229,31,78,31,154,31,69,31,150,31,131,31,28,31,167,31,75,31,174,31,200,31,54,31,112,31,247,31,247,30,76,31,9,31,27,31,12,31,22,31,22,30,128,31,32,31,44,31,212,31,156,31,126,31,104,31,104,30,104,29,52,31,52,30,59,31,93,31,223,31,34,31,105,31,62,31,114,31,6,31,45,31,45,30,158,31,168,31,92,31,92,30,170,31,212,31,134,31,241,31,241,30,23,31,87,31,132,31,132,30,51,31,28,31,29,31,252,31,93,31,202,31,202,30,69,31,69,30,15,31,15,30,15,29,15,28,22,31,209,31,46,31,156,31,156,30,205,31,205,30,63,31,38,31,44,31,238,31,150,31,150,30,83,31,83,30,121,31,131,31,131,30,57,31,85,31,213,31,233,31,233,30,97,31,141,31,186,31,5,31,5,30,5,29,236,31,236,30,234,31,234,30,83,31,83,30,251,31,235,31,33,31,56,31,168,31,248,31,104,31,104,30,50,31,50,30,28,31,200,31,154,31,154,30,131,31,218,31,53,31,53,30,172,31,74,31,74,30,187,31,187,30,110,31,110,30,93,31,109,31,131,31,7,31,197,31,234,31,140,31,123,31,112,31,128,31,166,31,166,30,219,31,123,31,49,31,49,30,49,29,242,31,178,31,110,31,110,30,83,31,45,31,208,31,131,31,57,31,241,31,53,31,47,31,28,31,205,31,205,30,144,31,116,31,113,31,191,31,29,31,77,31,2,31,218,31,144,31,103,31,56,31,38,31,167,31,16,31,174,31,194,31,194,30,250,31,96,31,63,31,108,31,2,31,138,31,221,31,204,31,204,30,204,29,234,31,81,31,209,31,174,31,18,31,236,31,224,31,224,30,204,31,64,31,156,31,156,30,95,31,24,31,24,30,139,31,139,30,43,31,43,30,149,31,81,31,226,31,12,31,12,30,173,31,77,31,246,31,152,31,152,30,239,31,125,31,125,30,44,31,44,30,159,31,159,30,36,31,65,31,22,31,96,31,96,30,155,31,155,30,115,31,34,31,56,31,45,31,26,31,159,31,147,31,101,31,199,31,199,30,46,31,207,31,138,31,211,31,82,31,92,31,156,31,166,31,166,30,113,31,176,31,8,31,30,31,30,30,212,31,212,30,191,31,138,31,195,31,145,31,105,31,82,31,82,30,132,31,222,31,12,31,109,31,38,31,38,30,14,31,96,31,224,31,26,31,26,30,26,29,89,31,136,31,159,31,31,31,98,31,46,31,19,31,236,31,152,31,90,31,114,31,114,30,142,31,142,30,96,31,237,31,229,31,175,31,173,31,30,31,30,30,30,29,202,31,57,31,232,31,139,31,213,31,202,31,224,31,198,31,68,31,28,31,28,30,105,31,105,30,225,31,129,31,9,31,168,31,147,31,147,30,95,31,95,30,252,31,63,31,52,31,52,30,162,31,202,31,199,31,7,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
