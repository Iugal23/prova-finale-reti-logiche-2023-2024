-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 660;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,44,0,39,0,109,0,140,0,0,0,0,0,0,0,0,0,59,0,40,0,129,0,171,0,242,0,178,0,10,0,0,0,0,0,0,0,135,0,0,0,217,0,132,0,0,0,38,0,98,0,0,0,40,0,0,0,36,0,149,0,0,0,232,0,41,0,192,0,254,0,60,0,84,0,186,0,254,0,88,0,26,0,66,0,106,0,72,0,0,0,50,0,140,0,0,0,52,0,31,0,43,0,134,0,233,0,0,0,0,0,30,0,81,0,5,0,89,0,203,0,79,0,250,0,0,0,0,0,0,0,0,0,21,0,192,0,58,0,192,0,127,0,228,0,139,0,36,0,18,0,241,0,14,0,0,0,121,0,136,0,238,0,83,0,135,0,33,0,162,0,105,0,0,0,199,0,77,0,71,0,243,0,146,0,0,0,125,0,15,0,99,0,238,0,119,0,49,0,60,0,0,0,219,0,47,0,222,0,157,0,70,0,106,0,9,0,124,0,39,0,207,0,54,0,0,0,106,0,216,0,0,0,0,0,243,0,43,0,0,0,189,0,232,0,128,0,161,0,209,0,0,0,169,0,23,0,105,0,226,0,60,0,89,0,0,0,149,0,233,0,60,0,73,0,0,0,130,0,0,0,14,0,141,0,253,0,32,0,59,0,0,0,176,0,178,0,160,0,132,0,172,0,13,0,217,0,69,0,116,0,94,0,0,0,22,0,217,0,0,0,183,0,180,0,0,0,74,0,124,0,0,0,0,0,45,0,58,0,72,0,38,0,114,0,145,0,21,0,207,0,21,0,236,0,54,0,82,0,148,0,0,0,0,0,24,0,212,0,111,0,202,0,0,0,0,0,25,0,0,0,81,0,116,0,88,0,233,0,0,0,160,0,67,0,0,0,216,0,0,0,166,0,183,0,243,0,107,0,245,0,39,0,75,0,29,0,210,0,13,0,38,0,119,0,224,0,120,0,227,0,191,0,36,0,127,0,150,0,0,0,119,0,255,0,217,0,206,0,18,0,202,0,2,0,191,0,180,0,0,0,85,0,179,0,96,0,0,0,169,0,0,0,162,0,231,0,164,0,100,0,227,0,0,0,93,0,145,0,79,0,95,0,131,0,0,0,204,0,116,0,0,0,66,0,19,0,228,0,17,0,0,0,0,0,102,0,84,0,41,0,8,0,162,0,108,0,196,0,0,0,169,0,39,0,141,0,83,0,57,0,131,0,7,0,179,0,0,0,243,0,116,0,232,0,117,0,2,0,122,0,0,0,51,0,211,0,163,0,108,0,2,0,0,0,0,0,147,0,81,0,72,0,246,0,52,0,45,0,67,0,208,0,137,0,86,0,16,0,0,0,44,0,214,0,155,0,163,0,13,0,234,0,170,0,250,0,0,0,0,0,21,0,210,0,60,0,62,0,22,0,167,0,134,0,95,0,199,0,143,0,238,0,177,0,29,0,97,0,62,0,44,0,0,0,46,0,120,0,53,0,22,0,253,0,0,0,34,0,52,0,0,0,47,0,158,0,20,0,62,0,198,0,79,0,57,0,227,0,26,0,153,0,135,0,0,0,51,0,0,0,56,0,0,0,109,0,0,0,0,0,186,0,0,0,171,0,20,0,159,0,0,0,231,0,140,0,0,0,0,0,85,0,0,0,229,0,0,0,173,0,115,0,223,0,192,0,95,0,37,0,64,0,31,0,68,0,191,0,66,0,4,0,200,0,171,0,164,0,86,0,93,0,201,0,160,0,0,0,72,0,131,0,247,0,180,0,129,0,47,0,121,0,215,0,169,0,0,0,215,0,0,0,58,0,0,0,0,0,144,0,138,0,152,0,204,0,137,0,0,0,185,0,87,0,196,0,195,0,240,0,107,0,85,0,0,0,98,0,0,0,215,0,191,0,0,0,185,0,0,0,0,0,0,0,40,0,163,0,13,0,142,0,0,0,60,0,194,0,215,0,55,0,94,0,239,0,162,0,0,0,61,0,0,0,178,0,85,0,175,0,85,0,40,0,254,0,162,0,221,0,0,0,186,0,207,0,84,0,0,0,0,0,249,0,0,0,175,0,32,0,156,0,141,0,49,0,201,0,107,0,116,0,25,0,5,0,191,0,0,0,62,0,157,0,0,0,0,0,144,0,0,0,129,0,104,0,43,0,34,0,245,0,251,0,11,0,0,0,44,0,158,0,123,0,193,0,118,0,248,0,153,0,90,0,72,0,159,0,0,0,11,0,164,0,31,0,19,0,195,0,51,0,213,0,85,0,236,0,240,0,0,0,0,0,241,0,150,0,254,0,164,0,1,0,105,0,66,0,32,0,131,0,109,0,188,0,44,0,75,0,169,0,199,0,0,0,149,0,130,0,150,0,0,0,213,0,166,0,69,0,0,0,184,0,33,0,187,0,0,0,122,0,12,0,106,0,242,0,102,0,0,0,243,0,30,0,136,0,105,0,23,0,0,0,181,0,0,0,231,0,150,0,0,0,13,0,28,0,102,0,199,0,59,0,205,0,37,0,196,0,187,0,163,0,69,0,206,0,134,0,244,0,3,0,0,0,0,0,202,0,171,0,63,0,168,0,185,0,159,0,2,0,22,0,234,0,35,0,0,0,46,0,173,0,62,0,167,0,189,0,177,0,0,0,63,0,179,0,8,0,233,0,72,0,104,0,45,0,0,0,74,0,0,0,224,0,73,0,37,0,63,0,62,0,97,0,213,0,0,0,0,0,253,0,239,0,239,0,155,0,143,0,248,0,204,0,0,0,0,0,50,0,167,0,0,0,0,0,0,0,199,0,251,0,50,0,126,0,55,0,199,0,169,0,105,0,0,0,236,0,0,0,227,0,178,0,204,0,0,0,48,0,122,0,158,0,205,0,60,0,149,0,26,0,119,0,120,0,0,0,52,0,157,0,159,0,167,0,62,0,0,0,249,0,164,0,158,0,68,0,123,0,219,0,180,0);
signal scenario_full  : scenario_type := (0,0,0,0,44,31,39,31,109,31,140,31,140,30,140,29,140,28,140,27,59,31,40,31,129,31,171,31,242,31,178,31,10,31,10,30,10,29,10,28,135,31,135,30,217,31,132,31,132,30,38,31,98,31,98,30,40,31,40,30,36,31,149,31,149,30,232,31,41,31,192,31,254,31,60,31,84,31,186,31,254,31,88,31,26,31,66,31,106,31,72,31,72,30,50,31,140,31,140,30,52,31,31,31,43,31,134,31,233,31,233,30,233,29,30,31,81,31,5,31,89,31,203,31,79,31,250,31,250,30,250,29,250,28,250,27,21,31,192,31,58,31,192,31,127,31,228,31,139,31,36,31,18,31,241,31,14,31,14,30,121,31,136,31,238,31,83,31,135,31,33,31,162,31,105,31,105,30,199,31,77,31,71,31,243,31,146,31,146,30,125,31,15,31,99,31,238,31,119,31,49,31,60,31,60,30,219,31,47,31,222,31,157,31,70,31,106,31,9,31,124,31,39,31,207,31,54,31,54,30,106,31,216,31,216,30,216,29,243,31,43,31,43,30,189,31,232,31,128,31,161,31,209,31,209,30,169,31,23,31,105,31,226,31,60,31,89,31,89,30,149,31,233,31,60,31,73,31,73,30,130,31,130,30,14,31,141,31,253,31,32,31,59,31,59,30,176,31,178,31,160,31,132,31,172,31,13,31,217,31,69,31,116,31,94,31,94,30,22,31,217,31,217,30,183,31,180,31,180,30,74,31,124,31,124,30,124,29,45,31,58,31,72,31,38,31,114,31,145,31,21,31,207,31,21,31,236,31,54,31,82,31,148,31,148,30,148,29,24,31,212,31,111,31,202,31,202,30,202,29,25,31,25,30,81,31,116,31,88,31,233,31,233,30,160,31,67,31,67,30,216,31,216,30,166,31,183,31,243,31,107,31,245,31,39,31,75,31,29,31,210,31,13,31,38,31,119,31,224,31,120,31,227,31,191,31,36,31,127,31,150,31,150,30,119,31,255,31,217,31,206,31,18,31,202,31,2,31,191,31,180,31,180,30,85,31,179,31,96,31,96,30,169,31,169,30,162,31,231,31,164,31,100,31,227,31,227,30,93,31,145,31,79,31,95,31,131,31,131,30,204,31,116,31,116,30,66,31,19,31,228,31,17,31,17,30,17,29,102,31,84,31,41,31,8,31,162,31,108,31,196,31,196,30,169,31,39,31,141,31,83,31,57,31,131,31,7,31,179,31,179,30,243,31,116,31,232,31,117,31,2,31,122,31,122,30,51,31,211,31,163,31,108,31,2,31,2,30,2,29,147,31,81,31,72,31,246,31,52,31,45,31,67,31,208,31,137,31,86,31,16,31,16,30,44,31,214,31,155,31,163,31,13,31,234,31,170,31,250,31,250,30,250,29,21,31,210,31,60,31,62,31,22,31,167,31,134,31,95,31,199,31,143,31,238,31,177,31,29,31,97,31,62,31,44,31,44,30,46,31,120,31,53,31,22,31,253,31,253,30,34,31,52,31,52,30,47,31,158,31,20,31,62,31,198,31,79,31,57,31,227,31,26,31,153,31,135,31,135,30,51,31,51,30,56,31,56,30,109,31,109,30,109,29,186,31,186,30,171,31,20,31,159,31,159,30,231,31,140,31,140,30,140,29,85,31,85,30,229,31,229,30,173,31,115,31,223,31,192,31,95,31,37,31,64,31,31,31,68,31,191,31,66,31,4,31,200,31,171,31,164,31,86,31,93,31,201,31,160,31,160,30,72,31,131,31,247,31,180,31,129,31,47,31,121,31,215,31,169,31,169,30,215,31,215,30,58,31,58,30,58,29,144,31,138,31,152,31,204,31,137,31,137,30,185,31,87,31,196,31,195,31,240,31,107,31,85,31,85,30,98,31,98,30,215,31,191,31,191,30,185,31,185,30,185,29,185,28,40,31,163,31,13,31,142,31,142,30,60,31,194,31,215,31,55,31,94,31,239,31,162,31,162,30,61,31,61,30,178,31,85,31,175,31,85,31,40,31,254,31,162,31,221,31,221,30,186,31,207,31,84,31,84,30,84,29,249,31,249,30,175,31,32,31,156,31,141,31,49,31,201,31,107,31,116,31,25,31,5,31,191,31,191,30,62,31,157,31,157,30,157,29,144,31,144,30,129,31,104,31,43,31,34,31,245,31,251,31,11,31,11,30,44,31,158,31,123,31,193,31,118,31,248,31,153,31,90,31,72,31,159,31,159,30,11,31,164,31,31,31,19,31,195,31,51,31,213,31,85,31,236,31,240,31,240,30,240,29,241,31,150,31,254,31,164,31,1,31,105,31,66,31,32,31,131,31,109,31,188,31,44,31,75,31,169,31,199,31,199,30,149,31,130,31,150,31,150,30,213,31,166,31,69,31,69,30,184,31,33,31,187,31,187,30,122,31,12,31,106,31,242,31,102,31,102,30,243,31,30,31,136,31,105,31,23,31,23,30,181,31,181,30,231,31,150,31,150,30,13,31,28,31,102,31,199,31,59,31,205,31,37,31,196,31,187,31,163,31,69,31,206,31,134,31,244,31,3,31,3,30,3,29,202,31,171,31,63,31,168,31,185,31,159,31,2,31,22,31,234,31,35,31,35,30,46,31,173,31,62,31,167,31,189,31,177,31,177,30,63,31,179,31,8,31,233,31,72,31,104,31,45,31,45,30,74,31,74,30,224,31,73,31,37,31,63,31,62,31,97,31,213,31,213,30,213,29,253,31,239,31,239,31,155,31,143,31,248,31,204,31,204,30,204,29,50,31,167,31,167,30,167,29,167,28,199,31,251,31,50,31,126,31,55,31,199,31,169,31,105,31,105,30,236,31,236,30,227,31,178,31,204,31,204,30,48,31,122,31,158,31,205,31,60,31,149,31,26,31,119,31,120,31,120,30,52,31,157,31,159,31,167,31,62,31,62,30,249,31,164,31,158,31,68,31,123,31,219,31,180,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
