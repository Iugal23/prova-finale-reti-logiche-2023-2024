-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 178;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (59,0,0,0,63,0,0,0,85,0,0,0,98,0,122,0,201,0,45,0,226,0,229,0,131,0,43,0,59,0,0,0,101,0,89,0,145,0,132,0,42,0,167,0,174,0,120,0,210,0,12,0,63,0,189,0,166,0,189,0,222,0,27,0,8,0,88,0,18,0,174,0,97,0,13,0,0,0,29,0,157,0,189,0,153,0,114,0,35,0,0,0,5,0,115,0,0,0,0,0,202,0,176,0,0,0,236,0,65,0,65,0,76,0,0,0,116,0,25,0,51,0,108,0,0,0,164,0,135,0,0,0,0,0,215,0,214,0,85,0,88,0,15,0,217,0,159,0,49,0,32,0,129,0,168,0,25,0,0,0,213,0,119,0,122,0,0,0,37,0,202,0,103,0,141,0,113,0,81,0,0,0,231,0,0,0,191,0,225,0,2,0,129,0,0,0,195,0,103,0,114,0,60,0,0,0,84,0,29,0,243,0,71,0,53,0,162,0,213,0,226,0,0,0,0,0,129,0,122,0,0,0,250,0,34,0,0,0,33,0,0,0,132,0,0,0,235,0,160,0,132,0,3,0,230,0,18,0,48,0,136,0,0,0,241,0,130,0,23,0,175,0,209,0,152,0,160,0,62,0,0,0,78,0,41,0,0,0,243,0,167,0,146,0,0,0,0,0,0,0,40,0,80,0,111,0,188,0,220,0,95,0,144,0,24,0,115,0,30,0,0,0,29,0,175,0,0,0,131,0,0,0,24,0,0,0,218,0,131,0,15,0,20,0,25,0,67,0,186,0,186,0,75,0,11,0);
signal scenario_full  : scenario_type := (59,31,59,30,63,31,63,30,85,31,85,30,98,31,122,31,201,31,45,31,226,31,229,31,131,31,43,31,59,31,59,30,101,31,89,31,145,31,132,31,42,31,167,31,174,31,120,31,210,31,12,31,63,31,189,31,166,31,189,31,222,31,27,31,8,31,88,31,18,31,174,31,97,31,13,31,13,30,29,31,157,31,189,31,153,31,114,31,35,31,35,30,5,31,115,31,115,30,115,29,202,31,176,31,176,30,236,31,65,31,65,31,76,31,76,30,116,31,25,31,51,31,108,31,108,30,164,31,135,31,135,30,135,29,215,31,214,31,85,31,88,31,15,31,217,31,159,31,49,31,32,31,129,31,168,31,25,31,25,30,213,31,119,31,122,31,122,30,37,31,202,31,103,31,141,31,113,31,81,31,81,30,231,31,231,30,191,31,225,31,2,31,129,31,129,30,195,31,103,31,114,31,60,31,60,30,84,31,29,31,243,31,71,31,53,31,162,31,213,31,226,31,226,30,226,29,129,31,122,31,122,30,250,31,34,31,34,30,33,31,33,30,132,31,132,30,235,31,160,31,132,31,3,31,230,31,18,31,48,31,136,31,136,30,241,31,130,31,23,31,175,31,209,31,152,31,160,31,62,31,62,30,78,31,41,31,41,30,243,31,167,31,146,31,146,30,146,29,146,28,40,31,80,31,111,31,188,31,220,31,95,31,144,31,24,31,115,31,30,31,30,30,29,31,175,31,175,30,131,31,131,30,24,31,24,30,218,31,131,31,15,31,20,31,25,31,67,31,186,31,186,31,75,31,11,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
