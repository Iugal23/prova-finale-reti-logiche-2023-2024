-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_587 is
end project_tb_587;

architecture project_tb_arch_587 of project_tb_587 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 898;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,207,0,241,0,180,0,66,0,0,0,0,0,137,0,116,0,216,0,0,0,0,0,67,0,176,0,230,0,50,0,129,0,0,0,112,0,224,0,210,0,0,0,33,0,0,0,211,0,0,0,242,0,21,0,0,0,146,0,118,0,241,0,205,0,114,0,48,0,40,0,159,0,1,0,181,0,216,0,0,0,91,0,169,0,65,0,0,0,131,0,12,0,219,0,0,0,7,0,0,0,21,0,0,0,0,0,0,0,193,0,46,0,155,0,64,0,223,0,199,0,0,0,72,0,51,0,0,0,181,0,129,0,31,0,96,0,8,0,0,0,102,0,38,0,150,0,14,0,45,0,0,0,0,0,177,0,0,0,188,0,203,0,76,0,28,0,0,0,0,0,104,0,235,0,240,0,0,0,126,0,172,0,193,0,0,0,0,0,48,0,0,0,0,0,221,0,126,0,122,0,0,0,226,0,91,0,218,0,0,0,202,0,0,0,165,0,6,0,98,0,0,0,169,0,5,0,98,0,217,0,123,0,148,0,0,0,0,0,0,0,244,0,133,0,7,0,24,0,121,0,95,0,57,0,125,0,29,0,16,0,57,0,253,0,207,0,187,0,0,0,176,0,18,0,78,0,0,0,0,0,0,0,103,0,0,0,152,0,0,0,141,0,47,0,126,0,35,0,12,0,0,0,132,0,250,0,195,0,138,0,0,0,29,0,201,0,182,0,126,0,0,0,48,0,162,0,57,0,207,0,32,0,0,0,105,0,197,0,198,0,138,0,144,0,161,0,173,0,28,0,206,0,164,0,95,0,28,0,161,0,165,0,0,0,223,0,8,0,0,0,0,0,90,0,228,0,210,0,0,0,125,0,6,0,35,0,56,0,190,0,226,0,255,0,169,0,173,0,51,0,69,0,57,0,0,0,132,0,39,0,65,0,0,0,72,0,0,0,189,0,3,0,0,0,134,0,214,0,0,0,147,0,76,0,142,0,54,0,33,0,167,0,54,0,168,0,58,0,168,0,145,0,199,0,13,0,67,0,180,0,0,0,48,0,0,0,143,0,0,0,114,0,18,0,89,0,242,0,65,0,152,0,247,0,0,0,89,0,149,0,78,0,110,0,8,0,207,0,100,0,254,0,162,0,221,0,78,0,63,0,0,0,135,0,184,0,30,0,183,0,25,0,154,0,0,0,128,0,121,0,0,0,100,0,252,0,0,0,220,0,214,0,0,0,0,0,242,0,0,0,0,0,93,0,235,0,213,0,65,0,0,0,78,0,35,0,0,0,59,0,0,0,197,0,4,0,31,0,9,0,0,0,31,0,0,0,193,0,0,0,0,0,0,0,0,0,157,0,72,0,151,0,80,0,46,0,166,0,201,0,11,0,0,0,57,0,199,0,81,0,0,0,176,0,221,0,0,0,111,0,46,0,188,0,0,0,149,0,0,0,163,0,0,0,33,0,15,0,189,0,1,0,66,0,77,0,229,0,110,0,179,0,0,0,0,0,211,0,183,0,242,0,190,0,124,0,9,0,36,0,250,0,91,0,20,0,54,0,2,0,124,0,107,0,194,0,45,0,36,0,166,0,0,0,83,0,119,0,203,0,194,0,65,0,142,0,0,0,0,0,0,0,104,0,0,0,133,0,0,0,48,0,219,0,250,0,78,0,130,0,126,0,0,0,80,0,168,0,178,0,127,0,225,0,242,0,37,0,0,0,18,0,71,0,31,0,114,0,0,0,18,0,16,0,158,0,49,0,155,0,113,0,78,0,12,0,192,0,171,0,0,0,202,0,219,0,0,0,242,0,228,0,115,0,0,0,240,0,62,0,5,0,105,0,61,0,173,0,93,0,203,0,71,0,6,0,139,0,62,0,94,0,147,0,234,0,216,0,0,0,0,0,127,0,167,0,0,0,0,0,153,0,0,0,245,0,83,0,76,0,0,0,239,0,226,0,185,0,113,0,123,0,0,0,0,0,0,0,0,0,0,0,184,0,92,0,87,0,77,0,80,0,137,0,252,0,85,0,141,0,0,0,38,0,124,0,0,0,70,0,228,0,93,0,26,0,72,0,155,0,92,0,198,0,103,0,0,0,114,0,0,0,176,0,241,0,167,0,76,0,28,0,80,0,105,0,212,0,0,0,0,0,139,0,174,0,203,0,0,0,0,0,31,0,116,0,248,0,121,0,203,0,84,0,118,0,139,0,191,0,3,0,94,0,99,0,102,0,0,0,196,0,5,0,238,0,8,0,169,0,41,0,50,0,245,0,127,0,102,0,166,0,53,0,21,0,23,0,103,0,166,0,44,0,6,0,222,0,192,0,84,0,238,0,178,0,121,0,22,0,55,0,61,0,71,0,104,0,149,0,25,0,226,0,87,0,86,0,206,0,217,0,22,0,0,0,90,0,18,0,34,0,0,0,37,0,165,0,0,0,34,0,151,0,0,0,47,0,116,0,0,0,82,0,123,0,252,0,23,0,22,0,167,0,0,0,200,0,212,0,0,0,60,0,0,0,0,0,158,0,119,0,72,0,0,0,0,0,45,0,173,0,212,0,238,0,170,0,73,0,146,0,80,0,79,0,233,0,95,0,0,0,0,0,83,0,187,0,173,0,156,0,0,0,0,0,150,0,149,0,0,0,112,0,62,0,76,0,0,0,192,0,167,0,201,0,204,0,8,0,0,0,0,0,210,0,0,0,0,0,0,0,123,0,200,0,231,0,249,0,235,0,0,0,181,0,2,0,0,0,134,0,218,0,98,0,171,0,220,0,187,0,133,0,55,0,88,0,0,0,26,0,83,0,0,0,151,0,82,0,60,0,29,0,138,0,8,0,171,0,164,0,191,0,135,0,44,0,121,0,0,0,0,0,228,0,137,0,230,0,199,0,67,0,48,0,138,0,31,0,0,0,0,0,139,0,37,0,222,0,0,0,224,0,254,0,0,0,229,0,29,0,126,0,117,0,153,0,135,0,167,0,0,0,142,0,172,0,221,0,28,0,193,0,0,0,0,0,6,0,0,0,0,0,66,0,178,0,126,0,0,0,0,0,114,0,0,0,151,0,18,0,196,0,149,0,79,0,90,0,0,0,0,0,0,0,222,0,185,0,0,0,156,0,10,0,128,0,60,0,203,0,115,0,254,0,88,0,0,0,72,0,44,0,216,0,189,0,53,0,0,0,10,0,124,0,0,0,0,0,135,0,68,0,67,0,113,0,0,0,0,0,137,0,165,0,25,0,253,0,146,0,55,0,0,0,53,0,205,0,0,0,102,0,63,0,160,0,249,0,21,0,251,0,253,0,162,0,0,0,0,0,6,0,0,0,110,0,222,0,65,0,224,0,53,0,182,0,0,0,85,0,0,0,88,0,172,0,0,0,248,0,200,0,3,0,8,0,163,0,0,0,117,0,124,0,173,0,136,0,59,0,41,0,229,0,68,0,203,0,138,0,187,0,210,0,0,0,133,0,236,0,0,0,149,0,230,0,65,0,0,0,246,0,11,0,103,0,62,0,15,0,217,0,67,0,22,0,230,0,211,0,0,0,44,0,41,0,123,0,138,0,220,0,0,0,29,0,99,0,0,0,251,0,0,0,43,0,0,0,229,0,66,0,231,0,133,0,197,0,38,0,148,0,123,0,11,0,128,0,60,0,0,0,23,0,62,0,0,0,146,0,0,0,201,0,244,0,186,0,0,0,131,0,0,0,102,0,142,0,45,0,15,0,6,0,0,0,0,0,132,0,0,0,0,0,73,0,75,0,0,0,0,0,37,0,234,0,203,0,135,0,66,0,121,0,154,0,149,0,106,0,203,0,0,0,23,0,67,0,68,0,205,0,138,0,217,0,190,0,120,0,0,0,193,0,0,0,0,0,114,0,161,0,0,0,217,0,248,0,76,0,130,0,149,0,42,0,172,0,0,0,30,0,168,0,6,0,15,0,0,0,54,0,195,0,0,0,171,0,90,0,245,0,185,0,0,0,210,0,152,0,76,0,52,0,24,0,230,0,0,0,46,0,164,0,0,0,25,0,0,0,0,0);
signal scenario_full  : scenario_type := (0,0,207,31,241,31,180,31,66,31,66,30,66,29,137,31,116,31,216,31,216,30,216,29,67,31,176,31,230,31,50,31,129,31,129,30,112,31,224,31,210,31,210,30,33,31,33,30,211,31,211,30,242,31,21,31,21,30,146,31,118,31,241,31,205,31,114,31,48,31,40,31,159,31,1,31,181,31,216,31,216,30,91,31,169,31,65,31,65,30,131,31,12,31,219,31,219,30,7,31,7,30,21,31,21,30,21,29,21,28,193,31,46,31,155,31,64,31,223,31,199,31,199,30,72,31,51,31,51,30,181,31,129,31,31,31,96,31,8,31,8,30,102,31,38,31,150,31,14,31,45,31,45,30,45,29,177,31,177,30,188,31,203,31,76,31,28,31,28,30,28,29,104,31,235,31,240,31,240,30,126,31,172,31,193,31,193,30,193,29,48,31,48,30,48,29,221,31,126,31,122,31,122,30,226,31,91,31,218,31,218,30,202,31,202,30,165,31,6,31,98,31,98,30,169,31,5,31,98,31,217,31,123,31,148,31,148,30,148,29,148,28,244,31,133,31,7,31,24,31,121,31,95,31,57,31,125,31,29,31,16,31,57,31,253,31,207,31,187,31,187,30,176,31,18,31,78,31,78,30,78,29,78,28,103,31,103,30,152,31,152,30,141,31,47,31,126,31,35,31,12,31,12,30,132,31,250,31,195,31,138,31,138,30,29,31,201,31,182,31,126,31,126,30,48,31,162,31,57,31,207,31,32,31,32,30,105,31,197,31,198,31,138,31,144,31,161,31,173,31,28,31,206,31,164,31,95,31,28,31,161,31,165,31,165,30,223,31,8,31,8,30,8,29,90,31,228,31,210,31,210,30,125,31,6,31,35,31,56,31,190,31,226,31,255,31,169,31,173,31,51,31,69,31,57,31,57,30,132,31,39,31,65,31,65,30,72,31,72,30,189,31,3,31,3,30,134,31,214,31,214,30,147,31,76,31,142,31,54,31,33,31,167,31,54,31,168,31,58,31,168,31,145,31,199,31,13,31,67,31,180,31,180,30,48,31,48,30,143,31,143,30,114,31,18,31,89,31,242,31,65,31,152,31,247,31,247,30,89,31,149,31,78,31,110,31,8,31,207,31,100,31,254,31,162,31,221,31,78,31,63,31,63,30,135,31,184,31,30,31,183,31,25,31,154,31,154,30,128,31,121,31,121,30,100,31,252,31,252,30,220,31,214,31,214,30,214,29,242,31,242,30,242,29,93,31,235,31,213,31,65,31,65,30,78,31,35,31,35,30,59,31,59,30,197,31,4,31,31,31,9,31,9,30,31,31,31,30,193,31,193,30,193,29,193,28,193,27,157,31,72,31,151,31,80,31,46,31,166,31,201,31,11,31,11,30,57,31,199,31,81,31,81,30,176,31,221,31,221,30,111,31,46,31,188,31,188,30,149,31,149,30,163,31,163,30,33,31,15,31,189,31,1,31,66,31,77,31,229,31,110,31,179,31,179,30,179,29,211,31,183,31,242,31,190,31,124,31,9,31,36,31,250,31,91,31,20,31,54,31,2,31,124,31,107,31,194,31,45,31,36,31,166,31,166,30,83,31,119,31,203,31,194,31,65,31,142,31,142,30,142,29,142,28,104,31,104,30,133,31,133,30,48,31,219,31,250,31,78,31,130,31,126,31,126,30,80,31,168,31,178,31,127,31,225,31,242,31,37,31,37,30,18,31,71,31,31,31,114,31,114,30,18,31,16,31,158,31,49,31,155,31,113,31,78,31,12,31,192,31,171,31,171,30,202,31,219,31,219,30,242,31,228,31,115,31,115,30,240,31,62,31,5,31,105,31,61,31,173,31,93,31,203,31,71,31,6,31,139,31,62,31,94,31,147,31,234,31,216,31,216,30,216,29,127,31,167,31,167,30,167,29,153,31,153,30,245,31,83,31,76,31,76,30,239,31,226,31,185,31,113,31,123,31,123,30,123,29,123,28,123,27,123,26,184,31,92,31,87,31,77,31,80,31,137,31,252,31,85,31,141,31,141,30,38,31,124,31,124,30,70,31,228,31,93,31,26,31,72,31,155,31,92,31,198,31,103,31,103,30,114,31,114,30,176,31,241,31,167,31,76,31,28,31,80,31,105,31,212,31,212,30,212,29,139,31,174,31,203,31,203,30,203,29,31,31,116,31,248,31,121,31,203,31,84,31,118,31,139,31,191,31,3,31,94,31,99,31,102,31,102,30,196,31,5,31,238,31,8,31,169,31,41,31,50,31,245,31,127,31,102,31,166,31,53,31,21,31,23,31,103,31,166,31,44,31,6,31,222,31,192,31,84,31,238,31,178,31,121,31,22,31,55,31,61,31,71,31,104,31,149,31,25,31,226,31,87,31,86,31,206,31,217,31,22,31,22,30,90,31,18,31,34,31,34,30,37,31,165,31,165,30,34,31,151,31,151,30,47,31,116,31,116,30,82,31,123,31,252,31,23,31,22,31,167,31,167,30,200,31,212,31,212,30,60,31,60,30,60,29,158,31,119,31,72,31,72,30,72,29,45,31,173,31,212,31,238,31,170,31,73,31,146,31,80,31,79,31,233,31,95,31,95,30,95,29,83,31,187,31,173,31,156,31,156,30,156,29,150,31,149,31,149,30,112,31,62,31,76,31,76,30,192,31,167,31,201,31,204,31,8,31,8,30,8,29,210,31,210,30,210,29,210,28,123,31,200,31,231,31,249,31,235,31,235,30,181,31,2,31,2,30,134,31,218,31,98,31,171,31,220,31,187,31,133,31,55,31,88,31,88,30,26,31,83,31,83,30,151,31,82,31,60,31,29,31,138,31,8,31,171,31,164,31,191,31,135,31,44,31,121,31,121,30,121,29,228,31,137,31,230,31,199,31,67,31,48,31,138,31,31,31,31,30,31,29,139,31,37,31,222,31,222,30,224,31,254,31,254,30,229,31,29,31,126,31,117,31,153,31,135,31,167,31,167,30,142,31,172,31,221,31,28,31,193,31,193,30,193,29,6,31,6,30,6,29,66,31,178,31,126,31,126,30,126,29,114,31,114,30,151,31,18,31,196,31,149,31,79,31,90,31,90,30,90,29,90,28,222,31,185,31,185,30,156,31,10,31,128,31,60,31,203,31,115,31,254,31,88,31,88,30,72,31,44,31,216,31,189,31,53,31,53,30,10,31,124,31,124,30,124,29,135,31,68,31,67,31,113,31,113,30,113,29,137,31,165,31,25,31,253,31,146,31,55,31,55,30,53,31,205,31,205,30,102,31,63,31,160,31,249,31,21,31,251,31,253,31,162,31,162,30,162,29,6,31,6,30,110,31,222,31,65,31,224,31,53,31,182,31,182,30,85,31,85,30,88,31,172,31,172,30,248,31,200,31,3,31,8,31,163,31,163,30,117,31,124,31,173,31,136,31,59,31,41,31,229,31,68,31,203,31,138,31,187,31,210,31,210,30,133,31,236,31,236,30,149,31,230,31,65,31,65,30,246,31,11,31,103,31,62,31,15,31,217,31,67,31,22,31,230,31,211,31,211,30,44,31,41,31,123,31,138,31,220,31,220,30,29,31,99,31,99,30,251,31,251,30,43,31,43,30,229,31,66,31,231,31,133,31,197,31,38,31,148,31,123,31,11,31,128,31,60,31,60,30,23,31,62,31,62,30,146,31,146,30,201,31,244,31,186,31,186,30,131,31,131,30,102,31,142,31,45,31,15,31,6,31,6,30,6,29,132,31,132,30,132,29,73,31,75,31,75,30,75,29,37,31,234,31,203,31,135,31,66,31,121,31,154,31,149,31,106,31,203,31,203,30,23,31,67,31,68,31,205,31,138,31,217,31,190,31,120,31,120,30,193,31,193,30,193,29,114,31,161,31,161,30,217,31,248,31,76,31,130,31,149,31,42,31,172,31,172,30,30,31,168,31,6,31,15,31,15,30,54,31,195,31,195,30,171,31,90,31,245,31,185,31,185,30,210,31,152,31,76,31,52,31,24,31,230,31,230,30,46,31,164,31,164,30,25,31,25,30,25,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
