-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_628 is
end project_tb_628;

architecture project_tb_arch_628 of project_tb_628 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 821;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (128,0,251,0,75,0,50,0,152,0,7,0,0,0,0,0,228,0,0,0,231,0,0,0,147,0,185,0,73,0,153,0,213,0,224,0,43,0,155,0,0,0,38,0,146,0,0,0,18,0,0,0,0,0,0,0,50,0,0,0,232,0,0,0,190,0,216,0,0,0,67,0,112,0,208,0,0,0,0,0,204,0,175,0,229,0,136,0,0,0,0,0,174,0,5,0,148,0,248,0,240,0,0,0,0,0,0,0,139,0,36,0,20,0,5,0,0,0,150,0,70,0,0,0,114,0,108,0,141,0,103,0,20,0,245,0,234,0,62,0,58,0,0,0,109,0,193,0,208,0,169,0,0,0,17,0,65,0,17,0,198,0,62,0,192,0,203,0,75,0,0,0,114,0,229,0,178,0,4,0,10,0,152,0,0,0,50,0,27,0,85,0,119,0,0,0,60,0,11,0,0,0,0,0,139,0,0,0,69,0,0,0,104,0,36,0,158,0,30,0,235,0,138,0,0,0,0,0,40,0,115,0,61,0,236,0,0,0,187,0,83,0,134,0,103,0,198,0,186,0,227,0,0,0,0,0,183,0,0,0,68,0,0,0,91,0,202,0,104,0,0,0,0,0,11,0,0,0,147,0,0,0,38,0,0,0,192,0,84,0,221,0,157,0,150,0,0,0,164,0,179,0,233,0,249,0,95,0,1,0,104,0,30,0,0,0,46,0,41,0,0,0,177,0,146,0,143,0,20,0,2,0,0,0,58,0,153,0,109,0,236,0,238,0,32,0,68,0,69,0,43,0,30,0,253,0,63,0,178,0,0,0,0,0,60,0,0,0,230,0,0,0,0,0,126,0,174,0,70,0,231,0,228,0,37,0,0,0,173,0,128,0,81,0,136,0,233,0,111,0,0,0,155,0,0,0,189,0,0,0,155,0,184,0,133,0,124,0,111,0,241,0,0,0,145,0,164,0,183,0,18,0,119,0,1,0,98,0,160,0,41,0,129,0,235,0,19,0,94,0,227,0,43,0,249,0,13,0,59,0,0,0,247,0,58,0,61,0,243,0,130,0,111,0,23,0,245,0,21,0,87,0,141,0,0,0,17,0,229,0,30,0,124,0,115,0,84,0,96,0,203,0,0,0,0,0,241,0,192,0,0,0,167,0,0,0,187,0,112,0,230,0,64,0,203,0,5,0,145,0,123,0,17,0,0,0,143,0,225,0,66,0,201,0,215,0,164,0,132,0,212,0,121,0,156,0,107,0,0,0,97,0,111,0,141,0,50,0,238,0,0,0,165,0,102,0,98,0,87,0,87,0,209,0,230,0,96,0,69,0,0,0,147,0,255,0,240,0,85,0,91,0,212,0,191,0,0,0,50,0,201,0,22,0,193,0,151,0,123,0,71,0,55,0,112,0,69,0,181,0,197,0,25,0,210,0,141,0,186,0,119,0,148,0,0,0,0,0,218,0,161,0,235,0,40,0,114,0,0,0,3,0,244,0,20,0,0,0,238,0,84,0,251,0,41,0,195,0,0,0,0,0,0,0,180,0,0,0,227,0,145,0,86,0,43,0,53,0,90,0,0,0,0,0,135,0,227,0,52,0,0,0,214,0,149,0,90,0,106,0,39,0,170,0,164,0,0,0,0,0,67,0,198,0,0,0,2,0,244,0,202,0,252,0,0,0,28,0,126,0,0,0,160,0,0,0,203,0,143,0,67,0,116,0,136,0,135,0,0,0,234,0,142,0,80,0,28,0,94,0,115,0,114,0,161,0,37,0,252,0,190,0,188,0,69,0,9,0,61,0,216,0,235,0,87,0,189,0,0,0,131,0,36,0,205,0,45,0,44,0,93,0,248,0,24,0,118,0,1,0,58,0,0,0,0,0,231,0,94,0,244,0,240,0,0,0,244,0,246,0,150,0,35,0,253,0,200,0,58,0,250,0,0,0,101,0,7,0,177,0,159,0,242,0,0,0,7,0,157,0,198,0,72,0,74,0,0,0,0,0,177,0,24,0,0,0,253,0,0,0,150,0,172,0,0,0,0,0,161,0,160,0,245,0,227,0,236,0,0,0,188,0,35,0,0,0,227,0,149,0,67,0,26,0,154,0,0,0,107,0,149,0,20,0,204,0,0,0,111,0,0,0,237,0,0,0,191,0,190,0,0,0,218,0,181,0,143,0,58,0,63,0,0,0,0,0,224,0,0,0,246,0,136,0,3,0,0,0,0,0,215,0,224,0,144,0,49,0,66,0,0,0,28,0,242,0,79,0,241,0,251,0,139,0,0,0,0,0,118,0,191,0,208,0,0,0,118,0,0,0,104,0,216,0,221,0,70,0,215,0,0,0,109,0,167,0,24,0,157,0,105,0,48,0,119,0,12,0,169,0,22,0,97,0,122,0,164,0,0,0,46,0,194,0,116,0,0,0,0,0,0,0,5,0,18,0,219,0,238,0,235,0,147,0,23,0,184,0,28,0,54,0,33,0,151,0,33,0,220,0,226,0,132,0,52,0,69,0,226,0,35,0,7,0,224,0,236,0,12,0,0,0,128,0,0,0,197,0,121,0,240,0,240,0,248,0,52,0,240,0,219,0,78,0,214,0,121,0,242,0,0,0,160,0,220,0,24,0,192,0,130,0,3,0,45,0,70,0,109,0,150,0,26,0,0,0,0,0,163,0,0,0,186,0,0,0,0,0,131,0,89,0,209,0,119,0,168,0,0,0,50,0,162,0,189,0,185,0,0,0,221,0,0,0,238,0,2,0,48,0,0,0,86,0,0,0,62,0,221,0,121,0,153,0,20,0,207,0,0,0,37,0,0,0,0,0,0,0,80,0,144,0,8,0,135,0,216,0,127,0,0,0,75,0,17,0,251,0,245,0,150,0,229,0,75,0,228,0,0,0,137,0,22,0,48,0,95,0,205,0,246,0,177,0,123,0,241,0,151,0,96,0,235,0,112,0,141,0,0,0,0,0,84,0,115,0,49,0,136,0,15,0,184,0,249,0,182,0,242,0,250,0,114,0,0,0,1,0,0,0,181,0,120,0,212,0,0,0,195,0,172,0,237,0,100,0,109,0,233,0,109,0,183,0,0,0,0,0,233,0,0,0,96,0,0,0,120,0,82,0,6,0,0,0,0,0,192,0,237,0,236,0,160,0,114,0,32,0,61,0,53,0,159,0,165,0,121,0,156,0,0,0,232,0,102,0,36,0,140,0,0,0,250,0,36,0,116,0,230,0,162,0,0,0,102,0,0,0,133,0,0,0,208,0,90,0,9,0,210,0,114,0,51,0,70,0,217,0,144,0,0,0,132,0,4,0,0,0,75,0,58,0,59,0,194,0,214,0,106,0,131,0,207,0,191,0,27,0,80,0,184,0,93,0,0,0,17,0,90,0,217,0,232,0,83,0,59,0,159,0,207,0,66,0,156,0,29,0,11,0,62,0,74,0,93,0,250,0,249,0,0,0,97,0,45,0,232,0,106,0,218,0,186,0,0,0,40,0,164,0,51,0,21,0,242,0,253,0,0,0,3,0,128,0,80,0,108,0,133,0,102,0,78,0,44,0,229,0,25,0,129,0,187,0,113,0,77,0,7,0,184,0,125,0,18,0,0,0,149,0,123,0,80,0,0,0,252,0,148,0,0,0,6,0,170,0,164,0,24,0,80,0,139,0,179,0,149,0,67,0,44,0);
signal scenario_full  : scenario_type := (128,31,251,31,75,31,50,31,152,31,7,31,7,30,7,29,228,31,228,30,231,31,231,30,147,31,185,31,73,31,153,31,213,31,224,31,43,31,155,31,155,30,38,31,146,31,146,30,18,31,18,30,18,29,18,28,50,31,50,30,232,31,232,30,190,31,216,31,216,30,67,31,112,31,208,31,208,30,208,29,204,31,175,31,229,31,136,31,136,30,136,29,174,31,5,31,148,31,248,31,240,31,240,30,240,29,240,28,139,31,36,31,20,31,5,31,5,30,150,31,70,31,70,30,114,31,108,31,141,31,103,31,20,31,245,31,234,31,62,31,58,31,58,30,109,31,193,31,208,31,169,31,169,30,17,31,65,31,17,31,198,31,62,31,192,31,203,31,75,31,75,30,114,31,229,31,178,31,4,31,10,31,152,31,152,30,50,31,27,31,85,31,119,31,119,30,60,31,11,31,11,30,11,29,139,31,139,30,69,31,69,30,104,31,36,31,158,31,30,31,235,31,138,31,138,30,138,29,40,31,115,31,61,31,236,31,236,30,187,31,83,31,134,31,103,31,198,31,186,31,227,31,227,30,227,29,183,31,183,30,68,31,68,30,91,31,202,31,104,31,104,30,104,29,11,31,11,30,147,31,147,30,38,31,38,30,192,31,84,31,221,31,157,31,150,31,150,30,164,31,179,31,233,31,249,31,95,31,1,31,104,31,30,31,30,30,46,31,41,31,41,30,177,31,146,31,143,31,20,31,2,31,2,30,58,31,153,31,109,31,236,31,238,31,32,31,68,31,69,31,43,31,30,31,253,31,63,31,178,31,178,30,178,29,60,31,60,30,230,31,230,30,230,29,126,31,174,31,70,31,231,31,228,31,37,31,37,30,173,31,128,31,81,31,136,31,233,31,111,31,111,30,155,31,155,30,189,31,189,30,155,31,184,31,133,31,124,31,111,31,241,31,241,30,145,31,164,31,183,31,18,31,119,31,1,31,98,31,160,31,41,31,129,31,235,31,19,31,94,31,227,31,43,31,249,31,13,31,59,31,59,30,247,31,58,31,61,31,243,31,130,31,111,31,23,31,245,31,21,31,87,31,141,31,141,30,17,31,229,31,30,31,124,31,115,31,84,31,96,31,203,31,203,30,203,29,241,31,192,31,192,30,167,31,167,30,187,31,112,31,230,31,64,31,203,31,5,31,145,31,123,31,17,31,17,30,143,31,225,31,66,31,201,31,215,31,164,31,132,31,212,31,121,31,156,31,107,31,107,30,97,31,111,31,141,31,50,31,238,31,238,30,165,31,102,31,98,31,87,31,87,31,209,31,230,31,96,31,69,31,69,30,147,31,255,31,240,31,85,31,91,31,212,31,191,31,191,30,50,31,201,31,22,31,193,31,151,31,123,31,71,31,55,31,112,31,69,31,181,31,197,31,25,31,210,31,141,31,186,31,119,31,148,31,148,30,148,29,218,31,161,31,235,31,40,31,114,31,114,30,3,31,244,31,20,31,20,30,238,31,84,31,251,31,41,31,195,31,195,30,195,29,195,28,180,31,180,30,227,31,145,31,86,31,43,31,53,31,90,31,90,30,90,29,135,31,227,31,52,31,52,30,214,31,149,31,90,31,106,31,39,31,170,31,164,31,164,30,164,29,67,31,198,31,198,30,2,31,244,31,202,31,252,31,252,30,28,31,126,31,126,30,160,31,160,30,203,31,143,31,67,31,116,31,136,31,135,31,135,30,234,31,142,31,80,31,28,31,94,31,115,31,114,31,161,31,37,31,252,31,190,31,188,31,69,31,9,31,61,31,216,31,235,31,87,31,189,31,189,30,131,31,36,31,205,31,45,31,44,31,93,31,248,31,24,31,118,31,1,31,58,31,58,30,58,29,231,31,94,31,244,31,240,31,240,30,244,31,246,31,150,31,35,31,253,31,200,31,58,31,250,31,250,30,101,31,7,31,177,31,159,31,242,31,242,30,7,31,157,31,198,31,72,31,74,31,74,30,74,29,177,31,24,31,24,30,253,31,253,30,150,31,172,31,172,30,172,29,161,31,160,31,245,31,227,31,236,31,236,30,188,31,35,31,35,30,227,31,149,31,67,31,26,31,154,31,154,30,107,31,149,31,20,31,204,31,204,30,111,31,111,30,237,31,237,30,191,31,190,31,190,30,218,31,181,31,143,31,58,31,63,31,63,30,63,29,224,31,224,30,246,31,136,31,3,31,3,30,3,29,215,31,224,31,144,31,49,31,66,31,66,30,28,31,242,31,79,31,241,31,251,31,139,31,139,30,139,29,118,31,191,31,208,31,208,30,118,31,118,30,104,31,216,31,221,31,70,31,215,31,215,30,109,31,167,31,24,31,157,31,105,31,48,31,119,31,12,31,169,31,22,31,97,31,122,31,164,31,164,30,46,31,194,31,116,31,116,30,116,29,116,28,5,31,18,31,219,31,238,31,235,31,147,31,23,31,184,31,28,31,54,31,33,31,151,31,33,31,220,31,226,31,132,31,52,31,69,31,226,31,35,31,7,31,224,31,236,31,12,31,12,30,128,31,128,30,197,31,121,31,240,31,240,31,248,31,52,31,240,31,219,31,78,31,214,31,121,31,242,31,242,30,160,31,220,31,24,31,192,31,130,31,3,31,45,31,70,31,109,31,150,31,26,31,26,30,26,29,163,31,163,30,186,31,186,30,186,29,131,31,89,31,209,31,119,31,168,31,168,30,50,31,162,31,189,31,185,31,185,30,221,31,221,30,238,31,2,31,48,31,48,30,86,31,86,30,62,31,221,31,121,31,153,31,20,31,207,31,207,30,37,31,37,30,37,29,37,28,80,31,144,31,8,31,135,31,216,31,127,31,127,30,75,31,17,31,251,31,245,31,150,31,229,31,75,31,228,31,228,30,137,31,22,31,48,31,95,31,205,31,246,31,177,31,123,31,241,31,151,31,96,31,235,31,112,31,141,31,141,30,141,29,84,31,115,31,49,31,136,31,15,31,184,31,249,31,182,31,242,31,250,31,114,31,114,30,1,31,1,30,181,31,120,31,212,31,212,30,195,31,172,31,237,31,100,31,109,31,233,31,109,31,183,31,183,30,183,29,233,31,233,30,96,31,96,30,120,31,82,31,6,31,6,30,6,29,192,31,237,31,236,31,160,31,114,31,32,31,61,31,53,31,159,31,165,31,121,31,156,31,156,30,232,31,102,31,36,31,140,31,140,30,250,31,36,31,116,31,230,31,162,31,162,30,102,31,102,30,133,31,133,30,208,31,90,31,9,31,210,31,114,31,51,31,70,31,217,31,144,31,144,30,132,31,4,31,4,30,75,31,58,31,59,31,194,31,214,31,106,31,131,31,207,31,191,31,27,31,80,31,184,31,93,31,93,30,17,31,90,31,217,31,232,31,83,31,59,31,159,31,207,31,66,31,156,31,29,31,11,31,62,31,74,31,93,31,250,31,249,31,249,30,97,31,45,31,232,31,106,31,218,31,186,31,186,30,40,31,164,31,51,31,21,31,242,31,253,31,253,30,3,31,128,31,80,31,108,31,133,31,102,31,78,31,44,31,229,31,25,31,129,31,187,31,113,31,77,31,7,31,184,31,125,31,18,31,18,30,149,31,123,31,80,31,80,30,252,31,148,31,148,30,6,31,170,31,164,31,24,31,80,31,139,31,179,31,149,31,67,31,44,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
