-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_100 is
end project_tb_100;

architecture project_tb_arch_100 of project_tb_100 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 776;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (116,0,11,0,215,0,126,0,63,0,100,0,227,0,83,0,242,0,184,0,231,0,190,0,106,0,15,0,190,0,179,0,22,0,50,0,240,0,205,0,126,0,94,0,49,0,10,0,238,0,187,0,0,0,81,0,6,0,3,0,60,0,0,0,237,0,0,0,24,0,122,0,0,0,98,0,84,0,0,0,204,0,0,0,0,0,0,0,216,0,0,0,168,0,128,0,0,0,55,0,107,0,234,0,0,0,0,0,202,0,0,0,0,0,202,0,177,0,86,0,0,0,137,0,125,0,220,0,49,0,0,0,119,0,94,0,219,0,161,0,103,0,56,0,167,0,0,0,0,0,0,0,157,0,223,0,172,0,194,0,8,0,95,0,0,0,0,0,0,0,0,0,210,0,0,0,0,0,86,0,0,0,0,0,45,0,88,0,42,0,139,0,26,0,30,0,221,0,68,0,168,0,113,0,130,0,252,0,16,0,0,0,232,0,36,0,0,0,108,0,118,0,117,0,175,0,77,0,227,0,144,0,0,0,0,0,66,0,221,0,0,0,236,0,72,0,123,0,142,0,0,0,233,0,40,0,30,0,0,0,32,0,223,0,88,0,92,0,180,0,216,0,173,0,0,0,214,0,174,0,180,0,163,0,221,0,0,0,212,0,96,0,0,0,46,0,59,0,58,0,174,0,51,0,56,0,0,0,178,0,0,0,0,0,147,0,226,0,0,0,133,0,181,0,193,0,0,0,18,0,0,0,232,0,13,0,0,0,202,0,50,0,0,0,0,0,151,0,207,0,31,0,173,0,0,0,186,0,0,0,34,0,0,0,162,0,144,0,41,0,34,0,228,0,0,0,162,0,0,0,135,0,0,0,29,0,189,0,233,0,248,0,0,0,166,0,170,0,131,0,0,0,111,0,0,0,221,0,171,0,122,0,144,0,0,0,208,0,23,0,172,0,134,0,239,0,98,0,19,0,129,0,188,0,14,0,235,0,242,0,69,0,0,0,0,0,0,0,108,0,170,0,0,0,0,0,57,0,129,0,0,0,0,0,0,0,34,0,0,0,65,0,50,0,29,0,188,0,220,0,236,0,251,0,70,0,230,0,105,0,15,0,225,0,127,0,119,0,150,0,116,0,227,0,0,0,141,0,103,0,124,0,166,0,96,0,148,0,0,0,81,0,73,0,250,0,0,0,86,0,45,0,41,0,141,0,137,0,11,0,0,0,94,0,52,0,206,0,44,0,0,0,78,0,168,0,0,0,100,0,53,0,203,0,48,0,100,0,205,0,200,0,57,0,170,0,118,0,0,0,107,0,0,0,0,0,166,0,139,0,224,0,184,0,214,0,233,0,0,0,216,0,116,0,108,0,139,0,99,0,219,0,12,0,179,0,0,0,103,0,53,0,0,0,70,0,150,0,2,0,151,0,183,0,99,0,183,0,213,0,89,0,223,0,138,0,250,0,0,0,95,0,30,0,58,0,206,0,192,0,205,0,82,0,34,0,0,0,161,0,201,0,211,0,0,0,0,0,32,0,72,0,0,0,40,0,3,0,0,0,32,0,210,0,196,0,0,0,141,0,24,0,0,0,239,0,66,0,18,0,194,0,168,0,77,0,55,0,177,0,0,0,135,0,131,0,53,0,130,0,243,0,151,0,242,0,123,0,52,0,6,0,168,0,213,0,0,0,158,0,49,0,0,0,0,0,156,0,146,0,42,0,200,0,115,0,84,0,124,0,0,0,63,0,146,0,60,0,0,0,0,0,116,0,0,0,111,0,0,0,91,0,233,0,0,0,58,0,191,0,0,0,205,0,161,0,35,0,0,0,105,0,234,0,96,0,31,0,191,0,0,0,231,0,194,0,32,0,33,0,9,0,95,0,48,0,0,0,0,0,238,0,0,0,142,0,157,0,147,0,152,0,36,0,0,0,92,0,109,0,81,0,35,0,165,0,0,0,140,0,155,0,44,0,5,0,0,0,186,0,210,0,24,0,75,0,246,0,99,0,20,0,0,0,0,0,0,0,191,0,144,0,166,0,15,0,12,0,219,0,253,0,0,0,15,0,0,0,213,0,55,0,109,0,75,0,0,0,204,0,194,0,0,0,60,0,153,0,148,0,0,0,0,0,68,0,84,0,207,0,5,0,123,0,0,0,86,0,244,0,49,0,216,0,36,0,59,0,31,0,217,0,32,0,81,0,119,0,137,0,237,0,112,0,189,0,17,0,0,0,7,0,0,0,103,0,0,0,0,0,226,0,56,0,0,0,32,0,0,0,245,0,34,0,160,0,69,0,150,0,17,0,119,0,227,0,202,0,0,0,171,0,219,0,42,0,208,0,148,0,218,0,181,0,0,0,94,0,4,0,10,0,128,0,1,0,187,0,159,0,171,0,90,0,172,0,58,0,137,0,202,0,0,0,172,0,250,0,37,0,49,0,210,0,100,0,59,0,0,0,0,0,0,0,221,0,217,0,33,0,230,0,3,0,246,0,48,0,88,0,163,0,14,0,92,0,0,0,132,0,162,0,176,0,103,0,0,0,41,0,190,0,126,0,0,0,68,0,161,0,0,0,0,0,132,0,72,0,67,0,18,0,109,0,218,0,0,0,0,0,60,0,175,0,204,0,254,0,80,0,150,0,135,0,245,0,212,0,11,0,94,0,0,0,0,0,31,0,238,0,12,0,27,0,200,0,117,0,173,0,10,0,92,0,180,0,26,0,41,0,172,0,94,0,0,0,91,0,255,0,187,0,78,0,59,0,0,0,77,0,24,0,96,0,0,0,157,0,140,0,124,0,126,0,179,0,200,0,35,0,0,0,0,0,93,0,36,0,124,0,161,0,247,0,71,0,104,0,239,0,67,0,216,0,0,0,77,0,0,0,151,0,138,0,236,0,214,0,0,0,2,0,103,0,215,0,249,0,9,0,191,0,0,0,0,0,172,0,35,0,4,0,0,0,0,0,156,0,149,0,194,0,0,0,125,0,189,0,227,0,228,0,159,0,168,0,116,0,131,0,23,0,50,0,0,0,104,0,0,0,179,0,0,0,206,0,33,0,0,0,191,0,0,0,185,0,49,0,187,0,224,0,12,0,41,0,205,0,51,0,234,0,161,0,161,0,0,0,228,0,0,0,110,0,182,0,176,0,33,0,130,0,137,0,0,0,72,0,210,0,177,0,224,0,41,0,106,0,180,0,246,0,29,0,61,0,203,0,0,0,0,0,26,0,70,0,80,0,115,0,0,0,242,0,92,0,39,0,0,0,193,0,0,0,147,0,79,0,24,0,0,0,160,0,234,0,40,0,0,0,215,0,208,0,0,0,104,0,0,0,155,0,12,0,131,0,250,0,0,0,0,0,0,0,177,0,146,0,7,0,0,0,213,0,45,0,0,0,84,0,210,0,0,0,17,0,185,0,16,0,58,0,176,0,0,0,112,0,33,0,224,0,183,0,166,0,0,0,87,0,43,0,0,0,97,0,75,0,97,0,187,0);
signal scenario_full  : scenario_type := (116,31,11,31,215,31,126,31,63,31,100,31,227,31,83,31,242,31,184,31,231,31,190,31,106,31,15,31,190,31,179,31,22,31,50,31,240,31,205,31,126,31,94,31,49,31,10,31,238,31,187,31,187,30,81,31,6,31,3,31,60,31,60,30,237,31,237,30,24,31,122,31,122,30,98,31,84,31,84,30,204,31,204,30,204,29,204,28,216,31,216,30,168,31,128,31,128,30,55,31,107,31,234,31,234,30,234,29,202,31,202,30,202,29,202,31,177,31,86,31,86,30,137,31,125,31,220,31,49,31,49,30,119,31,94,31,219,31,161,31,103,31,56,31,167,31,167,30,167,29,167,28,157,31,223,31,172,31,194,31,8,31,95,31,95,30,95,29,95,28,95,27,210,31,210,30,210,29,86,31,86,30,86,29,45,31,88,31,42,31,139,31,26,31,30,31,221,31,68,31,168,31,113,31,130,31,252,31,16,31,16,30,232,31,36,31,36,30,108,31,118,31,117,31,175,31,77,31,227,31,144,31,144,30,144,29,66,31,221,31,221,30,236,31,72,31,123,31,142,31,142,30,233,31,40,31,30,31,30,30,32,31,223,31,88,31,92,31,180,31,216,31,173,31,173,30,214,31,174,31,180,31,163,31,221,31,221,30,212,31,96,31,96,30,46,31,59,31,58,31,174,31,51,31,56,31,56,30,178,31,178,30,178,29,147,31,226,31,226,30,133,31,181,31,193,31,193,30,18,31,18,30,232,31,13,31,13,30,202,31,50,31,50,30,50,29,151,31,207,31,31,31,173,31,173,30,186,31,186,30,34,31,34,30,162,31,144,31,41,31,34,31,228,31,228,30,162,31,162,30,135,31,135,30,29,31,189,31,233,31,248,31,248,30,166,31,170,31,131,31,131,30,111,31,111,30,221,31,171,31,122,31,144,31,144,30,208,31,23,31,172,31,134,31,239,31,98,31,19,31,129,31,188,31,14,31,235,31,242,31,69,31,69,30,69,29,69,28,108,31,170,31,170,30,170,29,57,31,129,31,129,30,129,29,129,28,34,31,34,30,65,31,50,31,29,31,188,31,220,31,236,31,251,31,70,31,230,31,105,31,15,31,225,31,127,31,119,31,150,31,116,31,227,31,227,30,141,31,103,31,124,31,166,31,96,31,148,31,148,30,81,31,73,31,250,31,250,30,86,31,45,31,41,31,141,31,137,31,11,31,11,30,94,31,52,31,206,31,44,31,44,30,78,31,168,31,168,30,100,31,53,31,203,31,48,31,100,31,205,31,200,31,57,31,170,31,118,31,118,30,107,31,107,30,107,29,166,31,139,31,224,31,184,31,214,31,233,31,233,30,216,31,116,31,108,31,139,31,99,31,219,31,12,31,179,31,179,30,103,31,53,31,53,30,70,31,150,31,2,31,151,31,183,31,99,31,183,31,213,31,89,31,223,31,138,31,250,31,250,30,95,31,30,31,58,31,206,31,192,31,205,31,82,31,34,31,34,30,161,31,201,31,211,31,211,30,211,29,32,31,72,31,72,30,40,31,3,31,3,30,32,31,210,31,196,31,196,30,141,31,24,31,24,30,239,31,66,31,18,31,194,31,168,31,77,31,55,31,177,31,177,30,135,31,131,31,53,31,130,31,243,31,151,31,242,31,123,31,52,31,6,31,168,31,213,31,213,30,158,31,49,31,49,30,49,29,156,31,146,31,42,31,200,31,115,31,84,31,124,31,124,30,63,31,146,31,60,31,60,30,60,29,116,31,116,30,111,31,111,30,91,31,233,31,233,30,58,31,191,31,191,30,205,31,161,31,35,31,35,30,105,31,234,31,96,31,31,31,191,31,191,30,231,31,194,31,32,31,33,31,9,31,95,31,48,31,48,30,48,29,238,31,238,30,142,31,157,31,147,31,152,31,36,31,36,30,92,31,109,31,81,31,35,31,165,31,165,30,140,31,155,31,44,31,5,31,5,30,186,31,210,31,24,31,75,31,246,31,99,31,20,31,20,30,20,29,20,28,191,31,144,31,166,31,15,31,12,31,219,31,253,31,253,30,15,31,15,30,213,31,55,31,109,31,75,31,75,30,204,31,194,31,194,30,60,31,153,31,148,31,148,30,148,29,68,31,84,31,207,31,5,31,123,31,123,30,86,31,244,31,49,31,216,31,36,31,59,31,31,31,217,31,32,31,81,31,119,31,137,31,237,31,112,31,189,31,17,31,17,30,7,31,7,30,103,31,103,30,103,29,226,31,56,31,56,30,32,31,32,30,245,31,34,31,160,31,69,31,150,31,17,31,119,31,227,31,202,31,202,30,171,31,219,31,42,31,208,31,148,31,218,31,181,31,181,30,94,31,4,31,10,31,128,31,1,31,187,31,159,31,171,31,90,31,172,31,58,31,137,31,202,31,202,30,172,31,250,31,37,31,49,31,210,31,100,31,59,31,59,30,59,29,59,28,221,31,217,31,33,31,230,31,3,31,246,31,48,31,88,31,163,31,14,31,92,31,92,30,132,31,162,31,176,31,103,31,103,30,41,31,190,31,126,31,126,30,68,31,161,31,161,30,161,29,132,31,72,31,67,31,18,31,109,31,218,31,218,30,218,29,60,31,175,31,204,31,254,31,80,31,150,31,135,31,245,31,212,31,11,31,94,31,94,30,94,29,31,31,238,31,12,31,27,31,200,31,117,31,173,31,10,31,92,31,180,31,26,31,41,31,172,31,94,31,94,30,91,31,255,31,187,31,78,31,59,31,59,30,77,31,24,31,96,31,96,30,157,31,140,31,124,31,126,31,179,31,200,31,35,31,35,30,35,29,93,31,36,31,124,31,161,31,247,31,71,31,104,31,239,31,67,31,216,31,216,30,77,31,77,30,151,31,138,31,236,31,214,31,214,30,2,31,103,31,215,31,249,31,9,31,191,31,191,30,191,29,172,31,35,31,4,31,4,30,4,29,156,31,149,31,194,31,194,30,125,31,189,31,227,31,228,31,159,31,168,31,116,31,131,31,23,31,50,31,50,30,104,31,104,30,179,31,179,30,206,31,33,31,33,30,191,31,191,30,185,31,49,31,187,31,224,31,12,31,41,31,205,31,51,31,234,31,161,31,161,31,161,30,228,31,228,30,110,31,182,31,176,31,33,31,130,31,137,31,137,30,72,31,210,31,177,31,224,31,41,31,106,31,180,31,246,31,29,31,61,31,203,31,203,30,203,29,26,31,70,31,80,31,115,31,115,30,242,31,92,31,39,31,39,30,193,31,193,30,147,31,79,31,24,31,24,30,160,31,234,31,40,31,40,30,215,31,208,31,208,30,104,31,104,30,155,31,12,31,131,31,250,31,250,30,250,29,250,28,177,31,146,31,7,31,7,30,213,31,45,31,45,30,84,31,210,31,210,30,17,31,185,31,16,31,58,31,176,31,176,30,112,31,33,31,224,31,183,31,166,31,166,30,87,31,43,31,43,30,97,31,75,31,97,31,187,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
