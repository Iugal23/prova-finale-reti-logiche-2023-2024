-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_631 is
end project_tb_631;

architecture project_tb_arch_631 of project_tb_631 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 676;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (243,0,103,0,73,0,0,0,0,0,241,0,191,0,183,0,121,0,170,0,0,0,160,0,138,0,195,0,94,0,235,0,216,0,106,0,0,0,242,0,124,0,138,0,126,0,77,0,142,0,1,0,251,0,183,0,0,0,190,0,197,0,206,0,198,0,63,0,0,0,0,0,0,0,235,0,59,0,65,0,0,0,5,0,209,0,227,0,167,0,0,0,99,0,174,0,135,0,40,0,223,0,15,0,204,0,244,0,0,0,0,0,233,0,58,0,141,0,80,0,65,0,141,0,0,0,34,0,44,0,0,0,0,0,93,0,85,0,205,0,0,0,180,0,94,0,93,0,243,0,0,0,0,0,0,0,0,0,64,0,106,0,209,0,236,0,0,0,222,0,0,0,125,0,105,0,0,0,0,0,153,0,119,0,48,0,235,0,245,0,38,0,190,0,25,0,18,0,33,0,95,0,80,0,55,0,150,0,241,0,2,0,24,0,188,0,135,0,235,0,120,0,119,0,108,0,62,0,55,0,33,0,196,0,15,0,52,0,168,0,0,0,254,0,194,0,244,0,45,0,245,0,182,0,0,0,67,0,0,0,165,0,243,0,0,0,0,0,136,0,231,0,158,0,251,0,0,0,0,0,191,0,17,0,197,0,254,0,0,0,184,0,108,0,223,0,0,0,79,0,0,0,61,0,49,0,0,0,182,0,68,0,226,0,203,0,202,0,49,0,25,0,0,0,132,0,52,0,248,0,135,0,28,0,90,0,61,0,61,0,222,0,0,0,252,0,128,0,0,0,28,0,0,0,210,0,0,0,184,0,4,0,112,0,0,0,134,0,123,0,39,0,12,0,179,0,17,0,123,0,140,0,74,0,45,0,73,0,108,0,0,0,203,0,16,0,223,0,0,0,21,0,29,0,234,0,0,0,118,0,118,0,0,0,16,0,86,0,76,0,59,0,33,0,20,0,0,0,33,0,61,0,117,0,37,0,76,0,0,0,181,0,196,0,3,0,17,0,0,0,119,0,80,0,216,0,170,0,86,0,60,0,191,0,218,0,0,0,0,0,0,0,84,0,107,0,162,0,125,0,76,0,119,0,80,0,36,0,236,0,31,0,100,0,109,0,0,0,61,0,72,0,0,0,0,0,94,0,234,0,184,0,132,0,0,0,225,0,231,0,157,0,89,0,228,0,19,0,126,0,20,0,230,0,253,0,48,0,92,0,160,0,74,0,0,0,180,0,63,0,156,0,0,0,215,0,154,0,0,0,170,0,172,0,243,0,16,0,186,0,180,0,119,0,129,0,0,0,181,0,0,0,77,0,33,0,114,0,11,0,0,0,71,0,82,0,197,0,77,0,78,0,213,0,50,0,0,0,165,0,0,0,0,0,138,0,0,0,152,0,205,0,20,0,111,0,118,0,218,0,0,0,0,0,177,0,68,0,241,0,68,0,127,0,129,0,0,0,96,0,161,0,37,0,27,0,206,0,234,0,0,0,14,0,206,0,50,0,0,0,159,0,151,0,54,0,0,0,48,0,54,0,102,0,0,0,0,0,21,0,255,0,60,0,0,0,152,0,54,0,65,0,67,0,135,0,59,0,247,0,0,0,154,0,192,0,88,0,219,0,140,0,116,0,44,0,115,0,86,0,0,0,0,0,36,0,83,0,128,0,225,0,240,0,92,0,0,0,166,0,51,0,11,0,72,0,0,0,14,0,52,0,0,0,135,0,0,0,0,0,100,0,147,0,0,0,219,0,94,0,43,0,0,0,162,0,63,0,35,0,2,0,141,0,41,0,112,0,238,0,0,0,224,0,179,0,0,0,131,0,222,0,0,0,139,0,129,0,3,0,206,0,0,0,0,0,0,0,97,0,38,0,177,0,99,0,97,0,224,0,44,0,127,0,47,0,204,0,149,0,3,0,205,0,169,0,28,0,206,0,201,0,193,0,0,0,226,0,152,0,17,0,86,0,61,0,177,0,152,0,36,0,192,0,78,0,100,0,8,0,80,0,125,0,114,0,43,0,129,0,47,0,124,0,184,0,93,0,9,0,228,0,195,0,87,0,0,0,110,0,0,0,3,0,105,0,191,0,203,0,32,0,52,0,107,0,56,0,0,0,198,0,235,0,20,0,0,0,131,0,168,0,205,0,36,0,66,0,118,0,0,0,0,0,118,0,143,0,73,0,185,0,44,0,0,0,124,0,107,0,0,0,142,0,100,0,10,0,170,0,233,0,0,0,0,0,79,0,12,0,56,0,15,0,163,0,248,0,1,0,0,0,20,0,102,0,0,0,0,0,108,0,164,0,215,0,0,0,29,0,0,0,15,0,94,0,138,0,242,0,229,0,108,0,150,0,29,0,202,0,146,0,0,0,100,0,25,0,115,0,5,0,168,0,248,0,166,0,0,0,0,0,100,0,14,0,74,0,121,0,0,0,87,0,0,0,0,0,221,0,41,0,195,0,0,0,32,0,84,0,200,0,166,0,232,0,19,0,0,0,0,0,145,0,0,0,199,0,88,0,185,0,184,0,170,0,181,0,139,0,229,0,171,0,193,0,155,0,73,0,130,0,18,0,141,0,213,0,12,0,236,0,206,0,0,0,0,0,216,0,198,0,9,0,248,0,0,0,64,0,0,0,141,0,191,0,254,0,48,0,0,0,72,0,0,0,242,0,152,0,205,0,107,0,168,0,228,0,47,0,181,0,169,0,255,0,0,0,88,0,192,0,153,0,149,0,243,0,0,0,159,0,221,0,8,0,136,0,0,0,39,0,0,0,166,0,156,0,0,0,0,0,73,0,68,0,23,0,0,0,23,0,75,0,0,0,176,0,0,0,22,0,91,0,2,0,68,0,186,0,72,0,245,0,51,0,6,0,0,0,59,0,0,0,188,0,0,0,0,0,0,0,170,0,157,0,0,0,83,0,0,0,109,0,218,0,0,0,226,0,0,0,54,0,0,0,13,0,69,0,220,0,201,0,18,0,193,0,157,0,206,0,130,0,208,0,240,0,55,0,154,0,0,0,0,0,249,0,0,0,235,0);
signal scenario_full  : scenario_type := (243,31,103,31,73,31,73,30,73,29,241,31,191,31,183,31,121,31,170,31,170,30,160,31,138,31,195,31,94,31,235,31,216,31,106,31,106,30,242,31,124,31,138,31,126,31,77,31,142,31,1,31,251,31,183,31,183,30,190,31,197,31,206,31,198,31,63,31,63,30,63,29,63,28,235,31,59,31,65,31,65,30,5,31,209,31,227,31,167,31,167,30,99,31,174,31,135,31,40,31,223,31,15,31,204,31,244,31,244,30,244,29,233,31,58,31,141,31,80,31,65,31,141,31,141,30,34,31,44,31,44,30,44,29,93,31,85,31,205,31,205,30,180,31,94,31,93,31,243,31,243,30,243,29,243,28,243,27,64,31,106,31,209,31,236,31,236,30,222,31,222,30,125,31,105,31,105,30,105,29,153,31,119,31,48,31,235,31,245,31,38,31,190,31,25,31,18,31,33,31,95,31,80,31,55,31,150,31,241,31,2,31,24,31,188,31,135,31,235,31,120,31,119,31,108,31,62,31,55,31,33,31,196,31,15,31,52,31,168,31,168,30,254,31,194,31,244,31,45,31,245,31,182,31,182,30,67,31,67,30,165,31,243,31,243,30,243,29,136,31,231,31,158,31,251,31,251,30,251,29,191,31,17,31,197,31,254,31,254,30,184,31,108,31,223,31,223,30,79,31,79,30,61,31,49,31,49,30,182,31,68,31,226,31,203,31,202,31,49,31,25,31,25,30,132,31,52,31,248,31,135,31,28,31,90,31,61,31,61,31,222,31,222,30,252,31,128,31,128,30,28,31,28,30,210,31,210,30,184,31,4,31,112,31,112,30,134,31,123,31,39,31,12,31,179,31,17,31,123,31,140,31,74,31,45,31,73,31,108,31,108,30,203,31,16,31,223,31,223,30,21,31,29,31,234,31,234,30,118,31,118,31,118,30,16,31,86,31,76,31,59,31,33,31,20,31,20,30,33,31,61,31,117,31,37,31,76,31,76,30,181,31,196,31,3,31,17,31,17,30,119,31,80,31,216,31,170,31,86,31,60,31,191,31,218,31,218,30,218,29,218,28,84,31,107,31,162,31,125,31,76,31,119,31,80,31,36,31,236,31,31,31,100,31,109,31,109,30,61,31,72,31,72,30,72,29,94,31,234,31,184,31,132,31,132,30,225,31,231,31,157,31,89,31,228,31,19,31,126,31,20,31,230,31,253,31,48,31,92,31,160,31,74,31,74,30,180,31,63,31,156,31,156,30,215,31,154,31,154,30,170,31,172,31,243,31,16,31,186,31,180,31,119,31,129,31,129,30,181,31,181,30,77,31,33,31,114,31,11,31,11,30,71,31,82,31,197,31,77,31,78,31,213,31,50,31,50,30,165,31,165,30,165,29,138,31,138,30,152,31,205,31,20,31,111,31,118,31,218,31,218,30,218,29,177,31,68,31,241,31,68,31,127,31,129,31,129,30,96,31,161,31,37,31,27,31,206,31,234,31,234,30,14,31,206,31,50,31,50,30,159,31,151,31,54,31,54,30,48,31,54,31,102,31,102,30,102,29,21,31,255,31,60,31,60,30,152,31,54,31,65,31,67,31,135,31,59,31,247,31,247,30,154,31,192,31,88,31,219,31,140,31,116,31,44,31,115,31,86,31,86,30,86,29,36,31,83,31,128,31,225,31,240,31,92,31,92,30,166,31,51,31,11,31,72,31,72,30,14,31,52,31,52,30,135,31,135,30,135,29,100,31,147,31,147,30,219,31,94,31,43,31,43,30,162,31,63,31,35,31,2,31,141,31,41,31,112,31,238,31,238,30,224,31,179,31,179,30,131,31,222,31,222,30,139,31,129,31,3,31,206,31,206,30,206,29,206,28,97,31,38,31,177,31,99,31,97,31,224,31,44,31,127,31,47,31,204,31,149,31,3,31,205,31,169,31,28,31,206,31,201,31,193,31,193,30,226,31,152,31,17,31,86,31,61,31,177,31,152,31,36,31,192,31,78,31,100,31,8,31,80,31,125,31,114,31,43,31,129,31,47,31,124,31,184,31,93,31,9,31,228,31,195,31,87,31,87,30,110,31,110,30,3,31,105,31,191,31,203,31,32,31,52,31,107,31,56,31,56,30,198,31,235,31,20,31,20,30,131,31,168,31,205,31,36,31,66,31,118,31,118,30,118,29,118,31,143,31,73,31,185,31,44,31,44,30,124,31,107,31,107,30,142,31,100,31,10,31,170,31,233,31,233,30,233,29,79,31,12,31,56,31,15,31,163,31,248,31,1,31,1,30,20,31,102,31,102,30,102,29,108,31,164,31,215,31,215,30,29,31,29,30,15,31,94,31,138,31,242,31,229,31,108,31,150,31,29,31,202,31,146,31,146,30,100,31,25,31,115,31,5,31,168,31,248,31,166,31,166,30,166,29,100,31,14,31,74,31,121,31,121,30,87,31,87,30,87,29,221,31,41,31,195,31,195,30,32,31,84,31,200,31,166,31,232,31,19,31,19,30,19,29,145,31,145,30,199,31,88,31,185,31,184,31,170,31,181,31,139,31,229,31,171,31,193,31,155,31,73,31,130,31,18,31,141,31,213,31,12,31,236,31,206,31,206,30,206,29,216,31,198,31,9,31,248,31,248,30,64,31,64,30,141,31,191,31,254,31,48,31,48,30,72,31,72,30,242,31,152,31,205,31,107,31,168,31,228,31,47,31,181,31,169,31,255,31,255,30,88,31,192,31,153,31,149,31,243,31,243,30,159,31,221,31,8,31,136,31,136,30,39,31,39,30,166,31,156,31,156,30,156,29,73,31,68,31,23,31,23,30,23,31,75,31,75,30,176,31,176,30,22,31,91,31,2,31,68,31,186,31,72,31,245,31,51,31,6,31,6,30,59,31,59,30,188,31,188,30,188,29,188,28,170,31,157,31,157,30,83,31,83,30,109,31,218,31,218,30,226,31,226,30,54,31,54,30,13,31,69,31,220,31,201,31,18,31,193,31,157,31,206,31,130,31,208,31,240,31,55,31,154,31,154,30,154,29,249,31,249,30,235,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
