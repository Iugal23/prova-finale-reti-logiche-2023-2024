-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_823 is
end project_tb_823;

architecture project_tb_arch_823 of project_tb_823 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 258;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (34,0,109,0,0,0,216,0,199,0,65,0,158,0,0,0,101,0,0,0,120,0,96,0,248,0,170,0,0,0,105,0,0,0,47,0,38,0,28,0,0,0,156,0,208,0,0,0,55,0,207,0,244,0,144,0,112,0,136,0,25,0,234,0,40,0,46,0,0,0,0,0,44,0,161,0,122,0,139,0,79,0,232,0,0,0,91,0,91,0,184,0,148,0,12,0,244,0,12,0,7,0,47,0,47,0,163,0,234,0,238,0,0,0,98,0,0,0,0,0,50,0,0,0,0,0,0,0,0,0,12,0,74,0,157,0,194,0,0,0,237,0,135,0,221,0,127,0,198,0,209,0,0,0,73,0,81,0,145,0,13,0,87,0,93,0,246,0,166,0,0,0,104,0,244,0,188,0,142,0,188,0,0,0,146,0,43,0,0,0,193,0,85,0,160,0,146,0,0,0,144,0,0,0,205,0,209,0,91,0,48,0,20,0,98,0,202,0,153,0,132,0,199,0,14,0,0,0,39,0,97,0,21,0,91,0,217,0,77,0,199,0,84,0,0,0,0,0,55,0,235,0,0,0,111,0,0,0,0,0,223,0,0,0,0,0,0,0,223,0,214,0,108,0,59,0,61,0,143,0,143,0,131,0,211,0,196,0,153,0,203,0,239,0,20,0,111,0,142,0,129,0,33,0,239,0,144,0,0,0,0,0,70,0,242,0,106,0,63,0,52,0,0,0,198,0,156,0,101,0,113,0,120,0,222,0,0,0,108,0,30,0,174,0,0,0,17,0,138,0,74,0,5,0,72,0,244,0,127,0,40,0,0,0,244,0,53,0,0,0,19,0,128,0,49,0,110,0,154,0,16,0,63,0,125,0,166,0,39,0,61,0,148,0,244,0,82,0,67,0,0,0,193,0,0,0,0,0,92,0,238,0,169,0,143,0,0,0,217,0,253,0,241,0,48,0,216,0,122,0,244,0,166,0,140,0,115,0,195,0,205,0,131,0,16,0,208,0,0,0,0,0,16,0,125,0,154,0,123,0,0,0,87,0,238,0,218,0,171,0,0,0,44,0,0,0,210,0,0,0,203,0,172,0,132,0,0,0,0,0,226,0,135,0,141,0,100,0,0,0,0,0,59,0,178,0,96,0,0,0,148,0,0,0,0,0);
signal scenario_full  : scenario_type := (34,31,109,31,109,30,216,31,199,31,65,31,158,31,158,30,101,31,101,30,120,31,96,31,248,31,170,31,170,30,105,31,105,30,47,31,38,31,28,31,28,30,156,31,208,31,208,30,55,31,207,31,244,31,144,31,112,31,136,31,25,31,234,31,40,31,46,31,46,30,46,29,44,31,161,31,122,31,139,31,79,31,232,31,232,30,91,31,91,31,184,31,148,31,12,31,244,31,12,31,7,31,47,31,47,31,163,31,234,31,238,31,238,30,98,31,98,30,98,29,50,31,50,30,50,29,50,28,50,27,12,31,74,31,157,31,194,31,194,30,237,31,135,31,221,31,127,31,198,31,209,31,209,30,73,31,81,31,145,31,13,31,87,31,93,31,246,31,166,31,166,30,104,31,244,31,188,31,142,31,188,31,188,30,146,31,43,31,43,30,193,31,85,31,160,31,146,31,146,30,144,31,144,30,205,31,209,31,91,31,48,31,20,31,98,31,202,31,153,31,132,31,199,31,14,31,14,30,39,31,97,31,21,31,91,31,217,31,77,31,199,31,84,31,84,30,84,29,55,31,235,31,235,30,111,31,111,30,111,29,223,31,223,30,223,29,223,28,223,31,214,31,108,31,59,31,61,31,143,31,143,31,131,31,211,31,196,31,153,31,203,31,239,31,20,31,111,31,142,31,129,31,33,31,239,31,144,31,144,30,144,29,70,31,242,31,106,31,63,31,52,31,52,30,198,31,156,31,101,31,113,31,120,31,222,31,222,30,108,31,30,31,174,31,174,30,17,31,138,31,74,31,5,31,72,31,244,31,127,31,40,31,40,30,244,31,53,31,53,30,19,31,128,31,49,31,110,31,154,31,16,31,63,31,125,31,166,31,39,31,61,31,148,31,244,31,82,31,67,31,67,30,193,31,193,30,193,29,92,31,238,31,169,31,143,31,143,30,217,31,253,31,241,31,48,31,216,31,122,31,244,31,166,31,140,31,115,31,195,31,205,31,131,31,16,31,208,31,208,30,208,29,16,31,125,31,154,31,123,31,123,30,87,31,238,31,218,31,171,31,171,30,44,31,44,30,210,31,210,30,203,31,172,31,132,31,132,30,132,29,226,31,135,31,141,31,100,31,100,30,100,29,59,31,178,31,96,31,96,30,148,31,148,30,148,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
