-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 371;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (35,0,61,0,0,0,241,0,80,0,0,0,0,0,0,0,186,0,73,0,239,0,204,0,32,0,0,0,230,0,12,0,5,0,40,0,7,0,169,0,115,0,231,0,159,0,52,0,231,0,0,0,20,0,0,0,1,0,22,0,19,0,194,0,0,0,172,0,31,0,43,0,0,0,0,0,98,0,174,0,20,0,61,0,67,0,113,0,0,0,79,0,32,0,0,0,61,0,89,0,63,0,232,0,133,0,0,0,212,0,32,0,99,0,12,0,44,0,227,0,0,0,107,0,63,0,41,0,223,0,226,0,134,0,117,0,0,0,200,0,73,0,61,0,207,0,20,0,211,0,200,0,36,0,72,0,46,0,167,0,0,0,246,0,174,0,34,0,0,0,248,0,0,0,254,0,0,0,0,0,145,0,0,0,98,0,253,0,110,0,190,0,17,0,162,0,0,0,240,0,143,0,149,0,219,0,0,0,0,0,186,0,23,0,0,0,226,0,6,0,12,0,197,0,239,0,227,0,189,0,162,0,0,0,193,0,50,0,124,0,174,0,154,0,109,0,0,0,212,0,253,0,34,0,0,0,67,0,212,0,75,0,108,0,193,0,173,0,21,0,0,0,107,0,65,0,139,0,126,0,168,0,236,0,82,0,0,0,0,0,21,0,208,0,203,0,0,0,162,0,224,0,0,0,0,0,88,0,246,0,0,0,0,0,0,0,46,0,33,0,0,0,0,0,247,0,0,0,32,0,116,0,237,0,119,0,63,0,15,0,0,0,82,0,187,0,218,0,0,0,0,0,255,0,86,0,126,0,112,0,96,0,211,0,6,0,8,0,0,0,0,0,16,0,239,0,203,0,214,0,81,0,144,0,152,0,252,0,247,0,245,0,69,0,54,0,0,0,123,0,208,0,195,0,213,0,0,0,94,0,137,0,193,0,0,0,128,0,222,0,0,0,143,0,100,0,10,0,0,0,49,0,38,0,106,0,233,0,237,0,197,0,106,0,0,0,0,0,139,0,77,0,102,0,214,0,58,0,221,0,38,0,139,0,93,0,0,0,0,0,242,0,128,0,214,0,0,0,0,0,0,0,34,0,0,0,111,0,0,0,2,0,47,0,118,0,0,0,0,0,244,0,0,0,238,0,228,0,36,0,0,0,0,0,101,0,0,0,0,0,0,0,0,0,178,0,0,0,0,0,228,0,246,0,36,0,0,0,0,0,217,0,227,0,160,0,168,0,107,0,241,0,0,0,224,0,61,0,0,0,109,0,0,0,158,0,200,0,160,0,227,0,0,0,130,0,113,0,239,0,91,0,0,0,190,0,207,0,66,0,0,0,0,0,155,0,99,0,246,0,174,0,163,0,0,0,131,0,132,0,96,0,21,0,0,0,236,0,200,0,233,0,167,0,123,0,179,0,0,0,29,0,0,0,233,0,11,0,148,0,43,0,194,0,31,0,162,0,147,0,145,0,101,0,244,0,28,0,240,0,129,0,252,0,214,0,68,0,0,0,0,0,141,0,0,0,109,0,0,0,117,0,0,0,116,0,108,0,0,0,139,0,78,0,0,0,64,0,226,0,169,0,112,0,251,0,101,0,0,0,205,0,140,0,204,0,240,0,0,0,0,0,88,0,105,0,41,0,0,0,0,0,0,0,39,0,219,0,99,0,0,0);
signal scenario_full  : scenario_type := (35,31,61,31,61,30,241,31,80,31,80,30,80,29,80,28,186,31,73,31,239,31,204,31,32,31,32,30,230,31,12,31,5,31,40,31,7,31,169,31,115,31,231,31,159,31,52,31,231,31,231,30,20,31,20,30,1,31,22,31,19,31,194,31,194,30,172,31,31,31,43,31,43,30,43,29,98,31,174,31,20,31,61,31,67,31,113,31,113,30,79,31,32,31,32,30,61,31,89,31,63,31,232,31,133,31,133,30,212,31,32,31,99,31,12,31,44,31,227,31,227,30,107,31,63,31,41,31,223,31,226,31,134,31,117,31,117,30,200,31,73,31,61,31,207,31,20,31,211,31,200,31,36,31,72,31,46,31,167,31,167,30,246,31,174,31,34,31,34,30,248,31,248,30,254,31,254,30,254,29,145,31,145,30,98,31,253,31,110,31,190,31,17,31,162,31,162,30,240,31,143,31,149,31,219,31,219,30,219,29,186,31,23,31,23,30,226,31,6,31,12,31,197,31,239,31,227,31,189,31,162,31,162,30,193,31,50,31,124,31,174,31,154,31,109,31,109,30,212,31,253,31,34,31,34,30,67,31,212,31,75,31,108,31,193,31,173,31,21,31,21,30,107,31,65,31,139,31,126,31,168,31,236,31,82,31,82,30,82,29,21,31,208,31,203,31,203,30,162,31,224,31,224,30,224,29,88,31,246,31,246,30,246,29,246,28,46,31,33,31,33,30,33,29,247,31,247,30,32,31,116,31,237,31,119,31,63,31,15,31,15,30,82,31,187,31,218,31,218,30,218,29,255,31,86,31,126,31,112,31,96,31,211,31,6,31,8,31,8,30,8,29,16,31,239,31,203,31,214,31,81,31,144,31,152,31,252,31,247,31,245,31,69,31,54,31,54,30,123,31,208,31,195,31,213,31,213,30,94,31,137,31,193,31,193,30,128,31,222,31,222,30,143,31,100,31,10,31,10,30,49,31,38,31,106,31,233,31,237,31,197,31,106,31,106,30,106,29,139,31,77,31,102,31,214,31,58,31,221,31,38,31,139,31,93,31,93,30,93,29,242,31,128,31,214,31,214,30,214,29,214,28,34,31,34,30,111,31,111,30,2,31,47,31,118,31,118,30,118,29,244,31,244,30,238,31,228,31,36,31,36,30,36,29,101,31,101,30,101,29,101,28,101,27,178,31,178,30,178,29,228,31,246,31,36,31,36,30,36,29,217,31,227,31,160,31,168,31,107,31,241,31,241,30,224,31,61,31,61,30,109,31,109,30,158,31,200,31,160,31,227,31,227,30,130,31,113,31,239,31,91,31,91,30,190,31,207,31,66,31,66,30,66,29,155,31,99,31,246,31,174,31,163,31,163,30,131,31,132,31,96,31,21,31,21,30,236,31,200,31,233,31,167,31,123,31,179,31,179,30,29,31,29,30,233,31,11,31,148,31,43,31,194,31,31,31,162,31,147,31,145,31,101,31,244,31,28,31,240,31,129,31,252,31,214,31,68,31,68,30,68,29,141,31,141,30,109,31,109,30,117,31,117,30,116,31,108,31,108,30,139,31,78,31,78,30,64,31,226,31,169,31,112,31,251,31,101,31,101,30,205,31,140,31,204,31,240,31,240,30,240,29,88,31,105,31,41,31,41,30,41,29,41,28,39,31,219,31,99,31,99,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
