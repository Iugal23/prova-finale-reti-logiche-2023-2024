-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 544;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (255,0,144,0,0,0,78,0,0,0,0,0,110,0,59,0,180,0,236,0,150,0,0,0,92,0,122,0,135,0,0,0,0,0,14,0,173,0,230,0,27,0,63,0,0,0,119,0,127,0,90,0,200,0,101,0,0,0,74,0,191,0,145,0,104,0,154,0,0,0,68,0,39,0,12,0,121,0,86,0,216,0,179,0,0,0,8,0,193,0,207,0,117,0,26,0,127,0,14,0,159,0,193,0,104,0,128,0,132,0,117,0,84,0,89,0,0,0,11,0,39,0,0,0,233,0,197,0,175,0,11,0,0,0,92,0,83,0,94,0,0,0,170,0,238,0,128,0,4,0,205,0,40,0,249,0,208,0,61,0,172,0,80,0,0,0,0,0,92,0,0,0,0,0,0,0,49,0,156,0,181,0,105,0,0,0,138,0,213,0,0,0,190,0,227,0,0,0,25,0,60,0,41,0,11,0,253,0,100,0,116,0,121,0,77,0,102,0,225,0,42,0,226,0,119,0,125,0,25,0,0,0,0,0,173,0,0,0,0,0,0,0,80,0,87,0,127,0,171,0,42,0,0,0,128,0,176,0,160,0,60,0,153,0,0,0,48,0,63,0,161,0,207,0,130,0,110,0,105,0,230,0,78,0,198,0,194,0,171,0,43,0,48,0,156,0,19,0,0,0,251,0,195,0,220,0,145,0,184,0,70,0,187,0,82,0,0,0,94,0,106,0,70,0,160,0,216,0,53,0,231,0,0,0,85,0,205,0,80,0,62,0,226,0,202,0,0,0,136,0,43,0,71,0,0,0,232,0,177,0,37,0,138,0,129,0,28,0,16,0,18,0,112,0,55,0,0,0,32,0,144,0,11,0,226,0,218,0,0,0,166,0,0,0,59,0,216,0,116,0,136,0,2,0,39,0,252,0,224,0,201,0,0,0,195,0,29,0,0,0,16,0,196,0,244,0,9,0,126,0,14,0,189,0,0,0,105,0,103,0,8,0,74,0,182,0,125,0,98,0,0,0,14,0,58,0,26,0,74,0,0,0,122,0,112,0,88,0,0,0,102,0,240,0,41,0,96,0,75,0,185,0,207,0,227,0,178,0,103,0,0,0,0,0,0,0,135,0,198,0,102,0,198,0,245,0,0,0,163,0,150,0,0,0,221,0,95,0,0,0,185,0,83,0,0,0,0,0,0,0,50,0,18,0,86,0,206,0,124,0,86,0,0,0,166,0,0,0,185,0,245,0,16,0,217,0,20,0,152,0,41,0,193,0,0,0,186,0,19,0,0,0,252,0,187,0,203,0,41,0,37,0,86,0,0,0,118,0,34,0,190,0,100,0,19,0,70,0,57,0,8,0,102,0,176,0,22,0,23,0,7,0,212,0,0,0,78,0,247,0,0,0,6,0,195,0,0,0,64,0,0,0,12,0,47,0,19,0,30,0,8,0,29,0,18,0,73,0,109,0,0,0,97,0,208,0,78,0,3,0,0,0,194,0,0,0,152,0,191,0,0,0,38,0,162,0,98,0,0,0,58,0,0,0,0,0,0,0,135,0,181,0,236,0,232,0,61,0,239,0,195,0,0,0,22,0,107,0,40,0,158,0,0,0,229,0,0,0,94,0,0,0,252,0,101,0,185,0,73,0,100,0,70,0,197,0,194,0,36,0,246,0,0,0,62,0,228,0,19,0,210,0,84,0,106,0,106,0,89,0,219,0,0,0,239,0,181,0,169,0,141,0,158,0,141,0,0,0,60,0,185,0,149,0,12,0,150,0,69,0,42,0,24,0,131,0,254,0,220,0,0,0,221,0,101,0,154,0,0,0,0,0,0,0,0,0,233,0,70,0,167,0,246,0,174,0,52,0,173,0,135,0,0,0,151,0,146,0,160,0,38,0,47,0,193,0,96,0,0,0,0,0,109,0,3,0,246,0,193,0,0,0,87,0,0,0,18,0,66,0,74,0,100,0,4,0,36,0,188,0,101,0,0,0,217,0,0,0,0,0,101,0,174,0,236,0,220,0,101,0,58,0,240,0,145,0,194,0,0,0,0,0,69,0,205,0,137,0,69,0,137,0,243,0,0,0,0,0,114,0,99,0,162,0,1,0,183,0,191,0,250,0,0,0,255,0,176,0,239,0,0,0,0,0,157,0,173,0,156,0,9,0,91,0,177,0,76,0,213,0,0,0,0,0,0,0,0,0,80,0,14,0,222,0,0,0,58,0,151,0,156,0,145,0,0,0,0,0,123,0,134,0,252,0,0,0,24,0,172,0,58,0,186,0,93,0,218,0,158,0,214,0,0,0,199,0,165,0,115,0,53,0,72,0,19,0,0,0,39,0,183,0,206,0,146,0,0,0,4,0,94,0,138,0,0,0,0,0,141,0,32,0,255,0,6,0,176,0,89,0,219,0,0,0,196,0,0,0,0,0,255,0,95,0,0,0,121,0);
signal scenario_full  : scenario_type := (255,31,144,31,144,30,78,31,78,30,78,29,110,31,59,31,180,31,236,31,150,31,150,30,92,31,122,31,135,31,135,30,135,29,14,31,173,31,230,31,27,31,63,31,63,30,119,31,127,31,90,31,200,31,101,31,101,30,74,31,191,31,145,31,104,31,154,31,154,30,68,31,39,31,12,31,121,31,86,31,216,31,179,31,179,30,8,31,193,31,207,31,117,31,26,31,127,31,14,31,159,31,193,31,104,31,128,31,132,31,117,31,84,31,89,31,89,30,11,31,39,31,39,30,233,31,197,31,175,31,11,31,11,30,92,31,83,31,94,31,94,30,170,31,238,31,128,31,4,31,205,31,40,31,249,31,208,31,61,31,172,31,80,31,80,30,80,29,92,31,92,30,92,29,92,28,49,31,156,31,181,31,105,31,105,30,138,31,213,31,213,30,190,31,227,31,227,30,25,31,60,31,41,31,11,31,253,31,100,31,116,31,121,31,77,31,102,31,225,31,42,31,226,31,119,31,125,31,25,31,25,30,25,29,173,31,173,30,173,29,173,28,80,31,87,31,127,31,171,31,42,31,42,30,128,31,176,31,160,31,60,31,153,31,153,30,48,31,63,31,161,31,207,31,130,31,110,31,105,31,230,31,78,31,198,31,194,31,171,31,43,31,48,31,156,31,19,31,19,30,251,31,195,31,220,31,145,31,184,31,70,31,187,31,82,31,82,30,94,31,106,31,70,31,160,31,216,31,53,31,231,31,231,30,85,31,205,31,80,31,62,31,226,31,202,31,202,30,136,31,43,31,71,31,71,30,232,31,177,31,37,31,138,31,129,31,28,31,16,31,18,31,112,31,55,31,55,30,32,31,144,31,11,31,226,31,218,31,218,30,166,31,166,30,59,31,216,31,116,31,136,31,2,31,39,31,252,31,224,31,201,31,201,30,195,31,29,31,29,30,16,31,196,31,244,31,9,31,126,31,14,31,189,31,189,30,105,31,103,31,8,31,74,31,182,31,125,31,98,31,98,30,14,31,58,31,26,31,74,31,74,30,122,31,112,31,88,31,88,30,102,31,240,31,41,31,96,31,75,31,185,31,207,31,227,31,178,31,103,31,103,30,103,29,103,28,135,31,198,31,102,31,198,31,245,31,245,30,163,31,150,31,150,30,221,31,95,31,95,30,185,31,83,31,83,30,83,29,83,28,50,31,18,31,86,31,206,31,124,31,86,31,86,30,166,31,166,30,185,31,245,31,16,31,217,31,20,31,152,31,41,31,193,31,193,30,186,31,19,31,19,30,252,31,187,31,203,31,41,31,37,31,86,31,86,30,118,31,34,31,190,31,100,31,19,31,70,31,57,31,8,31,102,31,176,31,22,31,23,31,7,31,212,31,212,30,78,31,247,31,247,30,6,31,195,31,195,30,64,31,64,30,12,31,47,31,19,31,30,31,8,31,29,31,18,31,73,31,109,31,109,30,97,31,208,31,78,31,3,31,3,30,194,31,194,30,152,31,191,31,191,30,38,31,162,31,98,31,98,30,58,31,58,30,58,29,58,28,135,31,181,31,236,31,232,31,61,31,239,31,195,31,195,30,22,31,107,31,40,31,158,31,158,30,229,31,229,30,94,31,94,30,252,31,101,31,185,31,73,31,100,31,70,31,197,31,194,31,36,31,246,31,246,30,62,31,228,31,19,31,210,31,84,31,106,31,106,31,89,31,219,31,219,30,239,31,181,31,169,31,141,31,158,31,141,31,141,30,60,31,185,31,149,31,12,31,150,31,69,31,42,31,24,31,131,31,254,31,220,31,220,30,221,31,101,31,154,31,154,30,154,29,154,28,154,27,233,31,70,31,167,31,246,31,174,31,52,31,173,31,135,31,135,30,151,31,146,31,160,31,38,31,47,31,193,31,96,31,96,30,96,29,109,31,3,31,246,31,193,31,193,30,87,31,87,30,18,31,66,31,74,31,100,31,4,31,36,31,188,31,101,31,101,30,217,31,217,30,217,29,101,31,174,31,236,31,220,31,101,31,58,31,240,31,145,31,194,31,194,30,194,29,69,31,205,31,137,31,69,31,137,31,243,31,243,30,243,29,114,31,99,31,162,31,1,31,183,31,191,31,250,31,250,30,255,31,176,31,239,31,239,30,239,29,157,31,173,31,156,31,9,31,91,31,177,31,76,31,213,31,213,30,213,29,213,28,213,27,80,31,14,31,222,31,222,30,58,31,151,31,156,31,145,31,145,30,145,29,123,31,134,31,252,31,252,30,24,31,172,31,58,31,186,31,93,31,218,31,158,31,214,31,214,30,199,31,165,31,115,31,53,31,72,31,19,31,19,30,39,31,183,31,206,31,146,31,146,30,4,31,94,31,138,31,138,30,138,29,141,31,32,31,255,31,6,31,176,31,89,31,219,31,219,30,196,31,196,30,196,29,255,31,95,31,95,30,121,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
