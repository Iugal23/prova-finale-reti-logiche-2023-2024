-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_229 is
end project_tb_229;

architecture project_tb_arch_229 of project_tb_229 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 586;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,62,0,133,0,194,0,47,0,223,0,128,0,56,0,198,0,120,0,14,0,0,0,0,0,239,0,0,0,104,0,0,0,98,0,0,0,104,0,54,0,185,0,113,0,95,0,175,0,101,0,27,0,85,0,250,0,220,0,124,0,96,0,239,0,0,0,0,0,0,0,0,0,69,0,193,0,229,0,104,0,22,0,2,0,23,0,249,0,2,0,66,0,16,0,0,0,40,0,37,0,25,0,210,0,155,0,45,0,202,0,9,0,9,0,150,0,182,0,27,0,0,0,232,0,192,0,0,0,73,0,6,0,0,0,0,0,90,0,56,0,7,0,243,0,253,0,180,0,0,0,0,0,250,0,0,0,106,0,99,0,45,0,245,0,102,0,144,0,0,0,77,0,224,0,105,0,211,0,51,0,46,0,0,0,8,0,0,0,115,0,73,0,63,0,216,0,0,0,0,0,132,0,11,0,228,0,0,0,175,0,164,0,123,0,43,0,36,0,92,0,87,0,254,0,133,0,253,0,244,0,0,0,33,0,0,0,137,0,0,0,0,0,48,0,1,0,66,0,96,0,142,0,141,0,15,0,175,0,206,0,27,0,0,0,138,0,107,0,0,0,0,0,184,0,64,0,0,0,10,0,52,0,0,0,106,0,181,0,58,0,24,0,134,0,56,0,69,0,6,0,201,0,0,0,0,0,133,0,57,0,145,0,219,0,145,0,229,0,120,0,67,0,195,0,198,0,4,0,82,0,117,0,207,0,115,0,40,0,11,0,153,0,5,0,189,0,138,0,13,0,6,0,114,0,32,0,218,0,0,0,77,0,212,0,140,0,71,0,115,0,25,0,208,0,197,0,75,0,35,0,128,0,0,0,114,0,247,0,0,0,170,0,210,0,228,0,42,0,74,0,224,0,234,0,184,0,0,0,7,0,100,0,230,0,100,0,220,0,38,0,39,0,63,0,0,0,29,0,18,0,219,0,69,0,126,0,0,0,0,0,61,0,193,0,205,0,0,0,27,0,147,0,204,0,186,0,98,0,236,0,17,0,188,0,0,0,0,0,42,0,57,0,122,0,98,0,221,0,0,0,26,0,116,0,66,0,168,0,229,0,236,0,11,0,195,0,251,0,102,0,101,0,237,0,0,0,121,0,108,0,144,0,42,0,11,0,222,0,253,0,109,0,216,0,239,0,201,0,176,0,0,0,48,0,253,0,194,0,235,0,0,0,10,0,0,0,0,0,131,0,0,0,0,0,96,0,0,0,149,0,104,0,111,0,135,0,96,0,157,0,55,0,228,0,171,0,102,0,221,0,167,0,0,0,155,0,0,0,212,0,229,0,0,0,133,0,3,0,0,0,87,0,67,0,177,0,249,0,17,0,0,0,181,0,59,0,109,0,143,0,109,0,0,0,96,0,0,0,177,0,0,0,83,0,81,0,115,0,207,0,0,0,0,0,195,0,0,0,184,0,0,0,189,0,174,0,0,0,88,0,62,0,31,0,178,0,69,0,176,0,0,0,69,0,37,0,187,0,0,0,244,0,120,0,57,0,215,0,0,0,167,0,0,0,255,0,77,0,0,0,0,0,169,0,35,0,161,0,0,0,88,0,13,0,191,0,95,0,169,0,66,0,94,0,0,0,73,0,216,0,228,0,215,0,70,0,115,0,112,0,117,0,105,0,169,0,0,0,151,0,181,0,123,0,0,0,11,0,10,0,234,0,132,0,151,0,0,0,130,0,223,0,9,0,158,0,0,0,0,0,108,0,237,0,68,0,42,0,84,0,0,0,135,0,87,0,212,0,144,0,106,0,23,0,0,0,211,0,211,0,0,0,252,0,0,0,70,0,85,0,42,0,59,0,0,0,0,0,54,0,179,0,111,0,98,0,29,0,165,0,230,0,161,0,227,0,160,0,0,0,59,0,9,0,172,0,69,0,0,0,243,0,0,0,252,0,229,0,55,0,66,0,186,0,199,0,95,0,170,0,0,0,168,0,140,0,18,0,0,0,70,0,134,0,44,0,138,0,156,0,218,0,104,0,0,0,131,0,68,0,0,0,44,0,0,0,104,0,60,0,199,0,225,0,243,0,0,0,236,0,149,0,0,0,4,0,66,0,168,0,0,0,190,0,0,0,38,0,135,0,234,0,86,0,55,0,0,0,180,0,0,0,185,0,3,0,19,0,106,0,0,0,171,0,71,0,151,0,110,0,12,0,222,0,201,0,0,0,159,0,167,0,0,0,34,0,30,0,109,0,0,0,239,0,222,0,27,0,155,0,194,0,38,0,23,0,190,0,231,0,255,0,198,0,130,0,120,0,110,0,139,0,224,0,75,0,218,0,52,0,232,0,0,0,225,0,26,0,0,0,173,0,86,0,240,0,0,0,241,0,122,0,204,0,7,0,192,0,82,0,236,0,118,0,0,0,0,0,0,0,0,0,0,0,56,0,154,0,0,0,10,0,234,0,112,0,23,0,189,0,33,0,171,0,79,0,217,0,194,0,201,0,158,0,141,0,0,0,0,0,0,0,167,0,50,0,102,0,0,0,6,0,2,0,237,0,0,0,161,0,0,0,22,0,183,0,65,0,0,0,120,0,146,0,102,0,82,0,111,0,0,0,0,0,66,0,143,0,33,0);
signal scenario_full  : scenario_type := (0,0,62,31,133,31,194,31,47,31,223,31,128,31,56,31,198,31,120,31,14,31,14,30,14,29,239,31,239,30,104,31,104,30,98,31,98,30,104,31,54,31,185,31,113,31,95,31,175,31,101,31,27,31,85,31,250,31,220,31,124,31,96,31,239,31,239,30,239,29,239,28,239,27,69,31,193,31,229,31,104,31,22,31,2,31,23,31,249,31,2,31,66,31,16,31,16,30,40,31,37,31,25,31,210,31,155,31,45,31,202,31,9,31,9,31,150,31,182,31,27,31,27,30,232,31,192,31,192,30,73,31,6,31,6,30,6,29,90,31,56,31,7,31,243,31,253,31,180,31,180,30,180,29,250,31,250,30,106,31,99,31,45,31,245,31,102,31,144,31,144,30,77,31,224,31,105,31,211,31,51,31,46,31,46,30,8,31,8,30,115,31,73,31,63,31,216,31,216,30,216,29,132,31,11,31,228,31,228,30,175,31,164,31,123,31,43,31,36,31,92,31,87,31,254,31,133,31,253,31,244,31,244,30,33,31,33,30,137,31,137,30,137,29,48,31,1,31,66,31,96,31,142,31,141,31,15,31,175,31,206,31,27,31,27,30,138,31,107,31,107,30,107,29,184,31,64,31,64,30,10,31,52,31,52,30,106,31,181,31,58,31,24,31,134,31,56,31,69,31,6,31,201,31,201,30,201,29,133,31,57,31,145,31,219,31,145,31,229,31,120,31,67,31,195,31,198,31,4,31,82,31,117,31,207,31,115,31,40,31,11,31,153,31,5,31,189,31,138,31,13,31,6,31,114,31,32,31,218,31,218,30,77,31,212,31,140,31,71,31,115,31,25,31,208,31,197,31,75,31,35,31,128,31,128,30,114,31,247,31,247,30,170,31,210,31,228,31,42,31,74,31,224,31,234,31,184,31,184,30,7,31,100,31,230,31,100,31,220,31,38,31,39,31,63,31,63,30,29,31,18,31,219,31,69,31,126,31,126,30,126,29,61,31,193,31,205,31,205,30,27,31,147,31,204,31,186,31,98,31,236,31,17,31,188,31,188,30,188,29,42,31,57,31,122,31,98,31,221,31,221,30,26,31,116,31,66,31,168,31,229,31,236,31,11,31,195,31,251,31,102,31,101,31,237,31,237,30,121,31,108,31,144,31,42,31,11,31,222,31,253,31,109,31,216,31,239,31,201,31,176,31,176,30,48,31,253,31,194,31,235,31,235,30,10,31,10,30,10,29,131,31,131,30,131,29,96,31,96,30,149,31,104,31,111,31,135,31,96,31,157,31,55,31,228,31,171,31,102,31,221,31,167,31,167,30,155,31,155,30,212,31,229,31,229,30,133,31,3,31,3,30,87,31,67,31,177,31,249,31,17,31,17,30,181,31,59,31,109,31,143,31,109,31,109,30,96,31,96,30,177,31,177,30,83,31,81,31,115,31,207,31,207,30,207,29,195,31,195,30,184,31,184,30,189,31,174,31,174,30,88,31,62,31,31,31,178,31,69,31,176,31,176,30,69,31,37,31,187,31,187,30,244,31,120,31,57,31,215,31,215,30,167,31,167,30,255,31,77,31,77,30,77,29,169,31,35,31,161,31,161,30,88,31,13,31,191,31,95,31,169,31,66,31,94,31,94,30,73,31,216,31,228,31,215,31,70,31,115,31,112,31,117,31,105,31,169,31,169,30,151,31,181,31,123,31,123,30,11,31,10,31,234,31,132,31,151,31,151,30,130,31,223,31,9,31,158,31,158,30,158,29,108,31,237,31,68,31,42,31,84,31,84,30,135,31,87,31,212,31,144,31,106,31,23,31,23,30,211,31,211,31,211,30,252,31,252,30,70,31,85,31,42,31,59,31,59,30,59,29,54,31,179,31,111,31,98,31,29,31,165,31,230,31,161,31,227,31,160,31,160,30,59,31,9,31,172,31,69,31,69,30,243,31,243,30,252,31,229,31,55,31,66,31,186,31,199,31,95,31,170,31,170,30,168,31,140,31,18,31,18,30,70,31,134,31,44,31,138,31,156,31,218,31,104,31,104,30,131,31,68,31,68,30,44,31,44,30,104,31,60,31,199,31,225,31,243,31,243,30,236,31,149,31,149,30,4,31,66,31,168,31,168,30,190,31,190,30,38,31,135,31,234,31,86,31,55,31,55,30,180,31,180,30,185,31,3,31,19,31,106,31,106,30,171,31,71,31,151,31,110,31,12,31,222,31,201,31,201,30,159,31,167,31,167,30,34,31,30,31,109,31,109,30,239,31,222,31,27,31,155,31,194,31,38,31,23,31,190,31,231,31,255,31,198,31,130,31,120,31,110,31,139,31,224,31,75,31,218,31,52,31,232,31,232,30,225,31,26,31,26,30,173,31,86,31,240,31,240,30,241,31,122,31,204,31,7,31,192,31,82,31,236,31,118,31,118,30,118,29,118,28,118,27,118,26,56,31,154,31,154,30,10,31,234,31,112,31,23,31,189,31,33,31,171,31,79,31,217,31,194,31,201,31,158,31,141,31,141,30,141,29,141,28,167,31,50,31,102,31,102,30,6,31,2,31,237,31,237,30,161,31,161,30,22,31,183,31,65,31,65,30,120,31,146,31,102,31,82,31,111,31,111,30,111,29,66,31,143,31,33,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
