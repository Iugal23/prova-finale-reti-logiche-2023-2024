-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 689;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (62,0,51,0,0,0,228,0,167,0,0,0,11,0,88,0,69,0,104,0,160,0,196,0,150,0,0,0,0,0,82,0,64,0,2,0,17,0,21,0,214,0,27,0,35,0,249,0,222,0,76,0,148,0,221,0,137,0,118,0,158,0,250,0,243,0,179,0,0,0,251,0,98,0,235,0,2,0,124,0,225,0,77,0,137,0,152,0,125,0,201,0,65,0,106,0,103,0,214,0,0,0,40,0,193,0,207,0,238,0,178,0,38,0,201,0,16,0,0,0,52,0,18,0,232,0,64,0,198,0,193,0,0,0,72,0,0,0,0,0,53,0,221,0,205,0,0,0,236,0,32,0,3,0,151,0,115,0,235,0,116,0,0,0,154,0,0,0,57,0,14,0,248,0,0,0,14,0,0,0,0,0,0,0,207,0,251,0,222,0,0,0,0,0,50,0,13,0,161,0,198,0,23,0,62,0,58,0,76,0,134,0,0,0,0,0,0,0,0,0,39,0,232,0,157,0,118,0,0,0,233,0,75,0,0,0,237,0,0,0,36,0,21,0,0,0,222,0,122,0,250,0,188,0,165,0,58,0,251,0,218,0,191,0,193,0,2,0,60,0,175,0,254,0,194,0,144,0,15,0,0,0,92,0,85,0,178,0,186,0,0,0,86,0,127,0,8,0,12,0,0,0,0,0,0,0,173,0,27,0,151,0,227,0,80,0,169,0,176,0,0,0,34,0,55,0,151,0,0,0,132,0,124,0,90,0,0,0,176,0,22,0,188,0,67,0,116,0,48,0,72,0,0,0,0,0,218,0,111,0,225,0,232,0,95,0,0,0,0,0,169,0,119,0,76,0,118,0,199,0,136,0,255,0,120,0,0,0,17,0,157,0,42,0,13,0,237,0,142,0,198,0,201,0,122,0,194,0,40,0,0,0,162,0,2,0,133,0,154,0,71,0,225,0,238,0,3,0,112,0,233,0,121,0,33,0,65,0,108,0,131,0,205,0,197,0,220,0,100,0,59,0,92,0,161,0,178,0,74,0,28,0,192,0,55,0,191,0,211,0,111,0,112,0,0,0,78,0,155,0,195,0,0,0,225,0,0,0,104,0,192,0,105,0,12,0,20,0,161,0,35,0,174,0,138,0,159,0,0,0,182,0,0,0,116,0,61,0,17,0,1,0,0,0,138,0,126,0,144,0,172,0,218,0,13,0,107,0,195,0,4,0,0,0,185,0,210,0,0,0,0,0,17,0,92,0,205,0,6,0,249,0,195,0,212,0,135,0,28,0,89,0,116,0,215,0,0,0,125,0,15,0,0,0,0,0,218,0,250,0,197,0,124,0,122,0,33,0,0,0,0,0,137,0,0,0,253,0,116,0,234,0,161,0,109,0,0,0,0,0,0,0,175,0,59,0,0,0,219,0,45,0,0,0,96,0,0,0,10,0,122,0,10,0,118,0,245,0,99,0,246,0,49,0,181,0,204,0,214,0,173,0,0,0,62,0,182,0,135,0,26,0,0,0,225,0,0,0,27,0,0,0,120,0,144,0,0,0,168,0,137,0,9,0,235,0,146,0,205,0,162,0,0,0,239,0,149,0,77,0,33,0,98,0,18,0,0,0,158,0,0,0,0,0,0,0,2,0,35,0,29,0,26,0,54,0,87,0,21,0,254,0,212,0,0,0,0,0,224,0,4,0,153,0,0,0,129,0,241,0,106,0,178,0,97,0,101,0,0,0,0,0,191,0,149,0,80,0,217,0,194,0,145,0,199,0,118,0,75,0,238,0,191,0,0,0,107,0,52,0,7,0,188,0,64,0,0,0,0,0,93,0,121,0,47,0,108,0,0,0,71,0,98,0,168,0,214,0,0,0,0,0,132,0,97,0,0,0,136,0,193,0,130,0,28,0,0,0,118,0,157,0,42,0,118,0,82,0,0,0,167,0,149,0,250,0,127,0,42,0,2,0,0,0,119,0,0,0,78,0,198,0,107,0,113,0,60,0,13,0,0,0,106,0,109,0,56,0,94,0,206,0,231,0,1,0,182,0,221,0,0,0,26,0,219,0,221,0,153,0,31,0,6,0,111,0,239,0,0,0,131,0,77,0,211,0,49,0,137,0,113,0,91,0,214,0,22,0,171,0,0,0,0,0,201,0,94,0,245,0,58,0,249,0,22,0,227,0,215,0,47,0,208,0,0,0,40,0,0,0,0,0,238,0,122,0,86,0,0,0,19,0,51,0,157,0,227,0,0,0,155,0,179,0,133,0,23,0,78,0,0,0,242,0,238,0,254,0,63,0,174,0,81,0,163,0,225,0,46,0,30,0,22,0,209,0,252,0,252,0,0,0,189,0,0,0,233,0,122,0,42,0,148,0,162,0,64,0,0,0,61,0,0,0,191,0,144,0,81,0,234,0,114,0,0,0,242,0,229,0,0,0,247,0,0,0,205,0,31,0,247,0,156,0,136,0,141,0,0,0,225,0,114,0,11,0,144,0,0,0,0,0,17,0,227,0,203,0,145,0,41,0,0,0,193,0,141,0,42,0,114,0,26,0,0,0,0,0,0,0,60,0,182,0,177,0,207,0,182,0,0,0,3,0,104,0,152,0,155,0,94,0,0,0,187,0,47,0,75,0,217,0,40,0,132,0,0,0,0,0,0,0,81,0,124,0,248,0,74,0,0,0,37,0,0,0,10,0,250,0,243,0,231,0,81,0,65,0,0,0,42,0,181,0,150,0,243,0,0,0,179,0,83,0,0,0,237,0,166,0,0,0,54,0,204,0,71,0,219,0,0,0,0,0,0,0,11,0,26,0,162,0,21,0,0,0,0,0,0,0,35,0,21,0,163,0,0,0,211,0,100,0,0,0,231,0,101,0,246,0,0,0,229,0,215,0,127,0,202,0,234,0,216,0,12,0,85,0,1,0,60,0,182,0,98,0,48,0,227,0,218,0,0,0,55,0,1,0,91,0,221,0,219,0,195,0,108,0,172,0,0,0,0,0,0,0,223,0,0,0,25,0,244,0,230,0,0,0,34,0,58,0,26,0,41,0,114,0,0,0,0,0,68,0,0,0,0,0,141,0,164,0,189,0,0,0,40,0);
signal scenario_full  : scenario_type := (62,31,51,31,51,30,228,31,167,31,167,30,11,31,88,31,69,31,104,31,160,31,196,31,150,31,150,30,150,29,82,31,64,31,2,31,17,31,21,31,214,31,27,31,35,31,249,31,222,31,76,31,148,31,221,31,137,31,118,31,158,31,250,31,243,31,179,31,179,30,251,31,98,31,235,31,2,31,124,31,225,31,77,31,137,31,152,31,125,31,201,31,65,31,106,31,103,31,214,31,214,30,40,31,193,31,207,31,238,31,178,31,38,31,201,31,16,31,16,30,52,31,18,31,232,31,64,31,198,31,193,31,193,30,72,31,72,30,72,29,53,31,221,31,205,31,205,30,236,31,32,31,3,31,151,31,115,31,235,31,116,31,116,30,154,31,154,30,57,31,14,31,248,31,248,30,14,31,14,30,14,29,14,28,207,31,251,31,222,31,222,30,222,29,50,31,13,31,161,31,198,31,23,31,62,31,58,31,76,31,134,31,134,30,134,29,134,28,134,27,39,31,232,31,157,31,118,31,118,30,233,31,75,31,75,30,237,31,237,30,36,31,21,31,21,30,222,31,122,31,250,31,188,31,165,31,58,31,251,31,218,31,191,31,193,31,2,31,60,31,175,31,254,31,194,31,144,31,15,31,15,30,92,31,85,31,178,31,186,31,186,30,86,31,127,31,8,31,12,31,12,30,12,29,12,28,173,31,27,31,151,31,227,31,80,31,169,31,176,31,176,30,34,31,55,31,151,31,151,30,132,31,124,31,90,31,90,30,176,31,22,31,188,31,67,31,116,31,48,31,72,31,72,30,72,29,218,31,111,31,225,31,232,31,95,31,95,30,95,29,169,31,119,31,76,31,118,31,199,31,136,31,255,31,120,31,120,30,17,31,157,31,42,31,13,31,237,31,142,31,198,31,201,31,122,31,194,31,40,31,40,30,162,31,2,31,133,31,154,31,71,31,225,31,238,31,3,31,112,31,233,31,121,31,33,31,65,31,108,31,131,31,205,31,197,31,220,31,100,31,59,31,92,31,161,31,178,31,74,31,28,31,192,31,55,31,191,31,211,31,111,31,112,31,112,30,78,31,155,31,195,31,195,30,225,31,225,30,104,31,192,31,105,31,12,31,20,31,161,31,35,31,174,31,138,31,159,31,159,30,182,31,182,30,116,31,61,31,17,31,1,31,1,30,138,31,126,31,144,31,172,31,218,31,13,31,107,31,195,31,4,31,4,30,185,31,210,31,210,30,210,29,17,31,92,31,205,31,6,31,249,31,195,31,212,31,135,31,28,31,89,31,116,31,215,31,215,30,125,31,15,31,15,30,15,29,218,31,250,31,197,31,124,31,122,31,33,31,33,30,33,29,137,31,137,30,253,31,116,31,234,31,161,31,109,31,109,30,109,29,109,28,175,31,59,31,59,30,219,31,45,31,45,30,96,31,96,30,10,31,122,31,10,31,118,31,245,31,99,31,246,31,49,31,181,31,204,31,214,31,173,31,173,30,62,31,182,31,135,31,26,31,26,30,225,31,225,30,27,31,27,30,120,31,144,31,144,30,168,31,137,31,9,31,235,31,146,31,205,31,162,31,162,30,239,31,149,31,77,31,33,31,98,31,18,31,18,30,158,31,158,30,158,29,158,28,2,31,35,31,29,31,26,31,54,31,87,31,21,31,254,31,212,31,212,30,212,29,224,31,4,31,153,31,153,30,129,31,241,31,106,31,178,31,97,31,101,31,101,30,101,29,191,31,149,31,80,31,217,31,194,31,145,31,199,31,118,31,75,31,238,31,191,31,191,30,107,31,52,31,7,31,188,31,64,31,64,30,64,29,93,31,121,31,47,31,108,31,108,30,71,31,98,31,168,31,214,31,214,30,214,29,132,31,97,31,97,30,136,31,193,31,130,31,28,31,28,30,118,31,157,31,42,31,118,31,82,31,82,30,167,31,149,31,250,31,127,31,42,31,2,31,2,30,119,31,119,30,78,31,198,31,107,31,113,31,60,31,13,31,13,30,106,31,109,31,56,31,94,31,206,31,231,31,1,31,182,31,221,31,221,30,26,31,219,31,221,31,153,31,31,31,6,31,111,31,239,31,239,30,131,31,77,31,211,31,49,31,137,31,113,31,91,31,214,31,22,31,171,31,171,30,171,29,201,31,94,31,245,31,58,31,249,31,22,31,227,31,215,31,47,31,208,31,208,30,40,31,40,30,40,29,238,31,122,31,86,31,86,30,19,31,51,31,157,31,227,31,227,30,155,31,179,31,133,31,23,31,78,31,78,30,242,31,238,31,254,31,63,31,174,31,81,31,163,31,225,31,46,31,30,31,22,31,209,31,252,31,252,31,252,30,189,31,189,30,233,31,122,31,42,31,148,31,162,31,64,31,64,30,61,31,61,30,191,31,144,31,81,31,234,31,114,31,114,30,242,31,229,31,229,30,247,31,247,30,205,31,31,31,247,31,156,31,136,31,141,31,141,30,225,31,114,31,11,31,144,31,144,30,144,29,17,31,227,31,203,31,145,31,41,31,41,30,193,31,141,31,42,31,114,31,26,31,26,30,26,29,26,28,60,31,182,31,177,31,207,31,182,31,182,30,3,31,104,31,152,31,155,31,94,31,94,30,187,31,47,31,75,31,217,31,40,31,132,31,132,30,132,29,132,28,81,31,124,31,248,31,74,31,74,30,37,31,37,30,10,31,250,31,243,31,231,31,81,31,65,31,65,30,42,31,181,31,150,31,243,31,243,30,179,31,83,31,83,30,237,31,166,31,166,30,54,31,204,31,71,31,219,31,219,30,219,29,219,28,11,31,26,31,162,31,21,31,21,30,21,29,21,28,35,31,21,31,163,31,163,30,211,31,100,31,100,30,231,31,101,31,246,31,246,30,229,31,215,31,127,31,202,31,234,31,216,31,12,31,85,31,1,31,60,31,182,31,98,31,48,31,227,31,218,31,218,30,55,31,1,31,91,31,221,31,219,31,195,31,108,31,172,31,172,30,172,29,172,28,223,31,223,30,25,31,244,31,230,31,230,30,34,31,58,31,26,31,41,31,114,31,114,30,114,29,68,31,68,30,68,29,141,31,164,31,189,31,189,30,40,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
