-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_845 is
end project_tb_845;

architecture project_tb_arch_845 of project_tb_845 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 729;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (20,0,92,0,76,0,27,0,135,0,121,0,118,0,99,0,84,0,0,0,22,0,238,0,40,0,0,0,42,0,58,0,109,0,90,0,17,0,90,0,4,0,255,0,12,0,0,0,202,0,0,0,185,0,189,0,0,0,129,0,157,0,0,0,196,0,210,0,114,0,216,0,199,0,253,0,0,0,54,0,122,0,177,0,175,0,188,0,0,0,77,0,228,0,129,0,14,0,28,0,74,0,60,0,96,0,197,0,0,0,0,0,209,0,85,0,52,0,76,0,151,0,120,0,98,0,180,0,80,0,66,0,15,0,54,0,158,0,98,0,136,0,72,0,224,0,0,0,190,0,0,0,0,0,0,0,0,0,31,0,226,0,58,0,59,0,0,0,251,0,133,0,200,0,0,0,234,0,172,0,91,0,179,0,15,0,164,0,216,0,43,0,254,0,179,0,155,0,31,0,0,0,12,0,36,0,0,0,14,0,250,0,82,0,118,0,198,0,192,0,36,0,229,0,130,0,0,0,82,0,0,0,174,0,165,0,181,0,84,0,19,0,5,0,0,0,0,0,29,0,150,0,237,0,198,0,163,0,0,0,70,0,0,0,36,0,0,0,171,0,99,0,91,0,88,0,183,0,213,0,60,0,239,0,0,0,54,0,4,0,50,0,212,0,90,0,47,0,198,0,138,0,0,0,214,0,187,0,116,0,183,0,24,0,253,0,253,0,182,0,0,0,8,0,82,0,0,0,0,0,0,0,58,0,99,0,115,0,132,0,41,0,80,0,96,0,212,0,12,0,81,0,0,0,145,0,155,0,212,0,244,0,0,0,123,0,0,0,0,0,126,0,209,0,210,0,0,0,8,0,194,0,41,0,50,0,28,0,120,0,237,0,155,0,0,0,107,0,134,0,0,0,0,0,131,0,194,0,204,0,0,0,152,0,174,0,141,0,108,0,148,0,110,0,235,0,207,0,177,0,7,0,0,0,214,0,82,0,45,0,0,0,0,0,240,0,204,0,38,0,29,0,9,0,176,0,228,0,228,0,88,0,178,0,26,0,90,0,0,0,0,0,158,0,34,0,35,0,151,0,30,0,230,0,94,0,44,0,213,0,127,0,181,0,0,0,153,0,195,0,94,0,148,0,74,0,74,0,164,0,12,0,67,0,148,0,249,0,0,0,222,0,153,0,0,0,0,0,33,0,134,0,0,0,36,0,70,0,165,0,134,0,0,0,12,0,175,0,14,0,214,0,0,0,239,0,247,0,179,0,18,0,19,0,134,0,195,0,122,0,49,0,13,0,227,0,160,0,195,0,118,0,200,0,0,0,0,0,120,0,107,0,0,0,0,0,0,0,20,0,212,0,226,0,209,0,84,0,250,0,111,0,5,0,0,0,0,0,0,0,7,0,252,0,0,0,189,0,216,0,172,0,0,0,0,0,139,0,0,0,0,0,215,0,42,0,12,0,37,0,0,0,0,0,254,0,254,0,80,0,185,0,0,0,242,0,0,0,172,0,240,0,12,0,182,0,239,0,212,0,82,0,31,0,104,0,87,0,213,0,167,0,167,0,221,0,216,0,0,0,0,0,11,0,62,0,0,0,223,0,2,0,228,0,185,0,185,0,184,0,25,0,184,0,3,0,255,0,208,0,40,0,152,0,151,0,0,0,30,0,78,0,231,0,82,0,202,0,69,0,132,0,111,0,0,0,50,0,0,0,207,0,245,0,123,0,0,0,150,0,202,0,72,0,0,0,68,0,192,0,125,0,0,0,0,0,63,0,203,0,102,0,61,0,29,0,27,0,13,0,251,0,34,0,139,0,132,0,0,0,19,0,64,0,171,0,0,0,190,0,224,0,82,0,227,0,206,0,130,0,175,0,0,0,48,0,236,0,9,0,23,0,124,0,107,0,0,0,0,0,0,0,0,0,88,0,188,0,177,0,39,0,0,0,192,0,233,0,0,0,0,0,121,0,131,0,16,0,197,0,0,0,0,0,0,0,228,0,236,0,92,0,34,0,255,0,107,0,37,0,0,0,16,0,130,0,24,0,219,0,0,0,0,0,173,0,82,0,0,0,185,0,12,0,0,0,149,0,154,0,252,0,150,0,170,0,0,0,0,0,8,0,0,0,0,0,0,0,15,0,0,0,8,0,55,0,192,0,248,0,150,0,143,0,210,0,0,0,236,0,17,0,85,0,155,0,14,0,86,0,122,0,62,0,171,0,0,0,18,0,24,0,0,0,56,0,252,0,0,0,0,0,136,0,214,0,51,0,162,0,113,0,172,0,0,0,165,0,0,0,185,0,24,0,65,0,238,0,241,0,6,0,0,0,247,0,161,0,109,0,159,0,234,0,34,0,254,0,0,0,244,0,29,0,125,0,213,0,1,0,153,0,36,0,155,0,169,0,237,0,6,0,208,0,60,0,228,0,0,0,0,0,179,0,35,0,0,0,80,0,220,0,82,0,203,0,217,0,158,0,212,0,245,0,0,0,250,0,144,0,207,0,149,0,144,0,193,0,59,0,0,0,219,0,41,0,241,0,158,0,143,0,41,0,0,0,0,0,111,0,91,0,107,0,121,0,214,0,0,0,51,0,104,0,145,0,248,0,180,0,62,0,150,0,122,0,106,0,65,0,0,0,1,0,119,0,0,0,41,0,105,0,0,0,0,0,249,0,237,0,246,0,0,0,0,0,82,0,162,0,11,0,184,0,0,0,163,0,50,0,0,0,198,0,136,0,0,0,0,0,212,0,99,0,55,0,242,0,22,0,150,0,156,0,109,0,104,0,60,0,11,0,123,0,183,0,205,0,8,0,226,0,247,0,0,0,0,0,0,0,6,0,23,0,195,0,11,0,85,0,138,0,231,0,201,0,112,0,126,0,156,0,0,0,239,0,215,0,1,0,226,0,253,0,50,0,0,0,140,0,167,0,0,0,236,0,229,0,0,0,0,0,16,0,163,0,209,0,196,0,226,0,0,0,98,0,7,0,0,0,0,0,81,0,142,0,0,0,0,0,84,0,0,0,55,0,0,0,67,0,41,0,136,0,246,0,211,0,0,0,53,0,14,0,221,0,191,0,59,0,205,0,233,0,0,0,127,0,162,0,124,0,129,0,0,0,168,0,43,0,158,0,0,0,15,0,179,0,206,0,100,0,0,0,0,0,154,0,226,0,3,0,124,0,2,0,171,0,0,0,0,0,19,0,65,0,48,0,132,0,20,0,0,0,214,0,155,0,199,0,197,0,129,0,61,0,8,0,0,0,169,0,192,0,68,0,24,0);
signal scenario_full  : scenario_type := (20,31,92,31,76,31,27,31,135,31,121,31,118,31,99,31,84,31,84,30,22,31,238,31,40,31,40,30,42,31,58,31,109,31,90,31,17,31,90,31,4,31,255,31,12,31,12,30,202,31,202,30,185,31,189,31,189,30,129,31,157,31,157,30,196,31,210,31,114,31,216,31,199,31,253,31,253,30,54,31,122,31,177,31,175,31,188,31,188,30,77,31,228,31,129,31,14,31,28,31,74,31,60,31,96,31,197,31,197,30,197,29,209,31,85,31,52,31,76,31,151,31,120,31,98,31,180,31,80,31,66,31,15,31,54,31,158,31,98,31,136,31,72,31,224,31,224,30,190,31,190,30,190,29,190,28,190,27,31,31,226,31,58,31,59,31,59,30,251,31,133,31,200,31,200,30,234,31,172,31,91,31,179,31,15,31,164,31,216,31,43,31,254,31,179,31,155,31,31,31,31,30,12,31,36,31,36,30,14,31,250,31,82,31,118,31,198,31,192,31,36,31,229,31,130,31,130,30,82,31,82,30,174,31,165,31,181,31,84,31,19,31,5,31,5,30,5,29,29,31,150,31,237,31,198,31,163,31,163,30,70,31,70,30,36,31,36,30,171,31,99,31,91,31,88,31,183,31,213,31,60,31,239,31,239,30,54,31,4,31,50,31,212,31,90,31,47,31,198,31,138,31,138,30,214,31,187,31,116,31,183,31,24,31,253,31,253,31,182,31,182,30,8,31,82,31,82,30,82,29,82,28,58,31,99,31,115,31,132,31,41,31,80,31,96,31,212,31,12,31,81,31,81,30,145,31,155,31,212,31,244,31,244,30,123,31,123,30,123,29,126,31,209,31,210,31,210,30,8,31,194,31,41,31,50,31,28,31,120,31,237,31,155,31,155,30,107,31,134,31,134,30,134,29,131,31,194,31,204,31,204,30,152,31,174,31,141,31,108,31,148,31,110,31,235,31,207,31,177,31,7,31,7,30,214,31,82,31,45,31,45,30,45,29,240,31,204,31,38,31,29,31,9,31,176,31,228,31,228,31,88,31,178,31,26,31,90,31,90,30,90,29,158,31,34,31,35,31,151,31,30,31,230,31,94,31,44,31,213,31,127,31,181,31,181,30,153,31,195,31,94,31,148,31,74,31,74,31,164,31,12,31,67,31,148,31,249,31,249,30,222,31,153,31,153,30,153,29,33,31,134,31,134,30,36,31,70,31,165,31,134,31,134,30,12,31,175,31,14,31,214,31,214,30,239,31,247,31,179,31,18,31,19,31,134,31,195,31,122,31,49,31,13,31,227,31,160,31,195,31,118,31,200,31,200,30,200,29,120,31,107,31,107,30,107,29,107,28,20,31,212,31,226,31,209,31,84,31,250,31,111,31,5,31,5,30,5,29,5,28,7,31,252,31,252,30,189,31,216,31,172,31,172,30,172,29,139,31,139,30,139,29,215,31,42,31,12,31,37,31,37,30,37,29,254,31,254,31,80,31,185,31,185,30,242,31,242,30,172,31,240,31,12,31,182,31,239,31,212,31,82,31,31,31,104,31,87,31,213,31,167,31,167,31,221,31,216,31,216,30,216,29,11,31,62,31,62,30,223,31,2,31,228,31,185,31,185,31,184,31,25,31,184,31,3,31,255,31,208,31,40,31,152,31,151,31,151,30,30,31,78,31,231,31,82,31,202,31,69,31,132,31,111,31,111,30,50,31,50,30,207,31,245,31,123,31,123,30,150,31,202,31,72,31,72,30,68,31,192,31,125,31,125,30,125,29,63,31,203,31,102,31,61,31,29,31,27,31,13,31,251,31,34,31,139,31,132,31,132,30,19,31,64,31,171,31,171,30,190,31,224,31,82,31,227,31,206,31,130,31,175,31,175,30,48,31,236,31,9,31,23,31,124,31,107,31,107,30,107,29,107,28,107,27,88,31,188,31,177,31,39,31,39,30,192,31,233,31,233,30,233,29,121,31,131,31,16,31,197,31,197,30,197,29,197,28,228,31,236,31,92,31,34,31,255,31,107,31,37,31,37,30,16,31,130,31,24,31,219,31,219,30,219,29,173,31,82,31,82,30,185,31,12,31,12,30,149,31,154,31,252,31,150,31,170,31,170,30,170,29,8,31,8,30,8,29,8,28,15,31,15,30,8,31,55,31,192,31,248,31,150,31,143,31,210,31,210,30,236,31,17,31,85,31,155,31,14,31,86,31,122,31,62,31,171,31,171,30,18,31,24,31,24,30,56,31,252,31,252,30,252,29,136,31,214,31,51,31,162,31,113,31,172,31,172,30,165,31,165,30,185,31,24,31,65,31,238,31,241,31,6,31,6,30,247,31,161,31,109,31,159,31,234,31,34,31,254,31,254,30,244,31,29,31,125,31,213,31,1,31,153,31,36,31,155,31,169,31,237,31,6,31,208,31,60,31,228,31,228,30,228,29,179,31,35,31,35,30,80,31,220,31,82,31,203,31,217,31,158,31,212,31,245,31,245,30,250,31,144,31,207,31,149,31,144,31,193,31,59,31,59,30,219,31,41,31,241,31,158,31,143,31,41,31,41,30,41,29,111,31,91,31,107,31,121,31,214,31,214,30,51,31,104,31,145,31,248,31,180,31,62,31,150,31,122,31,106,31,65,31,65,30,1,31,119,31,119,30,41,31,105,31,105,30,105,29,249,31,237,31,246,31,246,30,246,29,82,31,162,31,11,31,184,31,184,30,163,31,50,31,50,30,198,31,136,31,136,30,136,29,212,31,99,31,55,31,242,31,22,31,150,31,156,31,109,31,104,31,60,31,11,31,123,31,183,31,205,31,8,31,226,31,247,31,247,30,247,29,247,28,6,31,23,31,195,31,11,31,85,31,138,31,231,31,201,31,112,31,126,31,156,31,156,30,239,31,215,31,1,31,226,31,253,31,50,31,50,30,140,31,167,31,167,30,236,31,229,31,229,30,229,29,16,31,163,31,209,31,196,31,226,31,226,30,98,31,7,31,7,30,7,29,81,31,142,31,142,30,142,29,84,31,84,30,55,31,55,30,67,31,41,31,136,31,246,31,211,31,211,30,53,31,14,31,221,31,191,31,59,31,205,31,233,31,233,30,127,31,162,31,124,31,129,31,129,30,168,31,43,31,158,31,158,30,15,31,179,31,206,31,100,31,100,30,100,29,154,31,226,31,3,31,124,31,2,31,171,31,171,30,171,29,19,31,65,31,48,31,132,31,20,31,20,30,214,31,155,31,199,31,197,31,129,31,61,31,8,31,8,30,169,31,192,31,68,31,24,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
