-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 807;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (184,0,142,0,224,0,193,0,0,0,91,0,179,0,149,0,70,0,247,0,14,0,0,0,67,0,176,0,0,0,0,0,0,0,0,0,247,0,254,0,88,0,136,0,0,0,6,0,211,0,0,0,0,0,0,0,238,0,56,0,65,0,22,0,31,0,0,0,159,0,74,0,201,0,53,0,214,0,0,0,183,0,98,0,110,0,122,0,130,0,218,0,37,0,0,0,133,0,124,0,223,0,0,0,238,0,184,0,76,0,208,0,0,0,0,0,190,0,165,0,255,0,161,0,82,0,36,0,0,0,57,0,194,0,154,0,238,0,64,0,189,0,115,0,68,0,168,0,0,0,241,0,90,0,0,0,0,0,196,0,6,0,211,0,164,0,99,0,223,0,12,0,92,0,198,0,241,0,112,0,93,0,114,0,30,0,108,0,177,0,0,0,0,0,140,0,0,0,155,0,0,0,171,0,71,0,0,0,211,0,249,0,236,0,178,0,216,0,213,0,171,0,174,0,63,0,0,0,0,0,70,0,158,0,46,0,225,0,102,0,0,0,12,0,0,0,0,0,206,0,12,0,46,0,181,0,76,0,82,0,210,0,227,0,95,0,0,0,88,0,0,0,147,0,7,0,100,0,21,0,12,0,17,0,0,0,0,0,189,0,0,0,201,0,0,0,0,0,151,0,169,0,84,0,160,0,151,0,157,0,72,0,0,0,9,0,255,0,6,0,0,0,12,0,0,0,90,0,0,0,138,0,112,0,204,0,236,0,229,0,0,0,149,0,0,0,30,0,103,0,159,0,0,0,20,0,230,0,40,0,0,0,62,0,169,0,164,0,0,0,86,0,79,0,0,0,251,0,0,0,41,0,154,0,20,0,97,0,197,0,10,0,87,0,0,0,108,0,0,0,81,0,237,0,0,0,169,0,58,0,173,0,214,0,242,0,185,0,128,0,86,0,113,0,92,0,225,0,0,0,12,0,15,0,0,0,240,0,0,0,9,0,0,0,40,0,45,0,0,0,36,0,227,0,126,0,38,0,7,0,179,0,100,0,95,0,161,0,233,0,249,0,138,0,16,0,235,0,254,0,160,0,0,0,0,0,24,0,237,0,0,0,142,0,75,0,115,0,0,0,234,0,143,0,3,0,0,0,137,0,0,0,220,0,54,0,0,0,171,0,246,0,14,0,42,0,0,0,129,0,222,0,0,0,152,0,0,0,51,0,237,0,128,0,254,0,178,0,34,0,2,0,160,0,29,0,16,0,242,0,15,0,7,0,151,0,43,0,91,0,201,0,150,0,226,0,156,0,223,0,97,0,10,0,215,0,66,0,64,0,97,0,251,0,132,0,37,0,243,0,95,0,179,0,0,0,0,0,145,0,71,0,0,0,237,0,51,0,0,0,110,0,108,0,13,0,172,0,150,0,47,0,244,0,205,0,23,0,94,0,192,0,0,0,49,0,40,0,135,0,67,0,2,0,234,0,16,0,0,0,42,0,116,0,43,0,239,0,160,0,95,0,160,0,241,0,50,0,203,0,106,0,254,0,200,0,0,0,142,0,55,0,190,0,7,0,92,0,187,0,0,0,60,0,102,0,66,0,0,0,77,0,225,0,189,0,0,0,245,0,66,0,0,0,0,0,146,0,61,0,255,0,110,0,51,0,45,0,230,0,207,0,0,0,0,0,72,0,0,0,0,0,104,0,178,0,0,0,204,0,116,0,35,0,41,0,13,0,49,0,18,0,0,0,105,0,150,0,192,0,117,0,150,0,170,0,133,0,224,0,44,0,0,0,76,0,225,0,206,0,0,0,0,0,0,0,25,0,0,0,9,0,0,0,35,0,17,0,167,0,0,0,88,0,24,0,17,0,28,0,202,0,198,0,219,0,157,0,0,0,128,0,0,0,0,0,233,0,82,0,40,0,130,0,43,0,224,0,80,0,204,0,49,0,0,0,96,0,131,0,251,0,111,0,172,0,253,0,63,0,227,0,55,0,93,0,17,0,90,0,38,0,82,0,203,0,113,0,46,0,0,0,239,0,129,0,198,0,223,0,169,0,106,0,20,0,47,0,0,0,174,0,0,0,17,0,60,0,238,0,182,0,0,0,24,0,0,0,69,0,72,0,0,0,50,0,246,0,0,0,14,0,0,0,175,0,0,0,211,0,0,0,244,0,57,0,236,0,253,0,73,0,0,0,166,0,196,0,201,0,190,0,150,0,27,0,220,0,35,0,235,0,150,0,0,0,0,0,213,0,3,0,27,0,0,0,0,0,53,0,196,0,209,0,195,0,134,0,6,0,251,0,225,0,134,0,150,0,86,0,235,0,80,0,0,0,39,0,87,0,250,0,201,0,0,0,168,0,117,0,133,0,52,0,0,0,179,0,124,0,92,0,200,0,5,0,216,0,47,0,0,0,141,0,180,0,45,0,0,0,0,0,35,0,69,0,0,0,0,0,236,0,103,0,0,0,0,0,0,0,232,0,222,0,214,0,0,0,53,0,11,0,252,0,184,0,246,0,0,0,146,0,233,0,0,0,184,0,41,0,218,0,205,0,0,0,13,0,0,0,52,0,41,0,0,0,0,0,95,0,29,0,0,0,247,0,122,0,180,0,178,0,135,0,8,0,0,0,100,0,220,0,0,0,177,0,133,0,0,0,3,0,45,0,143,0,18,0,199,0,48,0,62,0,184,0,240,0,53,0,255,0,125,0,90,0,80,0,7,0,166,0,19,0,8,0,252,0,149,0,30,0,173,0,211,0,0,0,252,0,25,0,0,0,214,0,0,0,249,0,0,0,0,0,0,0,188,0,73,0,41,0,178,0,185,0,74,0,0,0,0,0,195,0,207,0,179,0,138,0,207,0,49,0,23,0,35,0,157,0,185,0,30,0,172,0,127,0,106,0,0,0,222,0,47,0,98,0,27,0,240,0,164,0,203,0,0,0,240,0,166,0,203,0,128,0,81,0,102,0,0,0,51,0,3,0,254,0,165,0,216,0,63,0,62,0,134,0,116,0,108,0,192,0,116,0,95,0,212,0,34,0,0,0,19,0,184,0,79,0,120,0,55,0,15,0,255,0,41,0,20,0,0,0,138,0,165,0,191,0,115,0,53,0,227,0,0,0,184,0,199,0,19,0,129,0,255,0,15,0,22,0,0,0,225,0,0,0,0,0,148,0,0,0,0,0,229,0,165,0,42,0,48,0,1,0,177,0,0,0,145,0,206,0,237,0,1,0,0,0,156,0,27,0,77,0,55,0,94,0,10,0,206,0,25,0,137,0,0,0,0,0,200,0,163,0,55,0,230,0,202,0,121,0,21,0,95,0,240,0,126,0,102,0,229,0,80,0,86,0,0,0,2,0,173,0,196,0,225,0,0,0,0,0,0,0,104,0,0,0,34,0,99,0,0,0,232,0,128,0,180,0,102,0,0,0,11,0,0,0,206,0,182,0,193,0,35,0,26,0,144,0,76,0,79,0,60,0,0,0,0,0,76,0,158,0,149,0,180,0,101,0,104,0,79,0,0,0,142,0,106,0,172,0,25,0,84,0,93,0,12,0,253,0,150,0,0,0,254,0,31,0,3,0,140,0,34,0,50,0,78,0,67,0,169,0,245,0,0,0,131,0,0,0);
signal scenario_full  : scenario_type := (184,31,142,31,224,31,193,31,193,30,91,31,179,31,149,31,70,31,247,31,14,31,14,30,67,31,176,31,176,30,176,29,176,28,176,27,247,31,254,31,88,31,136,31,136,30,6,31,211,31,211,30,211,29,211,28,238,31,56,31,65,31,22,31,31,31,31,30,159,31,74,31,201,31,53,31,214,31,214,30,183,31,98,31,110,31,122,31,130,31,218,31,37,31,37,30,133,31,124,31,223,31,223,30,238,31,184,31,76,31,208,31,208,30,208,29,190,31,165,31,255,31,161,31,82,31,36,31,36,30,57,31,194,31,154,31,238,31,64,31,189,31,115,31,68,31,168,31,168,30,241,31,90,31,90,30,90,29,196,31,6,31,211,31,164,31,99,31,223,31,12,31,92,31,198,31,241,31,112,31,93,31,114,31,30,31,108,31,177,31,177,30,177,29,140,31,140,30,155,31,155,30,171,31,71,31,71,30,211,31,249,31,236,31,178,31,216,31,213,31,171,31,174,31,63,31,63,30,63,29,70,31,158,31,46,31,225,31,102,31,102,30,12,31,12,30,12,29,206,31,12,31,46,31,181,31,76,31,82,31,210,31,227,31,95,31,95,30,88,31,88,30,147,31,7,31,100,31,21,31,12,31,17,31,17,30,17,29,189,31,189,30,201,31,201,30,201,29,151,31,169,31,84,31,160,31,151,31,157,31,72,31,72,30,9,31,255,31,6,31,6,30,12,31,12,30,90,31,90,30,138,31,112,31,204,31,236,31,229,31,229,30,149,31,149,30,30,31,103,31,159,31,159,30,20,31,230,31,40,31,40,30,62,31,169,31,164,31,164,30,86,31,79,31,79,30,251,31,251,30,41,31,154,31,20,31,97,31,197,31,10,31,87,31,87,30,108,31,108,30,81,31,237,31,237,30,169,31,58,31,173,31,214,31,242,31,185,31,128,31,86,31,113,31,92,31,225,31,225,30,12,31,15,31,15,30,240,31,240,30,9,31,9,30,40,31,45,31,45,30,36,31,227,31,126,31,38,31,7,31,179,31,100,31,95,31,161,31,233,31,249,31,138,31,16,31,235,31,254,31,160,31,160,30,160,29,24,31,237,31,237,30,142,31,75,31,115,31,115,30,234,31,143,31,3,31,3,30,137,31,137,30,220,31,54,31,54,30,171,31,246,31,14,31,42,31,42,30,129,31,222,31,222,30,152,31,152,30,51,31,237,31,128,31,254,31,178,31,34,31,2,31,160,31,29,31,16,31,242,31,15,31,7,31,151,31,43,31,91,31,201,31,150,31,226,31,156,31,223,31,97,31,10,31,215,31,66,31,64,31,97,31,251,31,132,31,37,31,243,31,95,31,179,31,179,30,179,29,145,31,71,31,71,30,237,31,51,31,51,30,110,31,108,31,13,31,172,31,150,31,47,31,244,31,205,31,23,31,94,31,192,31,192,30,49,31,40,31,135,31,67,31,2,31,234,31,16,31,16,30,42,31,116,31,43,31,239,31,160,31,95,31,160,31,241,31,50,31,203,31,106,31,254,31,200,31,200,30,142,31,55,31,190,31,7,31,92,31,187,31,187,30,60,31,102,31,66,31,66,30,77,31,225,31,189,31,189,30,245,31,66,31,66,30,66,29,146,31,61,31,255,31,110,31,51,31,45,31,230,31,207,31,207,30,207,29,72,31,72,30,72,29,104,31,178,31,178,30,204,31,116,31,35,31,41,31,13,31,49,31,18,31,18,30,105,31,150,31,192,31,117,31,150,31,170,31,133,31,224,31,44,31,44,30,76,31,225,31,206,31,206,30,206,29,206,28,25,31,25,30,9,31,9,30,35,31,17,31,167,31,167,30,88,31,24,31,17,31,28,31,202,31,198,31,219,31,157,31,157,30,128,31,128,30,128,29,233,31,82,31,40,31,130,31,43,31,224,31,80,31,204,31,49,31,49,30,96,31,131,31,251,31,111,31,172,31,253,31,63,31,227,31,55,31,93,31,17,31,90,31,38,31,82,31,203,31,113,31,46,31,46,30,239,31,129,31,198,31,223,31,169,31,106,31,20,31,47,31,47,30,174,31,174,30,17,31,60,31,238,31,182,31,182,30,24,31,24,30,69,31,72,31,72,30,50,31,246,31,246,30,14,31,14,30,175,31,175,30,211,31,211,30,244,31,57,31,236,31,253,31,73,31,73,30,166,31,196,31,201,31,190,31,150,31,27,31,220,31,35,31,235,31,150,31,150,30,150,29,213,31,3,31,27,31,27,30,27,29,53,31,196,31,209,31,195,31,134,31,6,31,251,31,225,31,134,31,150,31,86,31,235,31,80,31,80,30,39,31,87,31,250,31,201,31,201,30,168,31,117,31,133,31,52,31,52,30,179,31,124,31,92,31,200,31,5,31,216,31,47,31,47,30,141,31,180,31,45,31,45,30,45,29,35,31,69,31,69,30,69,29,236,31,103,31,103,30,103,29,103,28,232,31,222,31,214,31,214,30,53,31,11,31,252,31,184,31,246,31,246,30,146,31,233,31,233,30,184,31,41,31,218,31,205,31,205,30,13,31,13,30,52,31,41,31,41,30,41,29,95,31,29,31,29,30,247,31,122,31,180,31,178,31,135,31,8,31,8,30,100,31,220,31,220,30,177,31,133,31,133,30,3,31,45,31,143,31,18,31,199,31,48,31,62,31,184,31,240,31,53,31,255,31,125,31,90,31,80,31,7,31,166,31,19,31,8,31,252,31,149,31,30,31,173,31,211,31,211,30,252,31,25,31,25,30,214,31,214,30,249,31,249,30,249,29,249,28,188,31,73,31,41,31,178,31,185,31,74,31,74,30,74,29,195,31,207,31,179,31,138,31,207,31,49,31,23,31,35,31,157,31,185,31,30,31,172,31,127,31,106,31,106,30,222,31,47,31,98,31,27,31,240,31,164,31,203,31,203,30,240,31,166,31,203,31,128,31,81,31,102,31,102,30,51,31,3,31,254,31,165,31,216,31,63,31,62,31,134,31,116,31,108,31,192,31,116,31,95,31,212,31,34,31,34,30,19,31,184,31,79,31,120,31,55,31,15,31,255,31,41,31,20,31,20,30,138,31,165,31,191,31,115,31,53,31,227,31,227,30,184,31,199,31,19,31,129,31,255,31,15,31,22,31,22,30,225,31,225,30,225,29,148,31,148,30,148,29,229,31,165,31,42,31,48,31,1,31,177,31,177,30,145,31,206,31,237,31,1,31,1,30,156,31,27,31,77,31,55,31,94,31,10,31,206,31,25,31,137,31,137,30,137,29,200,31,163,31,55,31,230,31,202,31,121,31,21,31,95,31,240,31,126,31,102,31,229,31,80,31,86,31,86,30,2,31,173,31,196,31,225,31,225,30,225,29,225,28,104,31,104,30,34,31,99,31,99,30,232,31,128,31,180,31,102,31,102,30,11,31,11,30,206,31,182,31,193,31,35,31,26,31,144,31,76,31,79,31,60,31,60,30,60,29,76,31,158,31,149,31,180,31,101,31,104,31,79,31,79,30,142,31,106,31,172,31,25,31,84,31,93,31,12,31,253,31,150,31,150,30,254,31,31,31,3,31,140,31,34,31,50,31,78,31,67,31,169,31,245,31,245,30,131,31,131,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
