-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 993;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (236,0,0,0,111,0,67,0,166,0,165,0,243,0,182,0,111,0,188,0,242,0,209,0,21,0,180,0,234,0,158,0,59,0,0,0,95,0,137,0,0,0,150,0,0,0,128,0,0,0,0,0,155,0,189,0,0,0,182,0,139,0,154,0,249,0,196,0,0,0,76,0,0,0,67,0,68,0,0,0,41,0,59,0,0,0,155,0,208,0,234,0,125,0,0,0,238,0,119,0,107,0,238,0,236,0,8,0,207,0,0,0,106,0,106,0,0,0,75,0,158,0,49,0,220,0,97,0,25,0,176,0,15,0,246,0,0,0,130,0,141,0,89,0,87,0,128,0,243,0,126,0,161,0,0,0,94,0,0,0,0,0,0,0,15,0,0,0,103,0,0,0,71,0,127,0,75,0,0,0,169,0,78,0,127,0,131,0,249,0,227,0,103,0,42,0,10,0,61,0,44,0,134,0,141,0,146,0,72,0,168,0,22,0,230,0,144,0,123,0,107,0,142,0,160,0,235,0,40,0,0,0,162,0,241,0,107,0,180,0,150,0,150,0,0,0,74,0,119,0,153,0,112,0,13,0,16,0,0,0,229,0,37,0,141,0,168,0,1,0,114,0,14,0,27,0,0,0,230,0,53,0,190,0,172,0,61,0,167,0,14,0,44,0,226,0,76,0,198,0,0,0,19,0,0,0,152,0,33,0,129,0,180,0,151,0,26,0,10,0,167,0,141,0,113,0,0,0,111,0,209,0,113,0,249,0,0,0,160,0,149,0,240,0,98,0,184,0,185,0,0,0,3,0,0,0,131,0,185,0,0,0,44,0,0,0,93,0,0,0,94,0,0,0,215,0,85,0,0,0,153,0,249,0,218,0,193,0,0,0,10,0,191,0,229,0,135,0,237,0,15,0,116,0,0,0,129,0,0,0,120,0,165,0,180,0,244,0,255,0,178,0,0,0,140,0,239,0,86,0,13,0,85,0,186,0,0,0,211,0,107,0,135,0,0,0,185,0,153,0,32,0,0,0,206,0,227,0,36,0,23,0,0,0,0,0,205,0,0,0,117,0,224,0,169,0,0,0,0,0,111,0,198,0,174,0,250,0,135,0,210,0,135,0,216,0,142,0,212,0,236,0,0,0,0,0,94,0,12,0,145,0,46,0,144,0,28,0,255,0,56,0,179,0,0,0,0,0,252,0,127,0,0,0,130,0,44,0,70,0,138,0,0,0,0,0,0,0,193,0,67,0,163,0,0,0,223,0,57,0,104,0,187,0,200,0,0,0,193,0,153,0,237,0,18,0,194,0,59,0,106,0,160,0,218,0,13,0,208,0,0,0,0,0,2,0,127,0,152,0,0,0,77,0,116,0,152,0,212,0,0,0,43,0,56,0,243,0,25,0,83,0,204,0,15,0,53,0,120,0,0,0,139,0,126,0,0,0,246,0,149,0,12,0,119,0,135,0,84,0,241,0,23,0,144,0,72,0,250,0,80,0,191,0,45,0,240,0,225,0,238,0,0,0,69,0,0,0,121,0,245,0,0,0,249,0,0,0,25,0,248,0,81,0,182,0,91,0,175,0,147,0,0,0,226,0,144,0,234,0,74,0,0,0,0,0,134,0,44,0,0,0,0,0,54,0,34,0,190,0,186,0,121,0,175,0,112,0,115,0,134,0,77,0,175,0,210,0,0,0,0,0,34,0,75,0,204,0,46,0,128,0,0,0,0,0,35,0,77,0,197,0,20,0,0,0,76,0,0,0,216,0,0,0,200,0,29,0,240,0,0,0,7,0,174,0,0,0,125,0,253,0,134,0,201,0,80,0,107,0,0,0,143,0,182,0,48,0,0,0,111,0,87,0,37,0,89,0,243,0,110,0,196,0,165,0,38,0,0,0,211,0,67,0,8,0,76,0,0,0,210,0,4,0,162,0,217,0,0,0,29,0,146,0,33,0,223,0,0,0,120,0,154,0,162,0,74,0,128,0,0,0,0,0,202,0,235,0,60,0,44,0,0,0,0,0,227,0,36,0,237,0,128,0,181,0,234,0,0,0,199,0,38,0,229,0,138,0,8,0,0,0,138,0,61,0,117,0,126,0,243,0,0,0,97,0,143,0,45,0,248,0,165,0,233,0,74,0,163,0,230,0,201,0,185,0,232,0,0,0,38,0,86,0,201,0,11,0,0,0,108,0,34,0,70,0,216,0,245,0,9,0,199,0,129,0,139,0,14,0,48,0,0,0,165,0,159,0,0,0,0,0,156,0,146,0,66,0,188,0,214,0,0,0,53,0,108,0,108,0,118,0,0,0,85,0,116,0,153,0,133,0,36,0,134,0,197,0,70,0,88,0,222,0,217,0,0,0,237,0,124,0,210,0,0,0,248,0,201,0,144,0,233,0,164,0,39,0,234,0,0,0,161,0,90,0,190,0,0,0,172,0,109,0,119,0,40,0,1,0,52,0,175,0,0,0,192,0,0,0,62,0,0,0,227,0,167,0,236,0,29,0,66,0,0,0,59,0,219,0,73,0,205,0,220,0,245,0,92,0,134,0,132,0,171,0,112,0,162,0,82,0,175,0,0,0,23,0,0,0,182,0,106,0,32,0,3,0,0,0,142,0,233,0,0,0,92,0,171,0,77,0,3,0,113,0,189,0,56,0,100,0,11,0,236,0,36,0,0,0,247,0,77,0,223,0,131,0,162,0,0,0,24,0,201,0,11,0,119,0,144,0,68,0,57,0,0,0,233,0,136,0,247,0,96,0,17,0,211,0,37,0,187,0,0,0,14,0,0,0,66,0,0,0,119,0,0,0,0,0,74,0,32,0,0,0,0,0,199,0,10,0,220,0,5,0,179,0,178,0,115,0,149,0,0,0,127,0,94,0,0,0,83,0,0,0,149,0,0,0,32,0,120,0,0,0,135,0,136,0,126,0,17,0,0,0,0,0,3,0,0,0,82,0,63,0,0,0,0,0,84,0,71,0,141,0,182,0,116,0,91,0,0,0,22,0,13,0,96,0,83,0,127,0,163,0,7,0,215,0,142,0,160,0,109,0,0,0,177,0,40,0,48,0,0,0,238,0,86,0,0,0,0,0,227,0,0,0,0,0,0,0,130,0,18,0,31,0,147,0,0,0,87,0,90,0,253,0,182,0,39,0,18,0,32,0,75,0,238,0,157,0,0,0,232,0,232,0,112,0,0,0,0,0,81,0,254,0,9,0,39,0,194,0,0,0,0,0,165,0,176,0,41,0,0,0,49,0,160,0,0,0,64,0,147,0,52,0,52,0,234,0,109,0,0,0,19,0,209,0,208,0,58,0,183,0,0,0,229,0,234,0,22,0,187,0,217,0,0,0,41,0,213,0,209,0,127,0,5,0,214,0,0,0,114,0,0,0,52,0,28,0,5,0,175,0,178,0,134,0,42,0,29,0,0,0,71,0,202,0,177,0,105,0,172,0,148,0,31,0,193,0,70,0,130,0,75,0,194,0,39,0,135,0,0,0,214,0,235,0,0,0,136,0,141,0,0,0,99,0,0,0,171,0,31,0,114,0,52,0,29,0,1,0,73,0,212,0,0,0,127,0,99,0,133,0,0,0,126,0,111,0,137,0,222,0,0,0,33,0,216,0,17,0,0,0,167,0,169,0,152,0,114,0,234,0,0,0,249,0,205,0,222,0,83,0,16,0,70,0,144,0,159,0,60,0,20,0,84,0,218,0,0,0,0,0,0,0,0,0,202,0,202,0,0,0,224,0,107,0,226,0,248,0,224,0,0,0,83,0,10,0,62,0,248,0,39,0,172,0,0,0,215,0,196,0,11,0,15,0,0,0,79,0,13,0,186,0,0,0,228,0,0,0,0,0,246,0,160,0,209,0,217,0,147,0,88,0,252,0,250,0,0,0,0,0,58,0,242,0,206,0,93,0,0,0,79,0,94,0,186,0,111,0,44,0,128,0,180,0,16,0,180,0,158,0,0,0,65,0,108,0,206,0,0,0,226,0,0,0,184,0,0,0,32,0,148,0,136,0,193,0,140,0,208,0,0,0,29,0,0,0,0,0,40,0,25,0,118,0,166,0,180,0,209,0,181,0,30,0,178,0,61,0,56,0,228,0,201,0,5,0,194,0,0,0,195,0,0,0,159,0,207,0,227,0,206,0,139,0,101,0,103,0,0,0,32,0,10,0,29,0,134,0,134,0,183,0,94,0,202,0,149,0,15,0,213,0,178,0,244,0,0,0,0,0,0,0,35,0,0,0,206,0,60,0,165,0,214,0,148,0,0,0,0,0,88,0,15,0,195,0,146,0,0,0,0,0,125,0,11,0,240,0,84,0,248,0,128,0,8,0,94,0,0,0,47,0,0,0,54,0,203,0,0,0,216,0,120,0,244,0,111,0,74,0,46,0,103,0,25,0,214,0,217,0,118,0,224,0,228,0,186,0,142,0,123,0,35,0,102,0,101,0,137,0);
signal scenario_full  : scenario_type := (236,31,236,30,111,31,67,31,166,31,165,31,243,31,182,31,111,31,188,31,242,31,209,31,21,31,180,31,234,31,158,31,59,31,59,30,95,31,137,31,137,30,150,31,150,30,128,31,128,30,128,29,155,31,189,31,189,30,182,31,139,31,154,31,249,31,196,31,196,30,76,31,76,30,67,31,68,31,68,30,41,31,59,31,59,30,155,31,208,31,234,31,125,31,125,30,238,31,119,31,107,31,238,31,236,31,8,31,207,31,207,30,106,31,106,31,106,30,75,31,158,31,49,31,220,31,97,31,25,31,176,31,15,31,246,31,246,30,130,31,141,31,89,31,87,31,128,31,243,31,126,31,161,31,161,30,94,31,94,30,94,29,94,28,15,31,15,30,103,31,103,30,71,31,127,31,75,31,75,30,169,31,78,31,127,31,131,31,249,31,227,31,103,31,42,31,10,31,61,31,44,31,134,31,141,31,146,31,72,31,168,31,22,31,230,31,144,31,123,31,107,31,142,31,160,31,235,31,40,31,40,30,162,31,241,31,107,31,180,31,150,31,150,31,150,30,74,31,119,31,153,31,112,31,13,31,16,31,16,30,229,31,37,31,141,31,168,31,1,31,114,31,14,31,27,31,27,30,230,31,53,31,190,31,172,31,61,31,167,31,14,31,44,31,226,31,76,31,198,31,198,30,19,31,19,30,152,31,33,31,129,31,180,31,151,31,26,31,10,31,167,31,141,31,113,31,113,30,111,31,209,31,113,31,249,31,249,30,160,31,149,31,240,31,98,31,184,31,185,31,185,30,3,31,3,30,131,31,185,31,185,30,44,31,44,30,93,31,93,30,94,31,94,30,215,31,85,31,85,30,153,31,249,31,218,31,193,31,193,30,10,31,191,31,229,31,135,31,237,31,15,31,116,31,116,30,129,31,129,30,120,31,165,31,180,31,244,31,255,31,178,31,178,30,140,31,239,31,86,31,13,31,85,31,186,31,186,30,211,31,107,31,135,31,135,30,185,31,153,31,32,31,32,30,206,31,227,31,36,31,23,31,23,30,23,29,205,31,205,30,117,31,224,31,169,31,169,30,169,29,111,31,198,31,174,31,250,31,135,31,210,31,135,31,216,31,142,31,212,31,236,31,236,30,236,29,94,31,12,31,145,31,46,31,144,31,28,31,255,31,56,31,179,31,179,30,179,29,252,31,127,31,127,30,130,31,44,31,70,31,138,31,138,30,138,29,138,28,193,31,67,31,163,31,163,30,223,31,57,31,104,31,187,31,200,31,200,30,193,31,153,31,237,31,18,31,194,31,59,31,106,31,160,31,218,31,13,31,208,31,208,30,208,29,2,31,127,31,152,31,152,30,77,31,116,31,152,31,212,31,212,30,43,31,56,31,243,31,25,31,83,31,204,31,15,31,53,31,120,31,120,30,139,31,126,31,126,30,246,31,149,31,12,31,119,31,135,31,84,31,241,31,23,31,144,31,72,31,250,31,80,31,191,31,45,31,240,31,225,31,238,31,238,30,69,31,69,30,121,31,245,31,245,30,249,31,249,30,25,31,248,31,81,31,182,31,91,31,175,31,147,31,147,30,226,31,144,31,234,31,74,31,74,30,74,29,134,31,44,31,44,30,44,29,54,31,34,31,190,31,186,31,121,31,175,31,112,31,115,31,134,31,77,31,175,31,210,31,210,30,210,29,34,31,75,31,204,31,46,31,128,31,128,30,128,29,35,31,77,31,197,31,20,31,20,30,76,31,76,30,216,31,216,30,200,31,29,31,240,31,240,30,7,31,174,31,174,30,125,31,253,31,134,31,201,31,80,31,107,31,107,30,143,31,182,31,48,31,48,30,111,31,87,31,37,31,89,31,243,31,110,31,196,31,165,31,38,31,38,30,211,31,67,31,8,31,76,31,76,30,210,31,4,31,162,31,217,31,217,30,29,31,146,31,33,31,223,31,223,30,120,31,154,31,162,31,74,31,128,31,128,30,128,29,202,31,235,31,60,31,44,31,44,30,44,29,227,31,36,31,237,31,128,31,181,31,234,31,234,30,199,31,38,31,229,31,138,31,8,31,8,30,138,31,61,31,117,31,126,31,243,31,243,30,97,31,143,31,45,31,248,31,165,31,233,31,74,31,163,31,230,31,201,31,185,31,232,31,232,30,38,31,86,31,201,31,11,31,11,30,108,31,34,31,70,31,216,31,245,31,9,31,199,31,129,31,139,31,14,31,48,31,48,30,165,31,159,31,159,30,159,29,156,31,146,31,66,31,188,31,214,31,214,30,53,31,108,31,108,31,118,31,118,30,85,31,116,31,153,31,133,31,36,31,134,31,197,31,70,31,88,31,222,31,217,31,217,30,237,31,124,31,210,31,210,30,248,31,201,31,144,31,233,31,164,31,39,31,234,31,234,30,161,31,90,31,190,31,190,30,172,31,109,31,119,31,40,31,1,31,52,31,175,31,175,30,192,31,192,30,62,31,62,30,227,31,167,31,236,31,29,31,66,31,66,30,59,31,219,31,73,31,205,31,220,31,245,31,92,31,134,31,132,31,171,31,112,31,162,31,82,31,175,31,175,30,23,31,23,30,182,31,106,31,32,31,3,31,3,30,142,31,233,31,233,30,92,31,171,31,77,31,3,31,113,31,189,31,56,31,100,31,11,31,236,31,36,31,36,30,247,31,77,31,223,31,131,31,162,31,162,30,24,31,201,31,11,31,119,31,144,31,68,31,57,31,57,30,233,31,136,31,247,31,96,31,17,31,211,31,37,31,187,31,187,30,14,31,14,30,66,31,66,30,119,31,119,30,119,29,74,31,32,31,32,30,32,29,199,31,10,31,220,31,5,31,179,31,178,31,115,31,149,31,149,30,127,31,94,31,94,30,83,31,83,30,149,31,149,30,32,31,120,31,120,30,135,31,136,31,126,31,17,31,17,30,17,29,3,31,3,30,82,31,63,31,63,30,63,29,84,31,71,31,141,31,182,31,116,31,91,31,91,30,22,31,13,31,96,31,83,31,127,31,163,31,7,31,215,31,142,31,160,31,109,31,109,30,177,31,40,31,48,31,48,30,238,31,86,31,86,30,86,29,227,31,227,30,227,29,227,28,130,31,18,31,31,31,147,31,147,30,87,31,90,31,253,31,182,31,39,31,18,31,32,31,75,31,238,31,157,31,157,30,232,31,232,31,112,31,112,30,112,29,81,31,254,31,9,31,39,31,194,31,194,30,194,29,165,31,176,31,41,31,41,30,49,31,160,31,160,30,64,31,147,31,52,31,52,31,234,31,109,31,109,30,19,31,209,31,208,31,58,31,183,31,183,30,229,31,234,31,22,31,187,31,217,31,217,30,41,31,213,31,209,31,127,31,5,31,214,31,214,30,114,31,114,30,52,31,28,31,5,31,175,31,178,31,134,31,42,31,29,31,29,30,71,31,202,31,177,31,105,31,172,31,148,31,31,31,193,31,70,31,130,31,75,31,194,31,39,31,135,31,135,30,214,31,235,31,235,30,136,31,141,31,141,30,99,31,99,30,171,31,31,31,114,31,52,31,29,31,1,31,73,31,212,31,212,30,127,31,99,31,133,31,133,30,126,31,111,31,137,31,222,31,222,30,33,31,216,31,17,31,17,30,167,31,169,31,152,31,114,31,234,31,234,30,249,31,205,31,222,31,83,31,16,31,70,31,144,31,159,31,60,31,20,31,84,31,218,31,218,30,218,29,218,28,218,27,202,31,202,31,202,30,224,31,107,31,226,31,248,31,224,31,224,30,83,31,10,31,62,31,248,31,39,31,172,31,172,30,215,31,196,31,11,31,15,31,15,30,79,31,13,31,186,31,186,30,228,31,228,30,228,29,246,31,160,31,209,31,217,31,147,31,88,31,252,31,250,31,250,30,250,29,58,31,242,31,206,31,93,31,93,30,79,31,94,31,186,31,111,31,44,31,128,31,180,31,16,31,180,31,158,31,158,30,65,31,108,31,206,31,206,30,226,31,226,30,184,31,184,30,32,31,148,31,136,31,193,31,140,31,208,31,208,30,29,31,29,30,29,29,40,31,25,31,118,31,166,31,180,31,209,31,181,31,30,31,178,31,61,31,56,31,228,31,201,31,5,31,194,31,194,30,195,31,195,30,159,31,207,31,227,31,206,31,139,31,101,31,103,31,103,30,32,31,10,31,29,31,134,31,134,31,183,31,94,31,202,31,149,31,15,31,213,31,178,31,244,31,244,30,244,29,244,28,35,31,35,30,206,31,60,31,165,31,214,31,148,31,148,30,148,29,88,31,15,31,195,31,146,31,146,30,146,29,125,31,11,31,240,31,84,31,248,31,128,31,8,31,94,31,94,30,47,31,47,30,54,31,203,31,203,30,216,31,120,31,244,31,111,31,74,31,46,31,103,31,25,31,214,31,217,31,118,31,224,31,228,31,186,31,142,31,123,31,35,31,102,31,101,31,137,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
