-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 334;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (32,0,125,0,29,0,43,0,0,0,0,0,59,0,204,0,190,0,6,0,0,0,44,0,225,0,33,0,96,0,64,0,52,0,0,0,1,0,0,0,221,0,0,0,0,0,0,0,0,0,82,0,147,0,85,0,48,0,19,0,225,0,249,0,138,0,112,0,69,0,31,0,170,0,0,0,57,0,181,0,46,0,58,0,0,0,0,0,40,0,173,0,0,0,229,0,213,0,144,0,139,0,9,0,0,0,15,0,168,0,103,0,20,0,141,0,189,0,232,0,71,0,52,0,97,0,200,0,116,0,110,0,0,0,242,0,0,0,209,0,179,0,28,0,0,0,173,0,41,0,16,0,90,0,185,0,130,0,0,0,209,0,72,0,70,0,177,0,178,0,0,0,101,0,0,0,0,0,0,0,223,0,0,0,32,0,132,0,0,0,154,0,0,0,16,0,229,0,49,0,199,0,245,0,166,0,0,0,93,0,0,0,0,0,135,0,134,0,0,0,170,0,193,0,0,0,131,0,24,0,17,0,101,0,15,0,148,0,250,0,0,0,212,0,102,0,0,0,190,0,67,0,138,0,0,0,0,0,232,0,115,0,100,0,73,0,0,0,0,0,225,0,0,0,232,0,199,0,221,0,90,0,0,0,25,0,108,0,0,0,179,0,9,0,0,0,126,0,113,0,176,0,191,0,46,0,134,0,125,0,28,0,0,0,0,0,97,0,211,0,101,0,36,0,172,0,149,0,220,0,43,0,213,0,229,0,216,0,192,0,11,0,25,0,0,0,25,0,0,0,47,0,220,0,0,0,8,0,0,0,4,0,229,0,0,0,44,0,67,0,103,0,0,0,123,0,0,0,36,0,92,0,71,0,153,0,247,0,151,0,17,0,0,0,124,0,235,0,0,0,6,0,71,0,0,0,42,0,123,0,89,0,71,0,172,0,35,0,114,0,193,0,229,0,0,0,217,0,23,0,255,0,199,0,4,0,133,0,84,0,239,0,0,0,201,0,101,0,0,0,17,0,162,0,249,0,0,0,218,0,196,0,213,0,197,0,24,0,165,0,4,0,9,0,88,0,17,0,147,0,170,0,38,0,67,0,167,0,73,0,55,0,137,0,0,0,87,0,0,0,189,0,205,0,0,0,169,0,104,0,157,0,213,0,125,0,0,0,109,0,9,0,197,0,105,0,0,0,193,0,0,0,124,0,10,0,93,0,238,0,124,0,74,0,190,0,199,0,198,0,81,0,147,0,0,0,0,0,87,0,203,0,0,0,183,0,109,0,248,0,125,0,0,0,90,0,253,0,0,0,0,0,91,0,64,0,2,0,143,0,0,0,127,0,5,0,0,0,39,0,56,0,74,0,119,0,125,0,88,0,243,0,203,0,180,0,0,0,97,0,35,0,126,0,0,0,0,0,75,0,212,0,109,0,1,0,48,0,128,0,63,0,109,0,12,0,23,0,0,0,165,0,140,0,9,0,6,0,251,0,152,0,96,0,174,0,124,0);
signal scenario_full  : scenario_type := (32,31,125,31,29,31,43,31,43,30,43,29,59,31,204,31,190,31,6,31,6,30,44,31,225,31,33,31,96,31,64,31,52,31,52,30,1,31,1,30,221,31,221,30,221,29,221,28,221,27,82,31,147,31,85,31,48,31,19,31,225,31,249,31,138,31,112,31,69,31,31,31,170,31,170,30,57,31,181,31,46,31,58,31,58,30,58,29,40,31,173,31,173,30,229,31,213,31,144,31,139,31,9,31,9,30,15,31,168,31,103,31,20,31,141,31,189,31,232,31,71,31,52,31,97,31,200,31,116,31,110,31,110,30,242,31,242,30,209,31,179,31,28,31,28,30,173,31,41,31,16,31,90,31,185,31,130,31,130,30,209,31,72,31,70,31,177,31,178,31,178,30,101,31,101,30,101,29,101,28,223,31,223,30,32,31,132,31,132,30,154,31,154,30,16,31,229,31,49,31,199,31,245,31,166,31,166,30,93,31,93,30,93,29,135,31,134,31,134,30,170,31,193,31,193,30,131,31,24,31,17,31,101,31,15,31,148,31,250,31,250,30,212,31,102,31,102,30,190,31,67,31,138,31,138,30,138,29,232,31,115,31,100,31,73,31,73,30,73,29,225,31,225,30,232,31,199,31,221,31,90,31,90,30,25,31,108,31,108,30,179,31,9,31,9,30,126,31,113,31,176,31,191,31,46,31,134,31,125,31,28,31,28,30,28,29,97,31,211,31,101,31,36,31,172,31,149,31,220,31,43,31,213,31,229,31,216,31,192,31,11,31,25,31,25,30,25,31,25,30,47,31,220,31,220,30,8,31,8,30,4,31,229,31,229,30,44,31,67,31,103,31,103,30,123,31,123,30,36,31,92,31,71,31,153,31,247,31,151,31,17,31,17,30,124,31,235,31,235,30,6,31,71,31,71,30,42,31,123,31,89,31,71,31,172,31,35,31,114,31,193,31,229,31,229,30,217,31,23,31,255,31,199,31,4,31,133,31,84,31,239,31,239,30,201,31,101,31,101,30,17,31,162,31,249,31,249,30,218,31,196,31,213,31,197,31,24,31,165,31,4,31,9,31,88,31,17,31,147,31,170,31,38,31,67,31,167,31,73,31,55,31,137,31,137,30,87,31,87,30,189,31,205,31,205,30,169,31,104,31,157,31,213,31,125,31,125,30,109,31,9,31,197,31,105,31,105,30,193,31,193,30,124,31,10,31,93,31,238,31,124,31,74,31,190,31,199,31,198,31,81,31,147,31,147,30,147,29,87,31,203,31,203,30,183,31,109,31,248,31,125,31,125,30,90,31,253,31,253,30,253,29,91,31,64,31,2,31,143,31,143,30,127,31,5,31,5,30,39,31,56,31,74,31,119,31,125,31,88,31,243,31,203,31,180,31,180,30,97,31,35,31,126,31,126,30,126,29,75,31,212,31,109,31,1,31,48,31,128,31,63,31,109,31,12,31,23,31,23,30,165,31,140,31,9,31,6,31,251,31,152,31,96,31,174,31,124,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
