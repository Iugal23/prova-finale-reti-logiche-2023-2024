-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 857;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (230,0,0,0,7,0,29,0,60,0,168,0,10,0,73,0,228,0,0,0,184,0,130,0,162,0,0,0,47,0,65,0,0,0,152,0,126,0,248,0,0,0,78,0,0,0,108,0,119,0,158,0,40,0,239,0,116,0,224,0,158,0,40,0,167,0,23,0,122,0,234,0,235,0,11,0,206,0,202,0,165,0,150,0,48,0,73,0,116,0,185,0,220,0,216,0,224,0,238,0,38,0,0,0,134,0,43,0,165,0,198,0,116,0,6,0,44,0,78,0,4,0,25,0,145,0,74,0,63,0,64,0,158,0,121,0,0,0,169,0,0,0,233,0,98,0,120,0,122,0,242,0,43,0,0,0,80,0,69,0,90,0,0,0,0,0,255,0,8,0,0,0,172,0,0,0,127,0,124,0,53,0,233,0,249,0,94,0,0,0,20,0,21,0,173,0,88,0,0,0,105,0,113,0,125,0,116,0,93,0,50,0,104,0,3,0,96,0,234,0,84,0,0,0,214,0,64,0,0,0,167,0,70,0,0,0,193,0,66,0,0,0,121,0,42,0,28,0,0,0,234,0,217,0,91,0,0,0,225,0,0,0,0,0,0,0,43,0,64,0,87,0,64,0,51,0,16,0,2,0,147,0,243,0,242,0,59,0,18,0,146,0,3,0,76,0,135,0,167,0,69,0,107,0,0,0,180,0,117,0,0,0,225,0,224,0,183,0,128,0,122,0,172,0,58,0,140,0,0,0,190,0,125,0,33,0,7,0,39,0,0,0,130,0,79,0,62,0,154,0,141,0,156,0,0,0,106,0,94,0,114,0,212,0,230,0,166,0,83,0,191,0,0,0,0,0,142,0,0,0,19,0,196,0,0,0,224,0,0,0,60,0,56,0,0,0,0,0,142,0,0,0,138,0,93,0,0,0,135,0,141,0,238,0,36,0,168,0,142,0,0,0,129,0,155,0,106,0,18,0,197,0,24,0,0,0,193,0,154,0,203,0,155,0,17,0,215,0,0,0,45,0,0,0,95,0,173,0,150,0,0,0,40,0,253,0,30,0,252,0,78,0,255,0,193,0,205,0,227,0,108,0,187,0,241,0,239,0,0,0,43,0,125,0,239,0,166,0,63,0,96,0,154,0,0,0,76,0,15,0,72,0,177,0,177,0,13,0,139,0,0,0,3,0,73,0,0,0,175,0,0,0,0,0,199,0,115,0,216,0,233,0,223,0,44,0,125,0,165,0,0,0,166,0,71,0,0,0,0,0,146,0,219,0,80,0,152,0,100,0,255,0,66,0,197,0,59,0,158,0,164,0,154,0,132,0,0,0,138,0,113,0,46,0,0,0,53,0,236,0,194,0,228,0,160,0,0,0,169,0,25,0,107,0,141,0,153,0,218,0,0,0,219,0,80,0,150,0,9,0,0,0,37,0,37,0,85,0,191,0,98,0,178,0,133,0,100,0,95,0,0,0,0,0,134,0,202,0,200,0,200,0,0,0,219,0,132,0,77,0,148,0,0,0,46,0,0,0,135,0,191,0,0,0,189,0,111,0,78,0,225,0,0,0,182,0,199,0,248,0,174,0,62,0,36,0,243,0,75,0,33,0,0,0,90,0,18,0,253,0,113,0,10,0,126,0,0,0,55,0,233,0,0,0,102,0,92,0,0,0,0,0,51,0,0,0,10,0,224,0,0,0,60,0,22,0,59,0,0,0,232,0,8,0,208,0,43,0,166,0,0,0,98,0,118,0,95,0,0,0,151,0,75,0,61,0,27,0,241,0,216,0,254,0,90,0,78,0,0,0,26,0,7,0,117,0,37,0,192,0,17,0,34,0,170,0,177,0,228,0,230,0,70,0,250,0,137,0,108,0,190,0,128,0,242,0,0,0,84,0,116,0,108,0,38,0,243,0,248,0,72,0,114,0,86,0,37,0,139,0,214,0,140,0,160,0,192,0,237,0,0,0,136,0,0,0,5,0,69,0,234,0,0,0,0,0,98,0,248,0,63,0,205,0,185,0,7,0,199,0,250,0,146,0,0,0,0,0,128,0,95,0,97,0,68,0,92,0,144,0,242,0,60,0,39,0,60,0,150,0,205,0,224,0,35,0,229,0,248,0,0,0,0,0,17,0,226,0,127,0,221,0,13,0,148,0,0,0,122,0,0,0,141,0,149,0,62,0,0,0,0,0,0,0,0,0,162,0,181,0,11,0,195,0,38,0,71,0,140,0,213,0,195,0,152,0,100,0,30,0,193,0,180,0,38,0,204,0,163,0,31,0,28,0,149,0,77,0,4,0,0,0,186,0,220,0,38,0,14,0,68,0,0,0,0,0,230,0,0,0,83,0,85,0,38,0,123,0,31,0,128,0,0,0,153,0,174,0,29,0,161,0,8,0,36,0,0,0,0,0,37,0,120,0,0,0,91,0,0,0,45,0,117,0,0,0,20,0,136,0,100,0,86,0,122,0,64,0,58,0,43,0,0,0,0,0,151,0,178,0,204,0,199,0,155,0,95,0,85,0,218,0,73,0,216,0,0,0,151,0,85,0,243,0,239,0,139,0,12,0,150,0,213,0,127,0,243,0,28,0,0,0,99,0,5,0,134,0,0,0,4,0,185,0,90,0,184,0,0,0,248,0,99,0,178,0,33,0,0,0,83,0,126,0,113,0,210,0,125,0,228,0,0,0,161,0,82,0,18,0,30,0,45,0,51,0,93,0,138,0,224,0,0,0,17,0,232,0,96,0,137,0,0,0,142,0,148,0,217,0,150,0,189,0,0,0,36,0,237,0,24,0,96,0,237,0,8,0,5,0,0,0,235,0,179,0,123,0,115,0,103,0,0,0,84,0,95,0,57,0,94,0,197,0,54,0,0,0,88,0,40,0,1,0,181,0,238,0,25,0,213,0,0,0,108,0,0,0,196,0,36,0,235,0,0,0,0,0,0,0,114,0,187,0,96,0,44,0,0,0,134,0,30,0,207,0,221,0,0,0,0,0,40,0,65,0,98,0,255,0,150,0,100,0,94,0,176,0,228,0,0,0,98,0,63,0,146,0,142,0,0,0,0,0,65,0,0,0,74,0,49,0,162,0,0,0,255,0,179,0,154,0,27,0,66,0,15,0,189,0,223,0,31,0,103,0,223,0,0,0,0,0,236,0,126,0,16,0,151,0,217,0,123,0,24,0,16,0,135,0,186,0,19,0,217,0,0,0,247,0,67,0,26,0,82,0,240,0,0,0,75,0,0,0,132,0,195,0,121,0,18,0,90,0,196,0,211,0,110,0,133,0,197,0,12,0,172,0,240,0,80,0,35,0,169,0,89,0,0,0,149,0,0,0,0,0,238,0,141,0,251,0,131,0,155,0,63,0,0,0,0,0,99,0,245,0,166,0,200,0,0,0,194,0,250,0,238,0,134,0,189,0,149,0,132,0,53,0,28,0,128,0,160,0,220,0,61,0,120,0,118,0,144,0,187,0,0,0,78,0,28,0,108,0,0,0,241,0,242,0,161,0,162,0,187,0,0,0,221,0,158,0,251,0,197,0,66,0,0,0,131,0,106,0,43,0,0,0,165,0,22,0,72,0,239,0,204,0,0,0,23,0,0,0,175,0,249,0,48,0,181,0,0,0,0,0,86,0,0,0,0,0,30,0,0,0,0,0,139,0,220,0,137,0,189,0,0,0,68,0,109,0,108,0,13,0,26,0,132,0,0,0,11,0,131,0,0,0,0,0,48,0,195,0,89,0,144,0,54,0,113,0,192,0,24,0,11,0,0,0,99,0,242,0,136,0,0,0,222,0,176,0,0,0,0,0,173,0,217,0,0,0,41,0,0,0,9,0,0,0,0,0,52,0);
signal scenario_full  : scenario_type := (230,31,230,30,7,31,29,31,60,31,168,31,10,31,73,31,228,31,228,30,184,31,130,31,162,31,162,30,47,31,65,31,65,30,152,31,126,31,248,31,248,30,78,31,78,30,108,31,119,31,158,31,40,31,239,31,116,31,224,31,158,31,40,31,167,31,23,31,122,31,234,31,235,31,11,31,206,31,202,31,165,31,150,31,48,31,73,31,116,31,185,31,220,31,216,31,224,31,238,31,38,31,38,30,134,31,43,31,165,31,198,31,116,31,6,31,44,31,78,31,4,31,25,31,145,31,74,31,63,31,64,31,158,31,121,31,121,30,169,31,169,30,233,31,98,31,120,31,122,31,242,31,43,31,43,30,80,31,69,31,90,31,90,30,90,29,255,31,8,31,8,30,172,31,172,30,127,31,124,31,53,31,233,31,249,31,94,31,94,30,20,31,21,31,173,31,88,31,88,30,105,31,113,31,125,31,116,31,93,31,50,31,104,31,3,31,96,31,234,31,84,31,84,30,214,31,64,31,64,30,167,31,70,31,70,30,193,31,66,31,66,30,121,31,42,31,28,31,28,30,234,31,217,31,91,31,91,30,225,31,225,30,225,29,225,28,43,31,64,31,87,31,64,31,51,31,16,31,2,31,147,31,243,31,242,31,59,31,18,31,146,31,3,31,76,31,135,31,167,31,69,31,107,31,107,30,180,31,117,31,117,30,225,31,224,31,183,31,128,31,122,31,172,31,58,31,140,31,140,30,190,31,125,31,33,31,7,31,39,31,39,30,130,31,79,31,62,31,154,31,141,31,156,31,156,30,106,31,94,31,114,31,212,31,230,31,166,31,83,31,191,31,191,30,191,29,142,31,142,30,19,31,196,31,196,30,224,31,224,30,60,31,56,31,56,30,56,29,142,31,142,30,138,31,93,31,93,30,135,31,141,31,238,31,36,31,168,31,142,31,142,30,129,31,155,31,106,31,18,31,197,31,24,31,24,30,193,31,154,31,203,31,155,31,17,31,215,31,215,30,45,31,45,30,95,31,173,31,150,31,150,30,40,31,253,31,30,31,252,31,78,31,255,31,193,31,205,31,227,31,108,31,187,31,241,31,239,31,239,30,43,31,125,31,239,31,166,31,63,31,96,31,154,31,154,30,76,31,15,31,72,31,177,31,177,31,13,31,139,31,139,30,3,31,73,31,73,30,175,31,175,30,175,29,199,31,115,31,216,31,233,31,223,31,44,31,125,31,165,31,165,30,166,31,71,31,71,30,71,29,146,31,219,31,80,31,152,31,100,31,255,31,66,31,197,31,59,31,158,31,164,31,154,31,132,31,132,30,138,31,113,31,46,31,46,30,53,31,236,31,194,31,228,31,160,31,160,30,169,31,25,31,107,31,141,31,153,31,218,31,218,30,219,31,80,31,150,31,9,31,9,30,37,31,37,31,85,31,191,31,98,31,178,31,133,31,100,31,95,31,95,30,95,29,134,31,202,31,200,31,200,31,200,30,219,31,132,31,77,31,148,31,148,30,46,31,46,30,135,31,191,31,191,30,189,31,111,31,78,31,225,31,225,30,182,31,199,31,248,31,174,31,62,31,36,31,243,31,75,31,33,31,33,30,90,31,18,31,253,31,113,31,10,31,126,31,126,30,55,31,233,31,233,30,102,31,92,31,92,30,92,29,51,31,51,30,10,31,224,31,224,30,60,31,22,31,59,31,59,30,232,31,8,31,208,31,43,31,166,31,166,30,98,31,118,31,95,31,95,30,151,31,75,31,61,31,27,31,241,31,216,31,254,31,90,31,78,31,78,30,26,31,7,31,117,31,37,31,192,31,17,31,34,31,170,31,177,31,228,31,230,31,70,31,250,31,137,31,108,31,190,31,128,31,242,31,242,30,84,31,116,31,108,31,38,31,243,31,248,31,72,31,114,31,86,31,37,31,139,31,214,31,140,31,160,31,192,31,237,31,237,30,136,31,136,30,5,31,69,31,234,31,234,30,234,29,98,31,248,31,63,31,205,31,185,31,7,31,199,31,250,31,146,31,146,30,146,29,128,31,95,31,97,31,68,31,92,31,144,31,242,31,60,31,39,31,60,31,150,31,205,31,224,31,35,31,229,31,248,31,248,30,248,29,17,31,226,31,127,31,221,31,13,31,148,31,148,30,122,31,122,30,141,31,149,31,62,31,62,30,62,29,62,28,62,27,162,31,181,31,11,31,195,31,38,31,71,31,140,31,213,31,195,31,152,31,100,31,30,31,193,31,180,31,38,31,204,31,163,31,31,31,28,31,149,31,77,31,4,31,4,30,186,31,220,31,38,31,14,31,68,31,68,30,68,29,230,31,230,30,83,31,85,31,38,31,123,31,31,31,128,31,128,30,153,31,174,31,29,31,161,31,8,31,36,31,36,30,36,29,37,31,120,31,120,30,91,31,91,30,45,31,117,31,117,30,20,31,136,31,100,31,86,31,122,31,64,31,58,31,43,31,43,30,43,29,151,31,178,31,204,31,199,31,155,31,95,31,85,31,218,31,73,31,216,31,216,30,151,31,85,31,243,31,239,31,139,31,12,31,150,31,213,31,127,31,243,31,28,31,28,30,99,31,5,31,134,31,134,30,4,31,185,31,90,31,184,31,184,30,248,31,99,31,178,31,33,31,33,30,83,31,126,31,113,31,210,31,125,31,228,31,228,30,161,31,82,31,18,31,30,31,45,31,51,31,93,31,138,31,224,31,224,30,17,31,232,31,96,31,137,31,137,30,142,31,148,31,217,31,150,31,189,31,189,30,36,31,237,31,24,31,96,31,237,31,8,31,5,31,5,30,235,31,179,31,123,31,115,31,103,31,103,30,84,31,95,31,57,31,94,31,197,31,54,31,54,30,88,31,40,31,1,31,181,31,238,31,25,31,213,31,213,30,108,31,108,30,196,31,36,31,235,31,235,30,235,29,235,28,114,31,187,31,96,31,44,31,44,30,134,31,30,31,207,31,221,31,221,30,221,29,40,31,65,31,98,31,255,31,150,31,100,31,94,31,176,31,228,31,228,30,98,31,63,31,146,31,142,31,142,30,142,29,65,31,65,30,74,31,49,31,162,31,162,30,255,31,179,31,154,31,27,31,66,31,15,31,189,31,223,31,31,31,103,31,223,31,223,30,223,29,236,31,126,31,16,31,151,31,217,31,123,31,24,31,16,31,135,31,186,31,19,31,217,31,217,30,247,31,67,31,26,31,82,31,240,31,240,30,75,31,75,30,132,31,195,31,121,31,18,31,90,31,196,31,211,31,110,31,133,31,197,31,12,31,172,31,240,31,80,31,35,31,169,31,89,31,89,30,149,31,149,30,149,29,238,31,141,31,251,31,131,31,155,31,63,31,63,30,63,29,99,31,245,31,166,31,200,31,200,30,194,31,250,31,238,31,134,31,189,31,149,31,132,31,53,31,28,31,128,31,160,31,220,31,61,31,120,31,118,31,144,31,187,31,187,30,78,31,28,31,108,31,108,30,241,31,242,31,161,31,162,31,187,31,187,30,221,31,158,31,251,31,197,31,66,31,66,30,131,31,106,31,43,31,43,30,165,31,22,31,72,31,239,31,204,31,204,30,23,31,23,30,175,31,249,31,48,31,181,31,181,30,181,29,86,31,86,30,86,29,30,31,30,30,30,29,139,31,220,31,137,31,189,31,189,30,68,31,109,31,108,31,13,31,26,31,132,31,132,30,11,31,131,31,131,30,131,29,48,31,195,31,89,31,144,31,54,31,113,31,192,31,24,31,11,31,11,30,99,31,242,31,136,31,136,30,222,31,176,31,176,30,176,29,173,31,217,31,217,30,41,31,41,30,9,31,9,30,9,29,52,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
