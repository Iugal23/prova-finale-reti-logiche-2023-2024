-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 777;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,128,0,124,0,150,0,0,0,194,0,182,0,237,0,184,0,0,0,224,0,0,0,0,0,156,0,70,0,0,0,118,0,182,0,221,0,83,0,150,0,168,0,242,0,37,0,78,0,192,0,77,0,82,0,69,0,109,0,22,0,20,0,37,0,69,0,0,0,0,0,0,0,226,0,0,0,30,0,236,0,117,0,238,0,137,0,117,0,66,0,9,0,78,0,117,0,0,0,172,0,177,0,123,0,68,0,117,0,223,0,179,0,52,0,118,0,126,0,196,0,108,0,101,0,68,0,110,0,254,0,55,0,251,0,114,0,102,0,137,0,24,0,221,0,0,0,239,0,189,0,226,0,0,0,213,0,36,0,109,0,111,0,85,0,18,0,148,0,230,0,0,0,0,0,215,0,174,0,64,0,93,0,0,0,94,0,102,0,104,0,234,0,57,0,0,0,109,0,229,0,99,0,168,0,137,0,251,0,141,0,0,0,0,0,179,0,184,0,0,0,131,0,107,0,59,0,14,0,0,0,190,0,66,0,57,0,134,0,182,0,0,0,96,0,199,0,247,0,63,0,212,0,17,0,8,0,202,0,10,0,157,0,120,0,0,0,1,0,170,0,0,0,0,0,130,0,0,0,178,0,232,0,30,0,0,0,131,0,147,0,136,0,82,0,186,0,25,0,0,0,37,0,236,0,0,0,0,0,0,0,119,0,75,0,90,0,87,0,0,0,215,0,247,0,138,0,239,0,156,0,68,0,11,0,54,0,163,0,214,0,73,0,88,0,11,0,0,0,85,0,236,0,94,0,43,0,147,0,49,0,0,0,121,0,0,0,110,0,75,0,43,0,7,0,92,0,27,0,0,0,223,0,214,0,148,0,141,0,147,0,0,0,224,0,236,0,115,0,0,0,19,0,0,0,22,0,120,0,49,0,37,0,69,0,100,0,213,0,221,0,146,0,245,0,204,0,0,0,27,0,82,0,168,0,107,0,144,0,206,0,0,0,0,0,0,0,145,0,0,0,186,0,140,0,132,0,216,0,0,0,228,0,185,0,14,0,193,0,207,0,9,0,210,0,21,0,55,0,0,0,100,0,227,0,21,0,236,0,71,0,214,0,39,0,0,0,14,0,149,0,116,0,0,0,0,0,62,0,18,0,138,0,198,0,0,0,81,0,213,0,177,0,73,0,155,0,0,0,80,0,249,0,151,0,0,0,57,0,7,0,25,0,0,0,0,0,200,0,229,0,39,0,237,0,201,0,47,0,211,0,40,0,0,0,178,0,164,0,28,0,0,0,154,0,201,0,26,0,4,0,213,0,71,0,118,0,217,0,130,0,62,0,166,0,109,0,239,0,246,0,76,0,0,0,13,0,0,0,55,0,0,0,14,0,0,0,49,0,89,0,217,0,229,0,96,0,124,0,249,0,0,0,3,0,211,0,78,0,107,0,21,0,167,0,0,0,34,0,0,0,86,0,118,0,64,0,123,0,118,0,104,0,57,0,0,0,19,0,87,0,128,0,177,0,59,0,95,0,183,0,111,0,0,0,184,0,164,0,50,0,0,0,246,0,0,0,0,0,58,0,159,0,81,0,144,0,126,0,58,0,185,0,36,0,250,0,105,0,223,0,132,0,0,0,53,0,21,0,115,0,0,0,61,0,70,0,38,0,140,0,92,0,71,0,254,0,80,0,74,0,119,0,0,0,248,0,179,0,168,0,26,0,109,0,0,0,145,0,122,0,0,0,0,0,67,0,118,0,242,0,0,0,34,0,0,0,40,0,104,0,14,0,139,0,18,0,0,0,74,0,0,0,22,0,35,0,0,0,81,0,59,0,17,0,136,0,6,0,232,0,46,0,202,0,0,0,87,0,209,0,196,0,230,0,46,0,0,0,136,0,52,0,57,0,69,0,0,0,191,0,155,0,215,0,192,0,119,0,0,0,248,0,182,0,41,0,232,0,62,0,63,0,123,0,235,0,121,0,111,0,104,0,141,0,0,0,85,0,0,0,0,0,0,0,21,0,16,0,0,0,175,0,0,0,56,0,45,0,6,0,41,0,5,0,0,0,113,0,119,0,163,0,238,0,141,0,221,0,0,0,18,0,97,0,243,0,208,0,233,0,238,0,133,0,36,0,136,0,249,0,0,0,0,0,240,0,93,0,38,0,175,0,39,0,101,0,148,0,0,0,229,0,39,0,0,0,225,0,118,0,0,0,59,0,30,0,0,0,199,0,130,0,40,0,73,0,212,0,0,0,204,0,40,0,124,0,0,0,22,0,219,0,119,0,66,0,42,0,212,0,0,0,65,0,0,0,0,0,125,0,51,0,8,0,72,0,12,0,164,0,214,0,0,0,158,0,0,0,0,0,255,0,11,0,12,0,179,0,14,0,224,0,0,0,0,0,0,0,225,0,17,0,229,0,175,0,0,0,177,0,152,0,11,0,143,0,0,0,134,0,98,0,202,0,0,0,50,0,0,0,250,0,0,0,252,0,150,0,95,0,0,0,190,0,194,0,228,0,0,0,231,0,114,0,19,0,0,0,198,0,250,0,0,0,123,0,20,0,186,0,0,0,250,0,164,0,83,0,41,0,0,0,67,0,0,0,74,0,0,0,156,0,51,0,67,0,152,0,0,0,15,0,240,0,51,0,0,0,11,0,153,0,212,0,144,0,165,0,24,0,236,0,157,0,255,0,205,0,3,0,162,0,38,0,202,0,0,0,23,0,98,0,0,0,0,0,239,0,209,0,0,0,195,0,66,0,137,0,0,0,187,0,98,0,209,0,40,0,62,0,167,0,0,0,73,0,214,0,0,0,0,0,168,0,0,0,188,0,0,0,168,0,0,0,0,0,122,0,105,0,102,0,144,0,23,0,39,0,0,0,220,0,207,0,4,0,45,0,190,0,0,0,9,0,192,0,244,0,242,0,108,0,23,0,3,0,0,0,164,0,78,0,249,0,219,0,0,0,206,0,57,0,13,0,46,0,23,0,20,0,104,0,0,0,141,0,14,0,158,0,136,0,225,0,242,0,0,0,215,0,247,0,10,0,0,0,64,0,255,0,233,0,235,0,177,0,191,0,90,0,192,0,129,0,0,0,0,0,135,0,121,0,178,0,69,0,0,0,81,0,99,0,100,0,209,0,108,0,204,0,232,0,89,0,235,0,193,0,235,0,252,0,159,0,229,0,59,0,0,0,190,0,207,0,96,0,51,0,4,0,12,0,28,0,213,0,0,0,93,0,0,0,0,0,32,0,0,0,222,0,177,0,34,0,106,0,171,0,212,0,72,0,144,0,92,0,247,0,20,0,85,0,0,0,167,0,74,0,0,0,219,0,114,0,0,0,181,0,22,0,232,0,0,0,0,0,239,0,202,0,145,0,56,0,91,0,37,0,87,0,184,0,7,0,2,0,5,0,163,0,0,0,110,0,197,0,7,0,43,0,48,0,46,0,215,0,206,0,244,0,0,0,0,0,197,0,111,0,0,0,158,0);
signal scenario_full  : scenario_type := (0,0,128,31,124,31,150,31,150,30,194,31,182,31,237,31,184,31,184,30,224,31,224,30,224,29,156,31,70,31,70,30,118,31,182,31,221,31,83,31,150,31,168,31,242,31,37,31,78,31,192,31,77,31,82,31,69,31,109,31,22,31,20,31,37,31,69,31,69,30,69,29,69,28,226,31,226,30,30,31,236,31,117,31,238,31,137,31,117,31,66,31,9,31,78,31,117,31,117,30,172,31,177,31,123,31,68,31,117,31,223,31,179,31,52,31,118,31,126,31,196,31,108,31,101,31,68,31,110,31,254,31,55,31,251,31,114,31,102,31,137,31,24,31,221,31,221,30,239,31,189,31,226,31,226,30,213,31,36,31,109,31,111,31,85,31,18,31,148,31,230,31,230,30,230,29,215,31,174,31,64,31,93,31,93,30,94,31,102,31,104,31,234,31,57,31,57,30,109,31,229,31,99,31,168,31,137,31,251,31,141,31,141,30,141,29,179,31,184,31,184,30,131,31,107,31,59,31,14,31,14,30,190,31,66,31,57,31,134,31,182,31,182,30,96,31,199,31,247,31,63,31,212,31,17,31,8,31,202,31,10,31,157,31,120,31,120,30,1,31,170,31,170,30,170,29,130,31,130,30,178,31,232,31,30,31,30,30,131,31,147,31,136,31,82,31,186,31,25,31,25,30,37,31,236,31,236,30,236,29,236,28,119,31,75,31,90,31,87,31,87,30,215,31,247,31,138,31,239,31,156,31,68,31,11,31,54,31,163,31,214,31,73,31,88,31,11,31,11,30,85,31,236,31,94,31,43,31,147,31,49,31,49,30,121,31,121,30,110,31,75,31,43,31,7,31,92,31,27,31,27,30,223,31,214,31,148,31,141,31,147,31,147,30,224,31,236,31,115,31,115,30,19,31,19,30,22,31,120,31,49,31,37,31,69,31,100,31,213,31,221,31,146,31,245,31,204,31,204,30,27,31,82,31,168,31,107,31,144,31,206,31,206,30,206,29,206,28,145,31,145,30,186,31,140,31,132,31,216,31,216,30,228,31,185,31,14,31,193,31,207,31,9,31,210,31,21,31,55,31,55,30,100,31,227,31,21,31,236,31,71,31,214,31,39,31,39,30,14,31,149,31,116,31,116,30,116,29,62,31,18,31,138,31,198,31,198,30,81,31,213,31,177,31,73,31,155,31,155,30,80,31,249,31,151,31,151,30,57,31,7,31,25,31,25,30,25,29,200,31,229,31,39,31,237,31,201,31,47,31,211,31,40,31,40,30,178,31,164,31,28,31,28,30,154,31,201,31,26,31,4,31,213,31,71,31,118,31,217,31,130,31,62,31,166,31,109,31,239,31,246,31,76,31,76,30,13,31,13,30,55,31,55,30,14,31,14,30,49,31,89,31,217,31,229,31,96,31,124,31,249,31,249,30,3,31,211,31,78,31,107,31,21,31,167,31,167,30,34,31,34,30,86,31,118,31,64,31,123,31,118,31,104,31,57,31,57,30,19,31,87,31,128,31,177,31,59,31,95,31,183,31,111,31,111,30,184,31,164,31,50,31,50,30,246,31,246,30,246,29,58,31,159,31,81,31,144,31,126,31,58,31,185,31,36,31,250,31,105,31,223,31,132,31,132,30,53,31,21,31,115,31,115,30,61,31,70,31,38,31,140,31,92,31,71,31,254,31,80,31,74,31,119,31,119,30,248,31,179,31,168,31,26,31,109,31,109,30,145,31,122,31,122,30,122,29,67,31,118,31,242,31,242,30,34,31,34,30,40,31,104,31,14,31,139,31,18,31,18,30,74,31,74,30,22,31,35,31,35,30,81,31,59,31,17,31,136,31,6,31,232,31,46,31,202,31,202,30,87,31,209,31,196,31,230,31,46,31,46,30,136,31,52,31,57,31,69,31,69,30,191,31,155,31,215,31,192,31,119,31,119,30,248,31,182,31,41,31,232,31,62,31,63,31,123,31,235,31,121,31,111,31,104,31,141,31,141,30,85,31,85,30,85,29,85,28,21,31,16,31,16,30,175,31,175,30,56,31,45,31,6,31,41,31,5,31,5,30,113,31,119,31,163,31,238,31,141,31,221,31,221,30,18,31,97,31,243,31,208,31,233,31,238,31,133,31,36,31,136,31,249,31,249,30,249,29,240,31,93,31,38,31,175,31,39,31,101,31,148,31,148,30,229,31,39,31,39,30,225,31,118,31,118,30,59,31,30,31,30,30,199,31,130,31,40,31,73,31,212,31,212,30,204,31,40,31,124,31,124,30,22,31,219,31,119,31,66,31,42,31,212,31,212,30,65,31,65,30,65,29,125,31,51,31,8,31,72,31,12,31,164,31,214,31,214,30,158,31,158,30,158,29,255,31,11,31,12,31,179,31,14,31,224,31,224,30,224,29,224,28,225,31,17,31,229,31,175,31,175,30,177,31,152,31,11,31,143,31,143,30,134,31,98,31,202,31,202,30,50,31,50,30,250,31,250,30,252,31,150,31,95,31,95,30,190,31,194,31,228,31,228,30,231,31,114,31,19,31,19,30,198,31,250,31,250,30,123,31,20,31,186,31,186,30,250,31,164,31,83,31,41,31,41,30,67,31,67,30,74,31,74,30,156,31,51,31,67,31,152,31,152,30,15,31,240,31,51,31,51,30,11,31,153,31,212,31,144,31,165,31,24,31,236,31,157,31,255,31,205,31,3,31,162,31,38,31,202,31,202,30,23,31,98,31,98,30,98,29,239,31,209,31,209,30,195,31,66,31,137,31,137,30,187,31,98,31,209,31,40,31,62,31,167,31,167,30,73,31,214,31,214,30,214,29,168,31,168,30,188,31,188,30,168,31,168,30,168,29,122,31,105,31,102,31,144,31,23,31,39,31,39,30,220,31,207,31,4,31,45,31,190,31,190,30,9,31,192,31,244,31,242,31,108,31,23,31,3,31,3,30,164,31,78,31,249,31,219,31,219,30,206,31,57,31,13,31,46,31,23,31,20,31,104,31,104,30,141,31,14,31,158,31,136,31,225,31,242,31,242,30,215,31,247,31,10,31,10,30,64,31,255,31,233,31,235,31,177,31,191,31,90,31,192,31,129,31,129,30,129,29,135,31,121,31,178,31,69,31,69,30,81,31,99,31,100,31,209,31,108,31,204,31,232,31,89,31,235,31,193,31,235,31,252,31,159,31,229,31,59,31,59,30,190,31,207,31,96,31,51,31,4,31,12,31,28,31,213,31,213,30,93,31,93,30,93,29,32,31,32,30,222,31,177,31,34,31,106,31,171,31,212,31,72,31,144,31,92,31,247,31,20,31,85,31,85,30,167,31,74,31,74,30,219,31,114,31,114,30,181,31,22,31,232,31,232,30,232,29,239,31,202,31,145,31,56,31,91,31,37,31,87,31,184,31,7,31,2,31,5,31,163,31,163,30,110,31,197,31,7,31,43,31,48,31,46,31,215,31,206,31,244,31,244,30,244,29,197,31,111,31,111,30,158,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
