-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 447;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (241,0,83,0,133,0,65,0,228,0,164,0,14,0,203,0,0,0,0,0,20,0,0,0,209,0,24,0,226,0,146,0,84,0,215,0,110,0,91,0,228,0,98,0,240,0,77,0,0,0,17,0,0,0,254,0,0,0,58,0,223,0,50,0,188,0,213,0,6,0,217,0,239,0,224,0,148,0,0,0,0,0,66,0,243,0,166,0,188,0,0,0,0,0,241,0,111,0,2,0,241,0,6,0,214,0,70,0,60,0,69,0,133,0,249,0,206,0,6,0,17,0,216,0,61,0,234,0,25,0,226,0,39,0,53,0,0,0,141,0,138,0,253,0,0,0,121,0,67,0,241,0,0,0,110,0,23,0,97,0,75,0,228,0,0,0,0,0,172,0,25,0,42,0,163,0,0,0,0,0,6,0,135,0,169,0,112,0,0,0,157,0,69,0,28,0,32,0,203,0,114,0,32,0,6,0,122,0,0,0,162,0,222,0,82,0,15,0,163,0,147,0,28,0,0,0,251,0,0,0,143,0,0,0,117,0,164,0,39,0,140,0,30,0,0,0,157,0,87,0,200,0,252,0,51,0,0,0,106,0,70,0,3,0,36,0,162,0,168,0,229,0,0,0,217,0,11,0,223,0,0,0,84,0,242,0,0,0,202,0,143,0,106,0,112,0,157,0,47,0,55,0,188,0,172,0,0,0,8,0,0,0,222,0,233,0,0,0,86,0,16,0,249,0,255,0,113,0,70,0,203,0,0,0,93,0,166,0,85,0,241,0,48,0,247,0,114,0,135,0,189,0,0,0,170,0,245,0,31,0,29,0,207,0,129,0,222,0,195,0,199,0,171,0,234,0,89,0,242,0,124,0,59,0,49,0,220,0,157,0,200,0,0,0,55,0,108,0,124,0,215,0,74,0,160,0,0,0,235,0,42,0,135,0,2,0,144,0,47,0,26,0,230,0,0,0,120,0,1,0,112,0,0,0,236,0,0,0,178,0,242,0,79,0,41,0,249,0,0,0,198,0,0,0,150,0,42,0,218,0,28,0,0,0,94,0,155,0,0,0,147,0,0,0,0,0,77,0,39,0,9,0,51,0,137,0,97,0,0,0,68,0,193,0,109,0,227,0,64,0,0,0,184,0,79,0,186,0,0,0,138,0,226,0,123,0,143,0,175,0,108,0,82,0,138,0,149,0,255,0,253,0,192,0,0,0,0,0,146,0,0,0,98,0,63,0,0,0,215,0,63,0,87,0,125,0,137,0,178,0,156,0,0,0,79,0,208,0,197,0,242,0,0,0,50,0,163,0,0,0,68,0,7,0,40,0,0,0,220,0,173,0,251,0,37,0,189,0,91,0,60,0,107,0,0,0,94,0,193,0,53,0,5,0,106,0,0,0,0,0,0,0,19,0,0,0,0,0,145,0,0,0,124,0,156,0,82,0,211,0,145,0,37,0,150,0,118,0,187,0,251,0,32,0,1,0,249,0,236,0,0,0,134,0,158,0,206,0,226,0,0,0,87,0,0,0,0,0,234,0,136,0,195,0,219,0,61,0,5,0,228,0,230,0,208,0,0,0,114,0,26,0,202,0,49,0,44,0,76,0,113,0,237,0,221,0,0,0,128,0,215,0,17,0,87,0,0,0,21,0,215,0,0,0,238,0,0,0,243,0,140,0,157,0,98,0,209,0,0,0,173,0,0,0,0,0,1,0,181,0,195,0,136,0,221,0,188,0,72,0,245,0,43,0,84,0,162,0,130,0,146,0,29,0,1,0,0,0,140,0,50,0,110,0,82,0,244,0,129,0,23,0,0,0,0,0,94,0,60,0,0,0,104,0,150,0,1,0,70,0,8,0,128,0,0,0,18,0,0,0,66,0,0,0,137,0,218,0,23,0,91,0,185,0,47,0,40,0,1,0,219,0,73,0,111,0,0,0,190,0,101,0,0,0,180,0,94,0,71,0,0,0,137,0,36,0,197,0,136,0,235,0,144,0,44,0,0,0,49,0,108,0,160,0);
signal scenario_full  : scenario_type := (241,31,83,31,133,31,65,31,228,31,164,31,14,31,203,31,203,30,203,29,20,31,20,30,209,31,24,31,226,31,146,31,84,31,215,31,110,31,91,31,228,31,98,31,240,31,77,31,77,30,17,31,17,30,254,31,254,30,58,31,223,31,50,31,188,31,213,31,6,31,217,31,239,31,224,31,148,31,148,30,148,29,66,31,243,31,166,31,188,31,188,30,188,29,241,31,111,31,2,31,241,31,6,31,214,31,70,31,60,31,69,31,133,31,249,31,206,31,6,31,17,31,216,31,61,31,234,31,25,31,226,31,39,31,53,31,53,30,141,31,138,31,253,31,253,30,121,31,67,31,241,31,241,30,110,31,23,31,97,31,75,31,228,31,228,30,228,29,172,31,25,31,42,31,163,31,163,30,163,29,6,31,135,31,169,31,112,31,112,30,157,31,69,31,28,31,32,31,203,31,114,31,32,31,6,31,122,31,122,30,162,31,222,31,82,31,15,31,163,31,147,31,28,31,28,30,251,31,251,30,143,31,143,30,117,31,164,31,39,31,140,31,30,31,30,30,157,31,87,31,200,31,252,31,51,31,51,30,106,31,70,31,3,31,36,31,162,31,168,31,229,31,229,30,217,31,11,31,223,31,223,30,84,31,242,31,242,30,202,31,143,31,106,31,112,31,157,31,47,31,55,31,188,31,172,31,172,30,8,31,8,30,222,31,233,31,233,30,86,31,16,31,249,31,255,31,113,31,70,31,203,31,203,30,93,31,166,31,85,31,241,31,48,31,247,31,114,31,135,31,189,31,189,30,170,31,245,31,31,31,29,31,207,31,129,31,222,31,195,31,199,31,171,31,234,31,89,31,242,31,124,31,59,31,49,31,220,31,157,31,200,31,200,30,55,31,108,31,124,31,215,31,74,31,160,31,160,30,235,31,42,31,135,31,2,31,144,31,47,31,26,31,230,31,230,30,120,31,1,31,112,31,112,30,236,31,236,30,178,31,242,31,79,31,41,31,249,31,249,30,198,31,198,30,150,31,42,31,218,31,28,31,28,30,94,31,155,31,155,30,147,31,147,30,147,29,77,31,39,31,9,31,51,31,137,31,97,31,97,30,68,31,193,31,109,31,227,31,64,31,64,30,184,31,79,31,186,31,186,30,138,31,226,31,123,31,143,31,175,31,108,31,82,31,138,31,149,31,255,31,253,31,192,31,192,30,192,29,146,31,146,30,98,31,63,31,63,30,215,31,63,31,87,31,125,31,137,31,178,31,156,31,156,30,79,31,208,31,197,31,242,31,242,30,50,31,163,31,163,30,68,31,7,31,40,31,40,30,220,31,173,31,251,31,37,31,189,31,91,31,60,31,107,31,107,30,94,31,193,31,53,31,5,31,106,31,106,30,106,29,106,28,19,31,19,30,19,29,145,31,145,30,124,31,156,31,82,31,211,31,145,31,37,31,150,31,118,31,187,31,251,31,32,31,1,31,249,31,236,31,236,30,134,31,158,31,206,31,226,31,226,30,87,31,87,30,87,29,234,31,136,31,195,31,219,31,61,31,5,31,228,31,230,31,208,31,208,30,114,31,26,31,202,31,49,31,44,31,76,31,113,31,237,31,221,31,221,30,128,31,215,31,17,31,87,31,87,30,21,31,215,31,215,30,238,31,238,30,243,31,140,31,157,31,98,31,209,31,209,30,173,31,173,30,173,29,1,31,181,31,195,31,136,31,221,31,188,31,72,31,245,31,43,31,84,31,162,31,130,31,146,31,29,31,1,31,1,30,140,31,50,31,110,31,82,31,244,31,129,31,23,31,23,30,23,29,94,31,60,31,60,30,104,31,150,31,1,31,70,31,8,31,128,31,128,30,18,31,18,30,66,31,66,30,137,31,218,31,23,31,91,31,185,31,47,31,40,31,1,31,219,31,73,31,111,31,111,30,190,31,101,31,101,30,180,31,94,31,71,31,71,30,137,31,36,31,197,31,136,31,235,31,144,31,44,31,44,30,49,31,108,31,160,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
