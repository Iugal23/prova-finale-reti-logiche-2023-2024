-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_56 is
end project_tb_56;

architecture project_tb_arch_56 of project_tb_56 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 221;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (9,0,1,0,0,0,245,0,1,0,239,0,232,0,223,0,14,0,85,0,37,0,171,0,90,0,97,0,252,0,38,0,55,0,135,0,0,0,196,0,0,0,153,0,191,0,194,0,85,0,0,0,7,0,0,0,34,0,199,0,93,0,104,0,0,0,0,0,207,0,122,0,76,0,37,0,0,0,113,0,64,0,214,0,122,0,5,0,139,0,200,0,0,0,0,0,87,0,123,0,216,0,0,0,184,0,217,0,248,0,160,0,12,0,111,0,0,0,0,0,146,0,130,0,208,0,0,0,130,0,145,0,114,0,200,0,173,0,189,0,119,0,93,0,101,0,24,0,0,0,237,0,78,0,162,0,88,0,144,0,0,0,63,0,189,0,162,0,198,0,202,0,235,0,77,0,0,0,129,0,0,0,79,0,0,0,0,0,12,0,202,0,43,0,199,0,188,0,0,0,0,0,78,0,244,0,0,0,121,0,189,0,0,0,0,0,9,0,101,0,115,0,53,0,29,0,102,0,0,0,73,0,221,0,203,0,0,0,0,0,251,0,229,0,0,0,25,0,0,0,27,0,108,0,0,0,147,0,31,0,0,0,0,0,1,0,95,0,96,0,0,0,89,0,211,0,75,0,150,0,201,0,0,0,62,0,239,0,61,0,7,0,0,0,59,0,245,0,161,0,0,0,40,0,2,0,0,0,171,0,18,0,193,0,183,0,254,0,45,0,236,0,0,0,107,0,131,0,117,0,33,0,0,0,149,0,223,0,106,0,19,0,97,0,128,0,90,0,0,0,25,0,4,0,16,0,55,0,137,0,74,0,122,0,149,0,123,0,13,0,223,0,235,0,12,0,202,0,171,0,88,0,34,0,107,0,176,0,92,0,70,0,110,0,42,0,229,0,164,0,53,0,137,0,172,0,170,0,253,0,0,0,224,0,69,0,103,0,26,0,19,0,47,0,0,0,61,0,220,0,130,0,237,0,92,0,173,0,145,0,68,0);
signal scenario_full  : scenario_type := (9,31,1,31,1,30,245,31,1,31,239,31,232,31,223,31,14,31,85,31,37,31,171,31,90,31,97,31,252,31,38,31,55,31,135,31,135,30,196,31,196,30,153,31,191,31,194,31,85,31,85,30,7,31,7,30,34,31,199,31,93,31,104,31,104,30,104,29,207,31,122,31,76,31,37,31,37,30,113,31,64,31,214,31,122,31,5,31,139,31,200,31,200,30,200,29,87,31,123,31,216,31,216,30,184,31,217,31,248,31,160,31,12,31,111,31,111,30,111,29,146,31,130,31,208,31,208,30,130,31,145,31,114,31,200,31,173,31,189,31,119,31,93,31,101,31,24,31,24,30,237,31,78,31,162,31,88,31,144,31,144,30,63,31,189,31,162,31,198,31,202,31,235,31,77,31,77,30,129,31,129,30,79,31,79,30,79,29,12,31,202,31,43,31,199,31,188,31,188,30,188,29,78,31,244,31,244,30,121,31,189,31,189,30,189,29,9,31,101,31,115,31,53,31,29,31,102,31,102,30,73,31,221,31,203,31,203,30,203,29,251,31,229,31,229,30,25,31,25,30,27,31,108,31,108,30,147,31,31,31,31,30,31,29,1,31,95,31,96,31,96,30,89,31,211,31,75,31,150,31,201,31,201,30,62,31,239,31,61,31,7,31,7,30,59,31,245,31,161,31,161,30,40,31,2,31,2,30,171,31,18,31,193,31,183,31,254,31,45,31,236,31,236,30,107,31,131,31,117,31,33,31,33,30,149,31,223,31,106,31,19,31,97,31,128,31,90,31,90,30,25,31,4,31,16,31,55,31,137,31,74,31,122,31,149,31,123,31,13,31,223,31,235,31,12,31,202,31,171,31,88,31,34,31,107,31,176,31,92,31,70,31,110,31,42,31,229,31,164,31,53,31,137,31,172,31,170,31,253,31,253,30,224,31,69,31,103,31,26,31,19,31,47,31,47,30,61,31,220,31,130,31,237,31,92,31,173,31,145,31,68,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
