-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_173 is
end project_tb_173;

architecture project_tb_arch_173 of project_tb_173 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 662;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,17,0,225,0,0,0,162,0,0,0,0,0,240,0,192,0,207,0,0,0,0,0,93,0,134,0,218,0,41,0,0,0,0,0,49,0,235,0,243,0,90,0,109,0,57,0,0,0,225,0,232,0,185,0,72,0,223,0,69,0,150,0,61,0,61,0,226,0,125,0,53,0,255,0,97,0,82,0,174,0,50,0,132,0,89,0,117,0,0,0,204,0,194,0,27,0,179,0,229,0,60,0,253,0,60,0,180,0,0,0,207,0,105,0,229,0,0,0,43,0,31,0,192,0,134,0,0,0,187,0,9,0,49,0,64,0,246,0,233,0,162,0,113,0,0,0,150,0,0,0,241,0,127,0,203,0,72,0,254,0,66,0,149,0,160,0,251,0,62,0,224,0,195,0,187,0,10,0,252,0,79,0,194,0,51,0,0,0,23,0,170,0,7,0,224,0,0,0,230,0,0,0,233,0,0,0,65,0,169,0,137,0,0,0,60,0,0,0,162,0,188,0,0,0,131,0,195,0,8,0,42,0,58,0,181,0,234,0,173,0,213,0,0,0,89,0,94,0,76,0,81,0,204,0,224,0,205,0,0,0,51,0,0,0,226,0,177,0,139,0,56,0,198,0,205,0,25,0,114,0,122,0,215,0,0,0,0,0,54,0,21,0,238,0,0,0,143,0,177,0,201,0,38,0,151,0,180,0,0,0,122,0,213,0,90,0,0,0,162,0,219,0,0,0,2,0,43,0,129,0,29,0,89,0,94,0,140,0,34,0,254,0,0,0,156,0,30,0,0,0,122,0,11,0,0,0,0,0,0,0,133,0,173,0,143,0,67,0,51,0,222,0,212,0,196,0,12,0,0,0,187,0,239,0,105,0,0,0,55,0,0,0,119,0,0,0,132,0,249,0,104,0,0,0,203,0,48,0,18,0,125,0,186,0,185,0,0,0,53,0,0,0,252,0,0,0,255,0,0,0,143,0,117,0,214,0,66,0,0,0,0,0,0,0,30,0,63,0,8,0,0,0,171,0,0,0,0,0,212,0,57,0,80,0,0,0,158,0,37,0,199,0,216,0,112,0,244,0,0,0,165,0,160,0,117,0,203,0,237,0,71,0,241,0,58,0,93,0,35,0,165,0,110,0,0,0,0,0,172,0,96,0,0,0,0,0,170,0,43,0,239,0,146,0,196,0,8,0,127,0,0,0,125,0,128,0,0,0,252,0,174,0,252,0,104,0,0,0,0,0,143,0,83,0,181,0,0,0,116,0,92,0,163,0,0,0,102,0,152,0,181,0,0,0,74,0,126,0,0,0,95,0,0,0,230,0,130,0,76,0,81,0,0,0,217,0,246,0,205,0,52,0,19,0,235,0,174,0,11,0,0,0,0,0,0,0,33,0,238,0,179,0,132,0,146,0,203,0,215,0,185,0,0,0,15,0,35,0,237,0,244,0,39,0,115,0,44,0,21,0,169,0,111,0,14,0,159,0,0,0,83,0,131,0,57,0,0,0,202,0,17,0,252,0,0,0,189,0,0,0,174,0,201,0,221,0,53,0,228,0,134,0,37,0,255,0,67,0,0,0,222,0,155,0,145,0,219,0,95,0,218,0,0,0,0,0,152,0,161,0,205,0,0,0,144,0,61,0,210,0,113,0,0,0,226,0,0,0,220,0,0,0,74,0,27,0,131,0,147,0,0,0,188,0,121,0,13,0,177,0,166,0,0,0,75,0,0,0,36,0,0,0,173,0,133,0,50,0,223,0,155,0,0,0,116,0,214,0,70,0,224,0,96,0,0,0,0,0,183,0,167,0,6,0,92,0,196,0,83,0,10,0,0,0,179,0,246,0,21,0,126,0,168,0,0,0,116,0,137,0,169,0,0,0,19,0,189,0,30,0,0,0,93,0,135,0,20,0,212,0,219,0,25,0,44,0,124,0,188,0,111,0,195,0,75,0,201,0,61,0,0,0,0,0,41,0,254,0,125,0,0,0,61,0,160,0,255,0,103,0,137,0,10,0,118,0,248,0,0,0,201,0,52,0,247,0,123,0,52,0,134,0,246,0,137,0,244,0,221,0,0,0,156,0,75,0,130,0,31,0,6,0,173,0,59,0,107,0,166,0,0,0,153,0,161,0,172,0,34,0,195,0,237,0,8,0,0,0,190,0,248,0,73,0,0,0,206,0,142,0,160,0,181,0,225,0,1,0,149,0,189,0,230,0,13,0,114,0,58,0,182,0,51,0,153,0,221,0,56,0,0,0,0,0,45,0,145,0,138,0,30,0,165,0,233,0,212,0,45,0,206,0,244,0,222,0,26,0,116,0,0,0,241,0,85,0,72,0,59,0,71,0,187,0,42,0,64,0,0,0,98,0,0,0,0,0,172,0,94,0,77,0,138,0,121,0,177,0,170,0,144,0,60,0,45,0,15,0,0,0,216,0,236,0,173,0,67,0,189,0,0,0,0,0,106,0,126,0,0,0,0,0,16,0,31,0,0,0,188,0,0,0,149,0,109,0,0,0,235,0,208,0,97,0,91,0,126,0,0,0,8,0,99,0,0,0,0,0,187,0,144,0,126,0,130,0,53,0,91,0,15,0,20,0,210,0,85,0,231,0,0,0,91,0,125,0,94,0,0,0,242,0,0,0,234,0,151,0,205,0,0,0,166,0,93,0,118,0,78,0,149,0,237,0,39,0,43,0,200,0,0,0,0,0,109,0,0,0,14,0,19,0,117,0,199,0,0,0,208,0,104,0,148,0,218,0,0,0,124,0,0,0,220,0,134,0,242,0,108,0,0,0,184,0,0,0,20,0,0,0,0,0,45,0,0,0,48,0,0,0,73,0,0,0,193,0,75,0,0,0,0,0,238,0,167,0,219,0,141,0,57,0,180,0,241,0,137,0,184,0,236,0,0,0,20,0,197,0,115,0,252,0,3,0,141,0,0,0,0,0,216,0,231,0,50,0,115,0,184,0,164,0);
signal scenario_full  : scenario_type := (0,0,17,31,225,31,225,30,162,31,162,30,162,29,240,31,192,31,207,31,207,30,207,29,93,31,134,31,218,31,41,31,41,30,41,29,49,31,235,31,243,31,90,31,109,31,57,31,57,30,225,31,232,31,185,31,72,31,223,31,69,31,150,31,61,31,61,31,226,31,125,31,53,31,255,31,97,31,82,31,174,31,50,31,132,31,89,31,117,31,117,30,204,31,194,31,27,31,179,31,229,31,60,31,253,31,60,31,180,31,180,30,207,31,105,31,229,31,229,30,43,31,31,31,192,31,134,31,134,30,187,31,9,31,49,31,64,31,246,31,233,31,162,31,113,31,113,30,150,31,150,30,241,31,127,31,203,31,72,31,254,31,66,31,149,31,160,31,251,31,62,31,224,31,195,31,187,31,10,31,252,31,79,31,194,31,51,31,51,30,23,31,170,31,7,31,224,31,224,30,230,31,230,30,233,31,233,30,65,31,169,31,137,31,137,30,60,31,60,30,162,31,188,31,188,30,131,31,195,31,8,31,42,31,58,31,181,31,234,31,173,31,213,31,213,30,89,31,94,31,76,31,81,31,204,31,224,31,205,31,205,30,51,31,51,30,226,31,177,31,139,31,56,31,198,31,205,31,25,31,114,31,122,31,215,31,215,30,215,29,54,31,21,31,238,31,238,30,143,31,177,31,201,31,38,31,151,31,180,31,180,30,122,31,213,31,90,31,90,30,162,31,219,31,219,30,2,31,43,31,129,31,29,31,89,31,94,31,140,31,34,31,254,31,254,30,156,31,30,31,30,30,122,31,11,31,11,30,11,29,11,28,133,31,173,31,143,31,67,31,51,31,222,31,212,31,196,31,12,31,12,30,187,31,239,31,105,31,105,30,55,31,55,30,119,31,119,30,132,31,249,31,104,31,104,30,203,31,48,31,18,31,125,31,186,31,185,31,185,30,53,31,53,30,252,31,252,30,255,31,255,30,143,31,117,31,214,31,66,31,66,30,66,29,66,28,30,31,63,31,8,31,8,30,171,31,171,30,171,29,212,31,57,31,80,31,80,30,158,31,37,31,199,31,216,31,112,31,244,31,244,30,165,31,160,31,117,31,203,31,237,31,71,31,241,31,58,31,93,31,35,31,165,31,110,31,110,30,110,29,172,31,96,31,96,30,96,29,170,31,43,31,239,31,146,31,196,31,8,31,127,31,127,30,125,31,128,31,128,30,252,31,174,31,252,31,104,31,104,30,104,29,143,31,83,31,181,31,181,30,116,31,92,31,163,31,163,30,102,31,152,31,181,31,181,30,74,31,126,31,126,30,95,31,95,30,230,31,130,31,76,31,81,31,81,30,217,31,246,31,205,31,52,31,19,31,235,31,174,31,11,31,11,30,11,29,11,28,33,31,238,31,179,31,132,31,146,31,203,31,215,31,185,31,185,30,15,31,35,31,237,31,244,31,39,31,115,31,44,31,21,31,169,31,111,31,14,31,159,31,159,30,83,31,131,31,57,31,57,30,202,31,17,31,252,31,252,30,189,31,189,30,174,31,201,31,221,31,53,31,228,31,134,31,37,31,255,31,67,31,67,30,222,31,155,31,145,31,219,31,95,31,218,31,218,30,218,29,152,31,161,31,205,31,205,30,144,31,61,31,210,31,113,31,113,30,226,31,226,30,220,31,220,30,74,31,27,31,131,31,147,31,147,30,188,31,121,31,13,31,177,31,166,31,166,30,75,31,75,30,36,31,36,30,173,31,133,31,50,31,223,31,155,31,155,30,116,31,214,31,70,31,224,31,96,31,96,30,96,29,183,31,167,31,6,31,92,31,196,31,83,31,10,31,10,30,179,31,246,31,21,31,126,31,168,31,168,30,116,31,137,31,169,31,169,30,19,31,189,31,30,31,30,30,93,31,135,31,20,31,212,31,219,31,25,31,44,31,124,31,188,31,111,31,195,31,75,31,201,31,61,31,61,30,61,29,41,31,254,31,125,31,125,30,61,31,160,31,255,31,103,31,137,31,10,31,118,31,248,31,248,30,201,31,52,31,247,31,123,31,52,31,134,31,246,31,137,31,244,31,221,31,221,30,156,31,75,31,130,31,31,31,6,31,173,31,59,31,107,31,166,31,166,30,153,31,161,31,172,31,34,31,195,31,237,31,8,31,8,30,190,31,248,31,73,31,73,30,206,31,142,31,160,31,181,31,225,31,1,31,149,31,189,31,230,31,13,31,114,31,58,31,182,31,51,31,153,31,221,31,56,31,56,30,56,29,45,31,145,31,138,31,30,31,165,31,233,31,212,31,45,31,206,31,244,31,222,31,26,31,116,31,116,30,241,31,85,31,72,31,59,31,71,31,187,31,42,31,64,31,64,30,98,31,98,30,98,29,172,31,94,31,77,31,138,31,121,31,177,31,170,31,144,31,60,31,45,31,15,31,15,30,216,31,236,31,173,31,67,31,189,31,189,30,189,29,106,31,126,31,126,30,126,29,16,31,31,31,31,30,188,31,188,30,149,31,109,31,109,30,235,31,208,31,97,31,91,31,126,31,126,30,8,31,99,31,99,30,99,29,187,31,144,31,126,31,130,31,53,31,91,31,15,31,20,31,210,31,85,31,231,31,231,30,91,31,125,31,94,31,94,30,242,31,242,30,234,31,151,31,205,31,205,30,166,31,93,31,118,31,78,31,149,31,237,31,39,31,43,31,200,31,200,30,200,29,109,31,109,30,14,31,19,31,117,31,199,31,199,30,208,31,104,31,148,31,218,31,218,30,124,31,124,30,220,31,134,31,242,31,108,31,108,30,184,31,184,30,20,31,20,30,20,29,45,31,45,30,48,31,48,30,73,31,73,30,193,31,75,31,75,30,75,29,238,31,167,31,219,31,141,31,57,31,180,31,241,31,137,31,184,31,236,31,236,30,20,31,197,31,115,31,252,31,3,31,141,31,141,30,141,29,216,31,231,31,50,31,115,31,184,31,164,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
