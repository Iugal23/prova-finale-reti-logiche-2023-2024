-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 888;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (160,0,0,0,0,0,0,0,140,0,104,0,0,0,131,0,125,0,218,0,0,0,134,0,73,0,0,0,225,0,189,0,61,0,0,0,9,0,207,0,0,0,11,0,83,0,91,0,176,0,78,0,80,0,16,0,246,0,0,0,252,0,120,0,234,0,15,0,107,0,149,0,42,0,0,0,0,0,123,0,224,0,0,0,140,0,0,0,215,0,208,0,220,0,48,0,114,0,127,0,30,0,96,0,0,0,0,0,180,0,194,0,57,0,198,0,115,0,163,0,35,0,144,0,78,0,147,0,62,0,149,0,45,0,95,0,0,0,174,0,0,0,161,0,255,0,133,0,179,0,73,0,153,0,0,0,166,0,124,0,6,0,36,0,26,0,56,0,0,0,0,0,36,0,156,0,155,0,118,0,78,0,235,0,224,0,116,0,196,0,0,0,0,0,79,0,4,0,0,0,199,0,88,0,187,0,0,0,13,0,170,0,0,0,47,0,31,0,98,0,0,0,0,0,37,0,148,0,28,0,216,0,238,0,41,0,177,0,99,0,0,0,13,0,0,0,207,0,225,0,247,0,54,0,204,0,16,0,0,0,153,0,13,0,112,0,81,0,234,0,114,0,2,0,43,0,84,0,177,0,205,0,153,0,0,0,31,0,238,0,0,0,216,0,14,0,94,0,0,0,0,0,107,0,0,0,10,0,223,0,80,0,250,0,81,0,132,0,0,0,0,0,196,0,53,0,0,0,139,0,0,0,129,0,90,0,54,0,84,0,141,0,0,0,137,0,110,0,60,0,189,0,106,0,0,0,0,0,1,0,162,0,0,0,32,0,152,0,79,0,56,0,87,0,216,0,165,0,0,0,0,0,88,0,201,0,84,0,20,0,192,0,187,0,232,0,24,0,112,0,28,0,192,0,165,0,181,0,71,0,105,0,244,0,0,0,230,0,181,0,40,0,242,0,74,0,0,0,114,0,0,0,0,0,155,0,173,0,90,0,132,0,59,0,0,0,171,0,40,0,0,0,30,0,202,0,162,0,192,0,227,0,0,0,172,0,0,0,114,0,71,0,254,0,206,0,0,0,0,0,100,0,79,0,60,0,222,0,106,0,166,0,71,0,79,0,2,0,183,0,4,0,85,0,0,0,254,0,190,0,224,0,0,0,39,0,166,0,109,0,78,0,125,0,22,0,5,0,69,0,51,0,104,0,171,0,189,0,87,0,160,0,86,0,0,0,101,0,21,0,0,0,77,0,103,0,15,0,70,0,187,0,151,0,101,0,111,0,0,0,138,0,226,0,162,0,125,0,1,0,156,0,123,0,170,0,0,0,0,0,0,0,5,0,9,0,106,0,189,0,134,0,150,0,103,0,182,0,59,0,148,0,113,0,81,0,0,0,3,0,64,0,218,0,151,0,54,0,220,0,42,0,176,0,35,0,78,0,71,0,210,0,233,0,111,0,214,0,196,0,67,0,156,0,244,0,181,0,179,0,213,0,0,0,248,0,115,0,247,0,1,0,122,0,111,0,186,0,0,0,32,0,0,0,54,0,98,0,237,0,130,0,115,0,253,0,0,0,0,0,4,0,177,0,0,0,0,0,0,0,0,0,72,0,244,0,97,0,0,0,0,0,15,0,0,0,177,0,68,0,23,0,0,0,78,0,0,0,0,0,48,0,71,0,0,0,117,0,188,0,121,0,119,0,102,0,229,0,0,0,229,0,20,0,0,0,150,0,191,0,45,0,160,0,237,0,208,0,0,0,245,0,0,0,123,0,0,0,0,0,165,0,0,0,0,0,17,0,236,0,192,0,175,0,209,0,0,0,142,0,35,0,250,0,203,0,44,0,196,0,83,0,110,0,140,0,0,0,204,0,0,0,148,0,5,0,147,0,83,0,204,0,77,0,241,0,214,0,97,0,48,0,175,0,245,0,148,0,95,0,123,0,0,0,102,0,0,0,171,0,223,0,209,0,118,0,148,0,232,0,219,0,162,0,180,0,162,0,147,0,166,0,179,0,0,0,140,0,27,0,153,0,11,0,156,0,0,0,0,0,45,0,10,0,170,0,224,0,211,0,181,0,0,0,228,0,0,0,0,0,202,0,145,0,43,0,94,0,237,0,103,0,116,0,24,0,145,0,145,0,71,0,132,0,193,0,0,0,6,0,0,0,96,0,116,0,126,0,103,0,234,0,245,0,137,0,0,0,220,0,68,0,235,0,57,0,35,0,0,0,86,0,168,0,229,0,99,0,45,0,125,0,218,0,0,0,135,0,111,0,0,0,167,0,54,0,0,0,147,0,253,0,0,0,0,0,250,0,124,0,42,0,0,0,223,0,171,0,123,0,0,0,111,0,189,0,16,0,198,0,78,0,211,0,0,0,0,0,207,0,192,0,0,0,135,0,0,0,246,0,208,0,36,0,0,0,86,0,100,0,0,0,92,0,217,0,137,0,66,0,198,0,190,0,233,0,66,0,0,0,78,0,0,0,7,0,212,0,214,0,106,0,88,0,186,0,19,0,130,0,181,0,146,0,0,0,134,0,174,0,55,0,139,0,19,0,73,0,0,0,244,0,185,0,0,0,189,0,0,0,110,0,0,0,156,0,141,0,118,0,0,0,44,0,142,0,84,0,0,0,123,0,195,0,0,0,228,0,34,0,172,0,194,0,0,0,100,0,218,0,114,0,216,0,157,0,20,0,254,0,23,0,182,0,233,0,248,0,0,0,6,0,0,0,54,0,28,0,102,0,64,0,0,0,12,0,0,0,164,0,69,0,40,0,237,0,20,0,13,0,4,0,0,0,231,0,126,0,219,0,232,0,255,0,58,0,90,0,181,0,0,0,106,0,107,0,113,0,0,0,62,0,0,0,48,0,173,0,158,0,0,0,206,0,232,0,162,0,249,0,0,0,18,0,18,0,0,0,59,0,0,0,92,0,0,0,218,0,139,0,162,0,0,0,220,0,219,0,242,0,80,0,0,0,221,0,195,0,43,0,0,0,95,0,245,0,31,0,10,0,218,0,0,0,65,0,15,0,0,0,18,0,0,0,80,0,0,0,141,0,88,0,231,0,65,0,119,0,126,0,188,0,253,0,0,0,175,0,215,0,97,0,0,0,59,0,204,0,0,0,0,0,19,0,69,0,0,0,0,0,31,0,0,0,0,0,53,0,41,0,240,0,0,0,87,0,71,0,0,0,203,0,210,0,199,0,29,0,109,0,100,0,239,0,55,0,236,0,191,0,204,0,184,0,89,0,105,0,45,0,99,0,22,0,52,0,92,0,119,0,2,0,8,0,82,0,0,0,0,0,5,0,5,0,183,0,230,0,79,0,93,0,226,0,100,0,48,0,159,0,210,0,128,0,122,0,155,0,0,0,0,0,71,0,0,0,224,0,178,0,14,0,0,0,0,0,99,0,0,0,252,0,81,0,251,0,48,0,0,0,0,0,171,0,200,0,176,0,191,0,197,0,57,0,27,0,183,0,21,0,137,0,167,0,54,0,14,0,44,0,152,0,160,0,57,0,49,0,20,0,193,0,0,0,111,0,131,0,0,0,14,0,5,0,29,0,147,0,122,0,199,0,70,0,217,0,198,0,178,0,0,0,245,0,232,0,29,0,206,0,7,0,147,0,186,0,51,0,129,0,0,0,153,0,179,0,102,0,90,0,0,0,45,0,78,0,143,0,176,0,154,0,111,0,200,0,7,0,0,0,107,0,70,0,0,0,248,0,148,0,144,0,149,0,254,0,0,0,179,0,64,0,137,0,63,0,190,0,116,0,0,0,177,0,72,0,160,0,46,0,145,0,57,0,16,0,176,0,0,0,73,0,208,0,0,0,98,0,229,0,152,0,60,0,0,0,0,0,152,0,146,0,0,0,0,0,100,0,197,0,78,0,45,0,186,0,136,0,131,0,31,0,243,0,0,0,24,0,199,0,224,0,66,0,38,0,0,0,67,0,99,0,0,0,222,0,5,0,233,0,164,0,45,0,0,0);
signal scenario_full  : scenario_type := (160,31,160,30,160,29,160,28,140,31,104,31,104,30,131,31,125,31,218,31,218,30,134,31,73,31,73,30,225,31,189,31,61,31,61,30,9,31,207,31,207,30,11,31,83,31,91,31,176,31,78,31,80,31,16,31,246,31,246,30,252,31,120,31,234,31,15,31,107,31,149,31,42,31,42,30,42,29,123,31,224,31,224,30,140,31,140,30,215,31,208,31,220,31,48,31,114,31,127,31,30,31,96,31,96,30,96,29,180,31,194,31,57,31,198,31,115,31,163,31,35,31,144,31,78,31,147,31,62,31,149,31,45,31,95,31,95,30,174,31,174,30,161,31,255,31,133,31,179,31,73,31,153,31,153,30,166,31,124,31,6,31,36,31,26,31,56,31,56,30,56,29,36,31,156,31,155,31,118,31,78,31,235,31,224,31,116,31,196,31,196,30,196,29,79,31,4,31,4,30,199,31,88,31,187,31,187,30,13,31,170,31,170,30,47,31,31,31,98,31,98,30,98,29,37,31,148,31,28,31,216,31,238,31,41,31,177,31,99,31,99,30,13,31,13,30,207,31,225,31,247,31,54,31,204,31,16,31,16,30,153,31,13,31,112,31,81,31,234,31,114,31,2,31,43,31,84,31,177,31,205,31,153,31,153,30,31,31,238,31,238,30,216,31,14,31,94,31,94,30,94,29,107,31,107,30,10,31,223,31,80,31,250,31,81,31,132,31,132,30,132,29,196,31,53,31,53,30,139,31,139,30,129,31,90,31,54,31,84,31,141,31,141,30,137,31,110,31,60,31,189,31,106,31,106,30,106,29,1,31,162,31,162,30,32,31,152,31,79,31,56,31,87,31,216,31,165,31,165,30,165,29,88,31,201,31,84,31,20,31,192,31,187,31,232,31,24,31,112,31,28,31,192,31,165,31,181,31,71,31,105,31,244,31,244,30,230,31,181,31,40,31,242,31,74,31,74,30,114,31,114,30,114,29,155,31,173,31,90,31,132,31,59,31,59,30,171,31,40,31,40,30,30,31,202,31,162,31,192,31,227,31,227,30,172,31,172,30,114,31,71,31,254,31,206,31,206,30,206,29,100,31,79,31,60,31,222,31,106,31,166,31,71,31,79,31,2,31,183,31,4,31,85,31,85,30,254,31,190,31,224,31,224,30,39,31,166,31,109,31,78,31,125,31,22,31,5,31,69,31,51,31,104,31,171,31,189,31,87,31,160,31,86,31,86,30,101,31,21,31,21,30,77,31,103,31,15,31,70,31,187,31,151,31,101,31,111,31,111,30,138,31,226,31,162,31,125,31,1,31,156,31,123,31,170,31,170,30,170,29,170,28,5,31,9,31,106,31,189,31,134,31,150,31,103,31,182,31,59,31,148,31,113,31,81,31,81,30,3,31,64,31,218,31,151,31,54,31,220,31,42,31,176,31,35,31,78,31,71,31,210,31,233,31,111,31,214,31,196,31,67,31,156,31,244,31,181,31,179,31,213,31,213,30,248,31,115,31,247,31,1,31,122,31,111,31,186,31,186,30,32,31,32,30,54,31,98,31,237,31,130,31,115,31,253,31,253,30,253,29,4,31,177,31,177,30,177,29,177,28,177,27,72,31,244,31,97,31,97,30,97,29,15,31,15,30,177,31,68,31,23,31,23,30,78,31,78,30,78,29,48,31,71,31,71,30,117,31,188,31,121,31,119,31,102,31,229,31,229,30,229,31,20,31,20,30,150,31,191,31,45,31,160,31,237,31,208,31,208,30,245,31,245,30,123,31,123,30,123,29,165,31,165,30,165,29,17,31,236,31,192,31,175,31,209,31,209,30,142,31,35,31,250,31,203,31,44,31,196,31,83,31,110,31,140,31,140,30,204,31,204,30,148,31,5,31,147,31,83,31,204,31,77,31,241,31,214,31,97,31,48,31,175,31,245,31,148,31,95,31,123,31,123,30,102,31,102,30,171,31,223,31,209,31,118,31,148,31,232,31,219,31,162,31,180,31,162,31,147,31,166,31,179,31,179,30,140,31,27,31,153,31,11,31,156,31,156,30,156,29,45,31,10,31,170,31,224,31,211,31,181,31,181,30,228,31,228,30,228,29,202,31,145,31,43,31,94,31,237,31,103,31,116,31,24,31,145,31,145,31,71,31,132,31,193,31,193,30,6,31,6,30,96,31,116,31,126,31,103,31,234,31,245,31,137,31,137,30,220,31,68,31,235,31,57,31,35,31,35,30,86,31,168,31,229,31,99,31,45,31,125,31,218,31,218,30,135,31,111,31,111,30,167,31,54,31,54,30,147,31,253,31,253,30,253,29,250,31,124,31,42,31,42,30,223,31,171,31,123,31,123,30,111,31,189,31,16,31,198,31,78,31,211,31,211,30,211,29,207,31,192,31,192,30,135,31,135,30,246,31,208,31,36,31,36,30,86,31,100,31,100,30,92,31,217,31,137,31,66,31,198,31,190,31,233,31,66,31,66,30,78,31,78,30,7,31,212,31,214,31,106,31,88,31,186,31,19,31,130,31,181,31,146,31,146,30,134,31,174,31,55,31,139,31,19,31,73,31,73,30,244,31,185,31,185,30,189,31,189,30,110,31,110,30,156,31,141,31,118,31,118,30,44,31,142,31,84,31,84,30,123,31,195,31,195,30,228,31,34,31,172,31,194,31,194,30,100,31,218,31,114,31,216,31,157,31,20,31,254,31,23,31,182,31,233,31,248,31,248,30,6,31,6,30,54,31,28,31,102,31,64,31,64,30,12,31,12,30,164,31,69,31,40,31,237,31,20,31,13,31,4,31,4,30,231,31,126,31,219,31,232,31,255,31,58,31,90,31,181,31,181,30,106,31,107,31,113,31,113,30,62,31,62,30,48,31,173,31,158,31,158,30,206,31,232,31,162,31,249,31,249,30,18,31,18,31,18,30,59,31,59,30,92,31,92,30,218,31,139,31,162,31,162,30,220,31,219,31,242,31,80,31,80,30,221,31,195,31,43,31,43,30,95,31,245,31,31,31,10,31,218,31,218,30,65,31,15,31,15,30,18,31,18,30,80,31,80,30,141,31,88,31,231,31,65,31,119,31,126,31,188,31,253,31,253,30,175,31,215,31,97,31,97,30,59,31,204,31,204,30,204,29,19,31,69,31,69,30,69,29,31,31,31,30,31,29,53,31,41,31,240,31,240,30,87,31,71,31,71,30,203,31,210,31,199,31,29,31,109,31,100,31,239,31,55,31,236,31,191,31,204,31,184,31,89,31,105,31,45,31,99,31,22,31,52,31,92,31,119,31,2,31,8,31,82,31,82,30,82,29,5,31,5,31,183,31,230,31,79,31,93,31,226,31,100,31,48,31,159,31,210,31,128,31,122,31,155,31,155,30,155,29,71,31,71,30,224,31,178,31,14,31,14,30,14,29,99,31,99,30,252,31,81,31,251,31,48,31,48,30,48,29,171,31,200,31,176,31,191,31,197,31,57,31,27,31,183,31,21,31,137,31,167,31,54,31,14,31,44,31,152,31,160,31,57,31,49,31,20,31,193,31,193,30,111,31,131,31,131,30,14,31,5,31,29,31,147,31,122,31,199,31,70,31,217,31,198,31,178,31,178,30,245,31,232,31,29,31,206,31,7,31,147,31,186,31,51,31,129,31,129,30,153,31,179,31,102,31,90,31,90,30,45,31,78,31,143,31,176,31,154,31,111,31,200,31,7,31,7,30,107,31,70,31,70,30,248,31,148,31,144,31,149,31,254,31,254,30,179,31,64,31,137,31,63,31,190,31,116,31,116,30,177,31,72,31,160,31,46,31,145,31,57,31,16,31,176,31,176,30,73,31,208,31,208,30,98,31,229,31,152,31,60,31,60,30,60,29,152,31,146,31,146,30,146,29,100,31,197,31,78,31,45,31,186,31,136,31,131,31,31,31,243,31,243,30,24,31,199,31,224,31,66,31,38,31,38,30,67,31,99,31,99,30,222,31,5,31,233,31,164,31,45,31,45,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
