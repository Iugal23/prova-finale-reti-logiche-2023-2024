-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 921;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (180,0,131,0,194,0,95,0,199,0,8,0,9,0,186,0,210,0,213,0,72,0,144,0,37,0,85,0,200,0,213,0,0,0,64,0,0,0,223,0,222,0,153,0,244,0,33,0,81,0,146,0,231,0,250,0,65,0,0,0,241,0,227,0,203,0,20,0,0,0,0,0,99,0,126,0,40,0,241,0,186,0,33,0,0,0,114,0,216,0,190,0,122,0,254,0,0,0,76,0,123,0,86,0,0,0,0,0,110,0,132,0,58,0,174,0,131,0,34,0,233,0,0,0,220,0,164,0,0,0,231,0,237,0,157,0,40,0,0,0,51,0,151,0,0,0,144,0,0,0,36,0,227,0,0,0,246,0,105,0,236,0,95,0,54,0,63,0,85,0,26,0,127,0,152,0,0,0,149,0,40,0,0,0,210,0,207,0,196,0,84,0,187,0,55,0,52,0,241,0,23,0,0,0,206,0,203,0,92,0,72,0,126,0,116,0,210,0,253,0,122,0,0,0,193,0,103,0,102,0,192,0,212,0,4,0,20,0,171,0,12,0,177,0,0,0,35,0,0,0,230,0,0,0,209,0,54,0,70,0,100,0,221,0,159,0,226,0,203,0,91,0,0,0,106,0,0,0,30,0,145,0,0,0,216,0,173,0,73,0,0,0,102,0,0,0,228,0,228,0,0,0,120,0,97,0,222,0,0,0,130,0,95,0,0,0,47,0,146,0,0,0,60,0,178,0,75,0,0,0,0,0,93,0,127,0,254,0,13,0,0,0,130,0,20,0,0,0,0,0,196,0,10,0,0,0,69,0,190,0,16,0,17,0,30,0,3,0,138,0,0,0,229,0,0,0,134,0,6,0,206,0,228,0,211,0,10,0,0,0,99,0,92,0,121,0,188,0,218,0,0,0,22,0,236,0,0,0,155,0,105,0,74,0,35,0,144,0,0,0,0,0,121,0,48,0,249,0,134,0,218,0,195,0,77,0,235,0,0,0,165,0,157,0,240,0,128,0,90,0,218,0,0,0,218,0,0,0,52,0,83,0,0,0,153,0,255,0,243,0,142,0,222,0,67,0,44,0,63,0,236,0,0,0,5,0,185,0,197,0,173,0,0,0,52,0,87,0,44,0,205,0,18,0,0,0,155,0,0,0,185,0,203,0,127,0,172,0,55,0,178,0,0,0,66,0,110,0,234,0,0,0,226,0,205,0,0,0,0,0,83,0,74,0,0,0,216,0,87,0,0,0,22,0,1,0,224,0,129,0,242,0,190,0,163,0,249,0,21,0,0,0,32,0,26,0,156,0,0,0,0,0,183,0,0,0,0,0,180,0,153,0,167,0,2,0,172,0,0,0,0,0,9,0,0,0,109,0,105,0,0,0,0,0,35,0,184,0,147,0,7,0,30,0,47,0,102,0,0,0,158,0,240,0,201,0,84,0,7,0,0,0,7,0,142,0,147,0,163,0,72,0,216,0,28,0,48,0,0,0,156,0,0,0,209,0,135,0,35,0,102,0,154,0,0,0,40,0,0,0,0,0,216,0,58,0,47,0,236,0,0,0,78,0,34,0,0,0,145,0,126,0,60,0,60,0,0,0,0,0,0,0,23,0,113,0,213,0,132,0,0,0,210,0,0,0,187,0,198,0,140,0,171,0,0,0,194,0,175,0,0,0,26,0,111,0,19,0,208,0,0,0,19,0,39,0,0,0,100,0,235,0,144,0,234,0,253,0,238,0,16,0,176,0,0,0,49,0,200,0,5,0,27,0,144,0,0,0,74,0,50,0,246,0,191,0,237,0,73,0,12,0,152,0,245,0,0,0,40,0,159,0,93,0,61,0,221,0,143,0,60,0,212,0,90,0,0,0,176,0,66,0,38,0,201,0,129,0,205,0,0,0,239,0,119,0,143,0,112,0,247,0,0,0,149,0,50,0,120,0,225,0,0,0,172,0,0,0,0,0,238,0,126,0,144,0,240,0,71,0,157,0,150,0,97,0,83,0,33,0,230,0,68,0,84,0,42,0,40,0,193,0,0,0,132,0,216,0,93,0,239,0,254,0,168,0,104,0,215,0,119,0,119,0,163,0,0,0,136,0,27,0,137,0,46,0,20,0,133,0,0,0,63,0,68,0,127,0,0,0,0,0,13,0,167,0,132,0,77,0,215,0,0,0,0,0,246,0,139,0,72,0,230,0,135,0,94,0,116,0,119,0,226,0,147,0,220,0,0,0,0,0,0,0,95,0,0,0,81,0,200,0,0,0,187,0,0,0,219,0,0,0,70,0,54,0,135,0,0,0,0,0,24,0,155,0,52,0,3,0,133,0,84,0,205,0,0,0,0,0,184,0,61,0,98,0,90,0,53,0,63,0,253,0,0,0,0,0,102,0,42,0,194,0,239,0,0,0,78,0,0,0,50,0,182,0,240,0,134,0,166,0,0,0,225,0,48,0,36,0,194,0,0,0,10,0,186,0,217,0,49,0,0,0,25,0,178,0,253,0,17,0,190,0,125,0,222,0,157,0,2,0,92,0,212,0,65,0,130,0,71,0,44,0,171,0,47,0,230,0,15,0,52,0,48,0,182,0,224,0,252,0,130,0,0,0,183,0,0,0,131,0,0,0,72,0,42,0,160,0,127,0,0,0,31,0,75,0,97,0,4,0,138,0,84,0,38,0,0,0,32,0,145,0,75,0,105,0,80,0,98,0,225,0,181,0,0,0,0,0,62,0,142,0,34,0,0,0,2,0,83,0,238,0,0,0,240,0,213,0,51,0,100,0,114,0,192,0,98,0,232,0,107,0,27,0,172,0,0,0,207,0,91,0,124,0,73,0,0,0,29,0,231,0,31,0,221,0,152,0,0,0,71,0,64,0,213,0,174,0,0,0,72,0,186,0,0,0,239,0,161,0,43,0,208,0,204,0,111,0,41,0,229,0,0,0,233,0,175,0,0,0,81,0,0,0,36,0,20,0,0,0,82,0,0,0,144,0,0,0,0,0,244,0,35,0,59,0,77,0,152,0,216,0,167,0,27,0,105,0,142,0,0,0,0,0,0,0,0,0,213,0,226,0,24,0,21,0,0,0,129,0,211,0,114,0,171,0,21,0,7,0,158,0,0,0,0,0,196,0,179,0,211,0,133,0,0,0,4,0,91,0,0,0,198,0,181,0,13,0,0,0,39,0,123,0,18,0,0,0,213,0,135,0,119,0,163,0,0,0,110,0,170,0,153,0,79,0,237,0,23,0,99,0,166,0,0,0,124,0,160,0,116,0,42,0,122,0,39,0,35,0,219,0,160,0,49,0,152,0,147,0,91,0,84,0,29,0,0,0,24,0,53,0,168,0,36,0,39,0,156,0,242,0,152,0,83,0,6,0,87,0,185,0,74,0,163,0,130,0,0,0,253,0,244,0,211,0,206,0,102,0,0,0,69,0,210,0,0,0,137,0,61,0,122,0,243,0,213,0,0,0,162,0,22,0,90,0,228,0,191,0,8,0,131,0,0,0,0,0,50,0,217,0,181,0,148,0,205,0,135,0,154,0,79,0,179,0,136,0,84,0,109,0,0,0,38,0,121,0,43,0,0,0,0,0,248,0,169,0,0,0,163,0,230,0,92,0,245,0,0,0,177,0,86,0,133,0,231,0,117,0,231,0,175,0,0,0,109,0,218,0,175,0,200,0,51,0,90,0,94,0,88,0,173,0,45,0,0,0,74,0,0,0,0,0,0,0,41,0,0,0,138,0,0,0,2,0,173,0,222,0,218,0,0,0,0,0,175,0,212,0,0,0,175,0,47,0,0,0,135,0,193,0,0,0,0,0,249,0,153,0,192,0,132,0,173,0,128,0,82,0,66,0,0,0,0,0,250,0,0,0,10,0,0,0,0,0,14,0,165,0,94,0,205,0,170,0,177,0,183,0,152,0,188,0,197,0,0,0,194,0,0,0,201,0,225,0,125,0,145,0,238,0,251,0,0,0,0,0,0,0,72,0,19,0,122,0,85,0,0,0,157,0,117,0,237,0,0,0,123,0,0,0,0,0,155,0,0,0,86,0,194,0,246,0,176,0,0,0,87,0,0,0,167,0,204,0,95,0,241,0,188,0,75,0,98,0,200,0,92,0,227,0,119,0,36,0,253,0,206,0);
signal scenario_full  : scenario_type := (180,31,131,31,194,31,95,31,199,31,8,31,9,31,186,31,210,31,213,31,72,31,144,31,37,31,85,31,200,31,213,31,213,30,64,31,64,30,223,31,222,31,153,31,244,31,33,31,81,31,146,31,231,31,250,31,65,31,65,30,241,31,227,31,203,31,20,31,20,30,20,29,99,31,126,31,40,31,241,31,186,31,33,31,33,30,114,31,216,31,190,31,122,31,254,31,254,30,76,31,123,31,86,31,86,30,86,29,110,31,132,31,58,31,174,31,131,31,34,31,233,31,233,30,220,31,164,31,164,30,231,31,237,31,157,31,40,31,40,30,51,31,151,31,151,30,144,31,144,30,36,31,227,31,227,30,246,31,105,31,236,31,95,31,54,31,63,31,85,31,26,31,127,31,152,31,152,30,149,31,40,31,40,30,210,31,207,31,196,31,84,31,187,31,55,31,52,31,241,31,23,31,23,30,206,31,203,31,92,31,72,31,126,31,116,31,210,31,253,31,122,31,122,30,193,31,103,31,102,31,192,31,212,31,4,31,20,31,171,31,12,31,177,31,177,30,35,31,35,30,230,31,230,30,209,31,54,31,70,31,100,31,221,31,159,31,226,31,203,31,91,31,91,30,106,31,106,30,30,31,145,31,145,30,216,31,173,31,73,31,73,30,102,31,102,30,228,31,228,31,228,30,120,31,97,31,222,31,222,30,130,31,95,31,95,30,47,31,146,31,146,30,60,31,178,31,75,31,75,30,75,29,93,31,127,31,254,31,13,31,13,30,130,31,20,31,20,30,20,29,196,31,10,31,10,30,69,31,190,31,16,31,17,31,30,31,3,31,138,31,138,30,229,31,229,30,134,31,6,31,206,31,228,31,211,31,10,31,10,30,99,31,92,31,121,31,188,31,218,31,218,30,22,31,236,31,236,30,155,31,105,31,74,31,35,31,144,31,144,30,144,29,121,31,48,31,249,31,134,31,218,31,195,31,77,31,235,31,235,30,165,31,157,31,240,31,128,31,90,31,218,31,218,30,218,31,218,30,52,31,83,31,83,30,153,31,255,31,243,31,142,31,222,31,67,31,44,31,63,31,236,31,236,30,5,31,185,31,197,31,173,31,173,30,52,31,87,31,44,31,205,31,18,31,18,30,155,31,155,30,185,31,203,31,127,31,172,31,55,31,178,31,178,30,66,31,110,31,234,31,234,30,226,31,205,31,205,30,205,29,83,31,74,31,74,30,216,31,87,31,87,30,22,31,1,31,224,31,129,31,242,31,190,31,163,31,249,31,21,31,21,30,32,31,26,31,156,31,156,30,156,29,183,31,183,30,183,29,180,31,153,31,167,31,2,31,172,31,172,30,172,29,9,31,9,30,109,31,105,31,105,30,105,29,35,31,184,31,147,31,7,31,30,31,47,31,102,31,102,30,158,31,240,31,201,31,84,31,7,31,7,30,7,31,142,31,147,31,163,31,72,31,216,31,28,31,48,31,48,30,156,31,156,30,209,31,135,31,35,31,102,31,154,31,154,30,40,31,40,30,40,29,216,31,58,31,47,31,236,31,236,30,78,31,34,31,34,30,145,31,126,31,60,31,60,31,60,30,60,29,60,28,23,31,113,31,213,31,132,31,132,30,210,31,210,30,187,31,198,31,140,31,171,31,171,30,194,31,175,31,175,30,26,31,111,31,19,31,208,31,208,30,19,31,39,31,39,30,100,31,235,31,144,31,234,31,253,31,238,31,16,31,176,31,176,30,49,31,200,31,5,31,27,31,144,31,144,30,74,31,50,31,246,31,191,31,237,31,73,31,12,31,152,31,245,31,245,30,40,31,159,31,93,31,61,31,221,31,143,31,60,31,212,31,90,31,90,30,176,31,66,31,38,31,201,31,129,31,205,31,205,30,239,31,119,31,143,31,112,31,247,31,247,30,149,31,50,31,120,31,225,31,225,30,172,31,172,30,172,29,238,31,126,31,144,31,240,31,71,31,157,31,150,31,97,31,83,31,33,31,230,31,68,31,84,31,42,31,40,31,193,31,193,30,132,31,216,31,93,31,239,31,254,31,168,31,104,31,215,31,119,31,119,31,163,31,163,30,136,31,27,31,137,31,46,31,20,31,133,31,133,30,63,31,68,31,127,31,127,30,127,29,13,31,167,31,132,31,77,31,215,31,215,30,215,29,246,31,139,31,72,31,230,31,135,31,94,31,116,31,119,31,226,31,147,31,220,31,220,30,220,29,220,28,95,31,95,30,81,31,200,31,200,30,187,31,187,30,219,31,219,30,70,31,54,31,135,31,135,30,135,29,24,31,155,31,52,31,3,31,133,31,84,31,205,31,205,30,205,29,184,31,61,31,98,31,90,31,53,31,63,31,253,31,253,30,253,29,102,31,42,31,194,31,239,31,239,30,78,31,78,30,50,31,182,31,240,31,134,31,166,31,166,30,225,31,48,31,36,31,194,31,194,30,10,31,186,31,217,31,49,31,49,30,25,31,178,31,253,31,17,31,190,31,125,31,222,31,157,31,2,31,92,31,212,31,65,31,130,31,71,31,44,31,171,31,47,31,230,31,15,31,52,31,48,31,182,31,224,31,252,31,130,31,130,30,183,31,183,30,131,31,131,30,72,31,42,31,160,31,127,31,127,30,31,31,75,31,97,31,4,31,138,31,84,31,38,31,38,30,32,31,145,31,75,31,105,31,80,31,98,31,225,31,181,31,181,30,181,29,62,31,142,31,34,31,34,30,2,31,83,31,238,31,238,30,240,31,213,31,51,31,100,31,114,31,192,31,98,31,232,31,107,31,27,31,172,31,172,30,207,31,91,31,124,31,73,31,73,30,29,31,231,31,31,31,221,31,152,31,152,30,71,31,64,31,213,31,174,31,174,30,72,31,186,31,186,30,239,31,161,31,43,31,208,31,204,31,111,31,41,31,229,31,229,30,233,31,175,31,175,30,81,31,81,30,36,31,20,31,20,30,82,31,82,30,144,31,144,30,144,29,244,31,35,31,59,31,77,31,152,31,216,31,167,31,27,31,105,31,142,31,142,30,142,29,142,28,142,27,213,31,226,31,24,31,21,31,21,30,129,31,211,31,114,31,171,31,21,31,7,31,158,31,158,30,158,29,196,31,179,31,211,31,133,31,133,30,4,31,91,31,91,30,198,31,181,31,13,31,13,30,39,31,123,31,18,31,18,30,213,31,135,31,119,31,163,31,163,30,110,31,170,31,153,31,79,31,237,31,23,31,99,31,166,31,166,30,124,31,160,31,116,31,42,31,122,31,39,31,35,31,219,31,160,31,49,31,152,31,147,31,91,31,84,31,29,31,29,30,24,31,53,31,168,31,36,31,39,31,156,31,242,31,152,31,83,31,6,31,87,31,185,31,74,31,163,31,130,31,130,30,253,31,244,31,211,31,206,31,102,31,102,30,69,31,210,31,210,30,137,31,61,31,122,31,243,31,213,31,213,30,162,31,22,31,90,31,228,31,191,31,8,31,131,31,131,30,131,29,50,31,217,31,181,31,148,31,205,31,135,31,154,31,79,31,179,31,136,31,84,31,109,31,109,30,38,31,121,31,43,31,43,30,43,29,248,31,169,31,169,30,163,31,230,31,92,31,245,31,245,30,177,31,86,31,133,31,231,31,117,31,231,31,175,31,175,30,109,31,218,31,175,31,200,31,51,31,90,31,94,31,88,31,173,31,45,31,45,30,74,31,74,30,74,29,74,28,41,31,41,30,138,31,138,30,2,31,173,31,222,31,218,31,218,30,218,29,175,31,212,31,212,30,175,31,47,31,47,30,135,31,193,31,193,30,193,29,249,31,153,31,192,31,132,31,173,31,128,31,82,31,66,31,66,30,66,29,250,31,250,30,10,31,10,30,10,29,14,31,165,31,94,31,205,31,170,31,177,31,183,31,152,31,188,31,197,31,197,30,194,31,194,30,201,31,225,31,125,31,145,31,238,31,251,31,251,30,251,29,251,28,72,31,19,31,122,31,85,31,85,30,157,31,117,31,237,31,237,30,123,31,123,30,123,29,155,31,155,30,86,31,194,31,246,31,176,31,176,30,87,31,87,30,167,31,204,31,95,31,241,31,188,31,75,31,98,31,200,31,92,31,227,31,119,31,36,31,253,31,206,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
