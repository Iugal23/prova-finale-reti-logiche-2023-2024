-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 912;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,198,0,242,0,180,0,0,0,111,0,68,0,103,0,251,0,163,0,234,0,21,0,223,0,154,0,0,0,15,0,147,0,128,0,0,0,102,0,243,0,37,0,74,0,27,0,0,0,58,0,197,0,222,0,151,0,218,0,149,0,68,0,144,0,185,0,227,0,190,0,188,0,131,0,188,0,254,0,194,0,70,0,10,0,0,0,196,0,231,0,0,0,163,0,12,0,0,0,119,0,86,0,0,0,64,0,216,0,126,0,217,0,2,0,0,0,0,0,0,0,8,0,48,0,20,0,92,0,97,0,99,0,0,0,21,0,86,0,198,0,0,0,16,0,234,0,18,0,5,0,0,0,220,0,152,0,244,0,36,0,227,0,230,0,225,0,0,0,15,0,86,0,0,0,252,0,26,0,2,0,240,0,149,0,110,0,241,0,233,0,20,0,0,0,237,0,52,0,31,0,240,0,0,0,0,0,93,0,12,0,25,0,153,0,186,0,214,0,185,0,0,0,147,0,111,0,0,0,120,0,212,0,161,0,201,0,74,0,228,0,208,0,0,0,91,0,180,0,116,0,234,0,101,0,80,0,0,0,19,0,0,0,36,0,136,0,13,0,187,0,17,0,0,0,0,0,167,0,0,0,210,0,113,0,73,0,83,0,228,0,0,0,90,0,57,0,187,0,234,0,107,0,220,0,133,0,118,0,81,0,103,0,61,0,96,0,2,0,226,0,68,0,17,0,28,0,0,0,104,0,200,0,49,0,184,0,103,0,155,0,64,0,8,0,111,0,43,0,114,0,195,0,251,0,225,0,254,0,119,0,38,0,3,0,15,0,85,0,124,0,132,0,142,0,207,0,14,0,111,0,224,0,168,0,0,0,236,0,250,0,195,0,138,0,164,0,0,0,157,0,212,0,10,0,194,0,146,0,182,0,151,0,166,0,19,0,129,0,139,0,116,0,61,0,59,0,240,0,123,0,0,0,72,0,177,0,59,0,44,0,0,0,37,0,34,0,145,0,237,0,0,0,27,0,0,0,138,0,109,0,31,0,133,0,68,0,95,0,0,0,0,0,0,0,0,0,176,0,167,0,96,0,165,0,165,0,40,0,199,0,187,0,150,0,201,0,112,0,186,0,85,0,0,0,21,0,40,0,99,0,149,0,51,0,48,0,0,0,14,0,211,0,12,0,207,0,56,0,131,0,72,0,253,0,127,0,0,0,0,0,0,0,7,0,53,0,201,0,91,0,0,0,0,0,0,0,189,0,64,0,242,0,253,0,0,0,72,0,9,0,43,0,184,0,89,0,15,0,32,0,185,0,132,0,252,0,21,0,70,0,142,0,0,0,128,0,5,0,0,0,28,0,16,0,215,0,163,0,253,0,92,0,115,0,234,0,0,0,90,0,140,0,217,0,224,0,150,0,155,0,128,0,61,0,148,0,160,0,188,0,135,0,16,0,99,0,89,0,94,0,242,0,151,0,205,0,121,0,162,0,211,0,183,0,187,0,240,0,239,0,216,0,134,0,146,0,0,0,132,0,113,0,72,0,250,0,187,0,144,0,203,0,83,0,62,0,54,0,224,0,39,0,29,0,0,0,199,0,251,0,0,0,101,0,237,0,150,0,210,0,93,0,46,0,83,0,41,0,208,0,70,0,248,0,180,0,115,0,89,0,102,0,33,0,141,0,14,0,73,0,19,0,5,0,89,0,174,0,211,0,183,0,84,0,0,0,177,0,0,0,11,0,0,0,0,0,70,0,180,0,148,0,242,0,140,0,27,0,155,0,255,0,51,0,0,0,30,0,4,0,64,0,214,0,83,0,29,0,110,0,9,0,24,0,108,0,242,0,171,0,123,0,0,0,129,0,58,0,157,0,149,0,249,0,115,0,9,0,70,0,104,0,0,0,64,0,16,0,103,0,0,0,1,0,53,0,47,0,121,0,231,0,181,0,54,0,5,0,83,0,134,0,168,0,117,0,236,0,199,0,235,0,196,0,109,0,42,0,0,0,240,0,1,0,51,0,163,0,0,0,233,0,191,0,146,0,29,0,221,0,0,0,215,0,164,0,212,0,238,0,91,0,0,0,65,0,0,0,21,0,94,0,213,0,187,0,195,0,182,0,0,0,200,0,232,0,143,0,0,0,247,0,136,0,0,0,0,0,0,0,243,0,43,0,7,0,0,0,72,0,83,0,111,0,16,0,209,0,149,0,141,0,7,0,28,0,0,0,94,0,0,0,0,0,53,0,0,0,83,0,252,0,231,0,247,0,31,0,4,0,243,0,0,0,239,0,0,0,78,0,0,0,16,0,0,0,32,0,87,0,61,0,69,0,181,0,0,0,101,0,200,0,0,0,158,0,179,0,116,0,0,0,137,0,133,0,0,0,140,0,186,0,217,0,131,0,88,0,121,0,111,0,11,0,146,0,214,0,255,0,151,0,0,0,0,0,30,0,60,0,0,0,0,0,0,0,113,0,254,0,167,0,0,0,171,0,105,0,156,0,243,0,0,0,0,0,54,0,130,0,23,0,227,0,215,0,190,0,172,0,153,0,8,0,44,0,231,0,38,0,0,0,224,0,57,0,29,0,99,0,108,0,0,0,121,0,90,0,0,0,89,0,233,0,254,0,222,0,185,0,94,0,241,0,0,0,148,0,82,0,84,0,70,0,71,0,0,0,231,0,18,0,70,0,89,0,225,0,7,0,106,0,0,0,237,0,195,0,103,0,0,0,27,0,131,0,137,0,246,0,198,0,121,0,0,0,0,0,0,0,216,0,202,0,0,0,36,0,187,0,191,0,224,0,215,0,85,0,0,0,209,0,53,0,204,0,182,0,255,0,31,0,2,0,83,0,254,0,0,0,172,0,177,0,138,0,195,0,0,0,121,0,133,0,89,0,165,0,140,0,212,0,0,0,192,0,178,0,0,0,222,0,142,0,98,0,40,0,93,0,89,0,186,0,128,0,134,0,100,0,93,0,246,0,0,0,0,0,45,0,98,0,31,0,190,0,252,0,58,0,156,0,94,0,208,0,0,0,0,0,137,0,0,0,173,0,0,0,203,0,68,0,127,0,0,0,83,0,194,0,245,0,175,0,227,0,202,0,176,0,67,0,3,0,243,0,22,0,187,0,227,0,0,0,146,0,154,0,170,0,95,0,84,0,0,0,212,0,240,0,156,0,235,0,0,0,106,0,164,0,209,0,112,0,4,0,206,0,128,0,246,0,126,0,201,0,75,0,0,0,98,0,211,0,247,0,176,0,114,0,0,0,87,0,67,0,153,0,191,0,107,0,34,0,0,0,0,0,0,0,0,0,0,0,30,0,64,0,27,0,130,0,71,0,0,0,0,0,174,0,61,0,81,0,66,0,0,0,7,0,0,0,176,0,204,0,119,0,0,0,0,0,186,0,0,0,137,0,179,0,37,0,0,0,80,0,184,0,0,0,157,0,25,0,192,0,250,0,0,0,36,0,22,0,0,0,0,0,56,0,0,0,121,0,0,0,0,0,74,0,0,0,199,0,0,0,119,0,172,0,115,0,110,0,237,0,0,0,0,0,0,0,81,0,0,0,151,0,97,0,100,0,118,0,22,0,0,0,150,0,133,0,0,0,142,0,0,0,206,0,123,0,131,0,0,0,138,0,0,0,74,0,230,0,92,0,168,0,71,0,148,0,32,0,148,0,221,0,41,0,0,0,231,0,122,0,73,0,143,0,166,0,1,0,34,0,103,0,0,0,168,0,111,0,6,0,0,0,18,0,134,0,139,0,169,0,34,0,146,0,0,0,29,0,29,0,0,0,0,0,220,0,138,0,0,0,192,0,0,0,59,0,32,0,93,0,189,0,83,0,166,0,21,0,42,0,246,0,166,0,0,0,0,0,0,0,244,0,88,0,45,0,249,0,77,0,192,0,151,0,116,0,37,0,74,0,244,0,26,0,129,0,232,0,145,0,48,0,0,0,39,0,252,0,37,0,67,0,114,0,205,0,0,0,124,0,115,0,43,0,209,0,249,0,117,0,133,0,140,0,61,0,104,0,38,0,0,0,131,0,58,0,23,0,146,0,98,0,135,0,254,0,4,0,161,0,0,0,212,0);
signal scenario_full  : scenario_type := (0,0,0,0,198,31,242,31,180,31,180,30,111,31,68,31,103,31,251,31,163,31,234,31,21,31,223,31,154,31,154,30,15,31,147,31,128,31,128,30,102,31,243,31,37,31,74,31,27,31,27,30,58,31,197,31,222,31,151,31,218,31,149,31,68,31,144,31,185,31,227,31,190,31,188,31,131,31,188,31,254,31,194,31,70,31,10,31,10,30,196,31,231,31,231,30,163,31,12,31,12,30,119,31,86,31,86,30,64,31,216,31,126,31,217,31,2,31,2,30,2,29,2,28,8,31,48,31,20,31,92,31,97,31,99,31,99,30,21,31,86,31,198,31,198,30,16,31,234,31,18,31,5,31,5,30,220,31,152,31,244,31,36,31,227,31,230,31,225,31,225,30,15,31,86,31,86,30,252,31,26,31,2,31,240,31,149,31,110,31,241,31,233,31,20,31,20,30,237,31,52,31,31,31,240,31,240,30,240,29,93,31,12,31,25,31,153,31,186,31,214,31,185,31,185,30,147,31,111,31,111,30,120,31,212,31,161,31,201,31,74,31,228,31,208,31,208,30,91,31,180,31,116,31,234,31,101,31,80,31,80,30,19,31,19,30,36,31,136,31,13,31,187,31,17,31,17,30,17,29,167,31,167,30,210,31,113,31,73,31,83,31,228,31,228,30,90,31,57,31,187,31,234,31,107,31,220,31,133,31,118,31,81,31,103,31,61,31,96,31,2,31,226,31,68,31,17,31,28,31,28,30,104,31,200,31,49,31,184,31,103,31,155,31,64,31,8,31,111,31,43,31,114,31,195,31,251,31,225,31,254,31,119,31,38,31,3,31,15,31,85,31,124,31,132,31,142,31,207,31,14,31,111,31,224,31,168,31,168,30,236,31,250,31,195,31,138,31,164,31,164,30,157,31,212,31,10,31,194,31,146,31,182,31,151,31,166,31,19,31,129,31,139,31,116,31,61,31,59,31,240,31,123,31,123,30,72,31,177,31,59,31,44,31,44,30,37,31,34,31,145,31,237,31,237,30,27,31,27,30,138,31,109,31,31,31,133,31,68,31,95,31,95,30,95,29,95,28,95,27,176,31,167,31,96,31,165,31,165,31,40,31,199,31,187,31,150,31,201,31,112,31,186,31,85,31,85,30,21,31,40,31,99,31,149,31,51,31,48,31,48,30,14,31,211,31,12,31,207,31,56,31,131,31,72,31,253,31,127,31,127,30,127,29,127,28,7,31,53,31,201,31,91,31,91,30,91,29,91,28,189,31,64,31,242,31,253,31,253,30,72,31,9,31,43,31,184,31,89,31,15,31,32,31,185,31,132,31,252,31,21,31,70,31,142,31,142,30,128,31,5,31,5,30,28,31,16,31,215,31,163,31,253,31,92,31,115,31,234,31,234,30,90,31,140,31,217,31,224,31,150,31,155,31,128,31,61,31,148,31,160,31,188,31,135,31,16,31,99,31,89,31,94,31,242,31,151,31,205,31,121,31,162,31,211,31,183,31,187,31,240,31,239,31,216,31,134,31,146,31,146,30,132,31,113,31,72,31,250,31,187,31,144,31,203,31,83,31,62,31,54,31,224,31,39,31,29,31,29,30,199,31,251,31,251,30,101,31,237,31,150,31,210,31,93,31,46,31,83,31,41,31,208,31,70,31,248,31,180,31,115,31,89,31,102,31,33,31,141,31,14,31,73,31,19,31,5,31,89,31,174,31,211,31,183,31,84,31,84,30,177,31,177,30,11,31,11,30,11,29,70,31,180,31,148,31,242,31,140,31,27,31,155,31,255,31,51,31,51,30,30,31,4,31,64,31,214,31,83,31,29,31,110,31,9,31,24,31,108,31,242,31,171,31,123,31,123,30,129,31,58,31,157,31,149,31,249,31,115,31,9,31,70,31,104,31,104,30,64,31,16,31,103,31,103,30,1,31,53,31,47,31,121,31,231,31,181,31,54,31,5,31,83,31,134,31,168,31,117,31,236,31,199,31,235,31,196,31,109,31,42,31,42,30,240,31,1,31,51,31,163,31,163,30,233,31,191,31,146,31,29,31,221,31,221,30,215,31,164,31,212,31,238,31,91,31,91,30,65,31,65,30,21,31,94,31,213,31,187,31,195,31,182,31,182,30,200,31,232,31,143,31,143,30,247,31,136,31,136,30,136,29,136,28,243,31,43,31,7,31,7,30,72,31,83,31,111,31,16,31,209,31,149,31,141,31,7,31,28,31,28,30,94,31,94,30,94,29,53,31,53,30,83,31,252,31,231,31,247,31,31,31,4,31,243,31,243,30,239,31,239,30,78,31,78,30,16,31,16,30,32,31,87,31,61,31,69,31,181,31,181,30,101,31,200,31,200,30,158,31,179,31,116,31,116,30,137,31,133,31,133,30,140,31,186,31,217,31,131,31,88,31,121,31,111,31,11,31,146,31,214,31,255,31,151,31,151,30,151,29,30,31,60,31,60,30,60,29,60,28,113,31,254,31,167,31,167,30,171,31,105,31,156,31,243,31,243,30,243,29,54,31,130,31,23,31,227,31,215,31,190,31,172,31,153,31,8,31,44,31,231,31,38,31,38,30,224,31,57,31,29,31,99,31,108,31,108,30,121,31,90,31,90,30,89,31,233,31,254,31,222,31,185,31,94,31,241,31,241,30,148,31,82,31,84,31,70,31,71,31,71,30,231,31,18,31,70,31,89,31,225,31,7,31,106,31,106,30,237,31,195,31,103,31,103,30,27,31,131,31,137,31,246,31,198,31,121,31,121,30,121,29,121,28,216,31,202,31,202,30,36,31,187,31,191,31,224,31,215,31,85,31,85,30,209,31,53,31,204,31,182,31,255,31,31,31,2,31,83,31,254,31,254,30,172,31,177,31,138,31,195,31,195,30,121,31,133,31,89,31,165,31,140,31,212,31,212,30,192,31,178,31,178,30,222,31,142,31,98,31,40,31,93,31,89,31,186,31,128,31,134,31,100,31,93,31,246,31,246,30,246,29,45,31,98,31,31,31,190,31,252,31,58,31,156,31,94,31,208,31,208,30,208,29,137,31,137,30,173,31,173,30,203,31,68,31,127,31,127,30,83,31,194,31,245,31,175,31,227,31,202,31,176,31,67,31,3,31,243,31,22,31,187,31,227,31,227,30,146,31,154,31,170,31,95,31,84,31,84,30,212,31,240,31,156,31,235,31,235,30,106,31,164,31,209,31,112,31,4,31,206,31,128,31,246,31,126,31,201,31,75,31,75,30,98,31,211,31,247,31,176,31,114,31,114,30,87,31,67,31,153,31,191,31,107,31,34,31,34,30,34,29,34,28,34,27,34,26,30,31,64,31,27,31,130,31,71,31,71,30,71,29,174,31,61,31,81,31,66,31,66,30,7,31,7,30,176,31,204,31,119,31,119,30,119,29,186,31,186,30,137,31,179,31,37,31,37,30,80,31,184,31,184,30,157,31,25,31,192,31,250,31,250,30,36,31,22,31,22,30,22,29,56,31,56,30,121,31,121,30,121,29,74,31,74,30,199,31,199,30,119,31,172,31,115,31,110,31,237,31,237,30,237,29,237,28,81,31,81,30,151,31,97,31,100,31,118,31,22,31,22,30,150,31,133,31,133,30,142,31,142,30,206,31,123,31,131,31,131,30,138,31,138,30,74,31,230,31,92,31,168,31,71,31,148,31,32,31,148,31,221,31,41,31,41,30,231,31,122,31,73,31,143,31,166,31,1,31,34,31,103,31,103,30,168,31,111,31,6,31,6,30,18,31,134,31,139,31,169,31,34,31,146,31,146,30,29,31,29,31,29,30,29,29,220,31,138,31,138,30,192,31,192,30,59,31,32,31,93,31,189,31,83,31,166,31,21,31,42,31,246,31,166,31,166,30,166,29,166,28,244,31,88,31,45,31,249,31,77,31,192,31,151,31,116,31,37,31,74,31,244,31,26,31,129,31,232,31,145,31,48,31,48,30,39,31,252,31,37,31,67,31,114,31,205,31,205,30,124,31,115,31,43,31,209,31,249,31,117,31,133,31,140,31,61,31,104,31,38,31,38,30,131,31,58,31,23,31,146,31,98,31,135,31,254,31,4,31,161,31,161,30,212,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
