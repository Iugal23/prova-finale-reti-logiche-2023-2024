-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_626 is
end project_tb_626;

architecture project_tb_arch_626 of project_tb_626 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 857;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (92,0,11,0,43,0,133,0,103,0,46,0,0,0,215,0,189,0,244,0,0,0,213,0,148,0,49,0,16,0,38,0,0,0,207,0,115,0,234,0,0,0,105,0,180,0,0,0,116,0,9,0,70,0,74,0,179,0,156,0,198,0,0,0,106,0,131,0,0,0,78,0,122,0,93,0,229,0,142,0,57,0,197,0,0,0,95,0,66,0,161,0,169,0,196,0,154,0,0,0,232,0,141,0,242,0,186,0,194,0,94,0,0,0,29,0,222,0,159,0,59,0,156,0,165,0,28,0,73,0,160,0,192,0,226,0,229,0,22,0,53,0,41,0,135,0,195,0,144,0,13,0,0,0,197,0,0,0,123,0,0,0,180,0,84,0,15,0,0,0,161,0,106,0,122,0,167,0,115,0,16,0,0,0,0,0,191,0,246,0,192,0,47,0,0,0,59,0,0,0,96,0,0,0,200,0,53,0,48,0,146,0,0,0,163,0,187,0,138,0,0,0,224,0,87,0,63,0,31,0,7,0,114,0,111,0,0,0,91,0,52,0,0,0,212,0,11,0,90,0,253,0,144,0,235,0,57,0,44,0,0,0,31,0,0,0,97,0,223,0,58,0,43,0,0,0,27,0,7,0,0,0,180,0,191,0,0,0,0,0,201,0,77,0,108,0,17,0,147,0,230,0,95,0,63,0,137,0,0,0,172,0,151,0,178,0,225,0,0,0,4,0,13,0,75,0,91,0,0,0,121,0,68,0,0,0,163,0,86,0,146,0,0,0,154,0,233,0,160,0,29,0,174,0,31,0,101,0,0,0,143,0,176,0,0,0,218,0,214,0,193,0,218,0,114,0,29,0,72,0,242,0,0,0,40,0,0,0,105,0,96,0,0,0,126,0,0,0,231,0,0,0,215,0,0,0,162,0,242,0,73,0,125,0,236,0,184,0,238,0,0,0,64,0,70,0,148,0,26,0,177,0,0,0,75,0,245,0,218,0,0,0,245,0,23,0,0,0,210,0,127,0,0,0,49,0,161,0,57,0,115,0,235,0,64,0,245,0,234,0,0,0,0,0,88,0,0,0,195,0,144,0,134,0,169,0,140,0,142,0,217,0,194,0,229,0,105,0,167,0,101,0,0,0,109,0,250,0,30,0,175,0,58,0,143,0,92,0,47,0,78,0,181,0,0,0,255,0,0,0,2,0,165,0,247,0,174,0,1,0,95,0,197,0,175,0,105,0,163,0,23,0,235,0,249,0,89,0,164,0,147,0,115,0,63,0,105,0,32,0,51,0,153,0,144,0,67,0,230,0,105,0,205,0,78,0,181,0,227,0,136,0,251,0,110,0,104,0,43,0,104,0,0,0,210,0,73,0,187,0,30,0,169,0,124,0,5,0,204,0,218,0,228,0,237,0,201,0,254,0,120,0,187,0,101,0,0,0,136,0,228,0,152,0,0,0,156,0,0,0,150,0,161,0,106,0,0,0,235,0,83,0,0,0,122,0,35,0,193,0,128,0,0,0,218,0,93,0,46,0,63,0,65,0,0,0,233,0,40,0,235,0,172,0,252,0,0,0,0,0,4,0,3,0,0,0,139,0,158,0,12,0,0,0,0,0,253,0,103,0,162,0,68,0,0,0,0,0,0,0,0,0,93,0,38,0,184,0,93,0,0,0,141,0,149,0,215,0,78,0,128,0,0,0,26,0,188,0,137,0,4,0,145,0,192,0,0,0,203,0,57,0,252,0,46,0,109,0,134,0,136,0,191,0,213,0,167,0,43,0,0,0,0,0,0,0,108,0,147,0,170,0,61,0,81,0,233,0,0,0,1,0,136,0,147,0,143,0,115,0,132,0,151,0,228,0,23,0,76,0,235,0,74,0,153,0,31,0,123,0,30,0,53,0,175,0,89,0,80,0,101,0,46,0,244,0,0,0,8,0,205,0,148,0,192,0,0,0,0,0,184,0,49,0,253,0,74,0,98,0,196,0,0,0,205,0,17,0,132,0,174,0,60,0,104,0,0,0,209,0,210,0,86,0,0,0,0,0,227,0,206,0,162,0,6,0,96,0,32,0,57,0,0,0,141,0,0,0,116,0,211,0,45,0,0,0,9,0,0,0,25,0,64,0,28,0,208,0,125,0,216,0,60,0,115,0,157,0,157,0,104,0,30,0,0,0,81,0,0,0,90,0,111,0,250,0,0,0,92,0,0,0,206,0,153,0,247,0,50,0,43,0,0,0,185,0,214,0,228,0,214,0,200,0,123,0,114,0,182,0,191,0,74,0,0,0,94,0,162,0,28,0,162,0,253,0,0,0,146,0,0,0,62,0,0,0,188,0,0,0,0,0,91,0,136,0,155,0,129,0,67,0,6,0,58,0,80,0,217,0,137,0,13,0,178,0,0,0,36,0,94,0,211,0,188,0,14,0,172,0,78,0,147,0,148,0,0,0,254,0,134,0,199,0,189,0,123,0,4,0,0,0,0,0,0,0,3,0,189,0,131,0,72,0,235,0,253,0,241,0,208,0,11,0,1,0,0,0,244,0,252,0,12,0,104,0,249,0,37,0,0,0,0,0,126,0,88,0,232,0,0,0,217,0,108,0,22,0,188,0,237,0,190,0,143,0,164,0,189,0,138,0,187,0,77,0,0,0,0,0,226,0,193,0,0,0,224,0,0,0,0,0,0,0,128,0,18,0,204,0,181,0,191,0,62,0,240,0,168,0,64,0,0,0,65,0,152,0,165,0,30,0,67,0,200,0,236,0,232,0,110,0,84,0,44,0,57,0,27,0,169,0,68,0,146,0,0,0,149,0,0,0,86,0,232,0,98,0,200,0,0,0,0,0,33,0,169,0,101,0,23,0,0,0,69,0,183,0,185,0,245,0,0,0,226,0,62,0,90,0,235,0,156,0,29,0,29,0,110,0,32,0,142,0,0,0,188,0,52,0,105,0,106,0,0,0,0,0,188,0,28,0,74,0,210,0,0,0,98,0,112,0,34,0,0,0,0,0,8,0,121,0,157,0,64,0,226,0,175,0,160,0,91,0,0,0,235,0,246,0,187,0,1,0,246,0,128,0,69,0,128,0,251,0,72,0,2,0,152,0,174,0,191,0,109,0,139,0,152,0,0,0,46,0,4,0,101,0,122,0,18,0,151,0,243,0,181,0,234,0,0,0,97,0,0,0,15,0,213,0,0,0,71,0,152,0,138,0,110,0,177,0,14,0,118,0,56,0,163,0,174,0,8,0,224,0,0,0,0,0,16,0,150,0,91,0,62,0,89,0,0,0,94,0,242,0,227,0,100,0,14,0,146,0,49,0,0,0,137,0,0,0,192,0,252,0,117,0,141,0,35,0,251,0,214,0,0,0,233,0,195,0,189,0,154,0,0,0,0,0,6,0,19,0,164,0,46,0,104,0,191,0,0,0,65,0,197,0,109,0,0,0,0,0,3,0,112,0,254,0,52,0,0,0,48,0,218,0,229,0,0,0,0,0,115,0,47,0,208,0,235,0,122,0,30,0,92,0,51,0,106,0,83,0,232,0,158,0,45,0,57,0,211,0,0,0,152,0,0,0,43,0,255,0,98,0,25,0,0,0,200,0,232,0,39,0,142,0,90,0,75,0,123,0,63,0,19,0,92,0,33,0,0,0,135,0,4,0,176,0,132,0,160,0,108,0,104,0,94,0,250,0,218,0,213,0,84,0,36,0,127,0,142,0,0,0,110,0,225,0,117,0,210,0,0,0,131,0,157,0,215,0,208,0,0,0,101,0,126,0,164,0,0,0,78,0,218,0,0,0,0,0,133,0,105,0,0,0,77,0,197,0,223,0,187,0,244,0,250,0,238,0,194,0);
signal scenario_full  : scenario_type := (92,31,11,31,43,31,133,31,103,31,46,31,46,30,215,31,189,31,244,31,244,30,213,31,148,31,49,31,16,31,38,31,38,30,207,31,115,31,234,31,234,30,105,31,180,31,180,30,116,31,9,31,70,31,74,31,179,31,156,31,198,31,198,30,106,31,131,31,131,30,78,31,122,31,93,31,229,31,142,31,57,31,197,31,197,30,95,31,66,31,161,31,169,31,196,31,154,31,154,30,232,31,141,31,242,31,186,31,194,31,94,31,94,30,29,31,222,31,159,31,59,31,156,31,165,31,28,31,73,31,160,31,192,31,226,31,229,31,22,31,53,31,41,31,135,31,195,31,144,31,13,31,13,30,197,31,197,30,123,31,123,30,180,31,84,31,15,31,15,30,161,31,106,31,122,31,167,31,115,31,16,31,16,30,16,29,191,31,246,31,192,31,47,31,47,30,59,31,59,30,96,31,96,30,200,31,53,31,48,31,146,31,146,30,163,31,187,31,138,31,138,30,224,31,87,31,63,31,31,31,7,31,114,31,111,31,111,30,91,31,52,31,52,30,212,31,11,31,90,31,253,31,144,31,235,31,57,31,44,31,44,30,31,31,31,30,97,31,223,31,58,31,43,31,43,30,27,31,7,31,7,30,180,31,191,31,191,30,191,29,201,31,77,31,108,31,17,31,147,31,230,31,95,31,63,31,137,31,137,30,172,31,151,31,178,31,225,31,225,30,4,31,13,31,75,31,91,31,91,30,121,31,68,31,68,30,163,31,86,31,146,31,146,30,154,31,233,31,160,31,29,31,174,31,31,31,101,31,101,30,143,31,176,31,176,30,218,31,214,31,193,31,218,31,114,31,29,31,72,31,242,31,242,30,40,31,40,30,105,31,96,31,96,30,126,31,126,30,231,31,231,30,215,31,215,30,162,31,242,31,73,31,125,31,236,31,184,31,238,31,238,30,64,31,70,31,148,31,26,31,177,31,177,30,75,31,245,31,218,31,218,30,245,31,23,31,23,30,210,31,127,31,127,30,49,31,161,31,57,31,115,31,235,31,64,31,245,31,234,31,234,30,234,29,88,31,88,30,195,31,144,31,134,31,169,31,140,31,142,31,217,31,194,31,229,31,105,31,167,31,101,31,101,30,109,31,250,31,30,31,175,31,58,31,143,31,92,31,47,31,78,31,181,31,181,30,255,31,255,30,2,31,165,31,247,31,174,31,1,31,95,31,197,31,175,31,105,31,163,31,23,31,235,31,249,31,89,31,164,31,147,31,115,31,63,31,105,31,32,31,51,31,153,31,144,31,67,31,230,31,105,31,205,31,78,31,181,31,227,31,136,31,251,31,110,31,104,31,43,31,104,31,104,30,210,31,73,31,187,31,30,31,169,31,124,31,5,31,204,31,218,31,228,31,237,31,201,31,254,31,120,31,187,31,101,31,101,30,136,31,228,31,152,31,152,30,156,31,156,30,150,31,161,31,106,31,106,30,235,31,83,31,83,30,122,31,35,31,193,31,128,31,128,30,218,31,93,31,46,31,63,31,65,31,65,30,233,31,40,31,235,31,172,31,252,31,252,30,252,29,4,31,3,31,3,30,139,31,158,31,12,31,12,30,12,29,253,31,103,31,162,31,68,31,68,30,68,29,68,28,68,27,93,31,38,31,184,31,93,31,93,30,141,31,149,31,215,31,78,31,128,31,128,30,26,31,188,31,137,31,4,31,145,31,192,31,192,30,203,31,57,31,252,31,46,31,109,31,134,31,136,31,191,31,213,31,167,31,43,31,43,30,43,29,43,28,108,31,147,31,170,31,61,31,81,31,233,31,233,30,1,31,136,31,147,31,143,31,115,31,132,31,151,31,228,31,23,31,76,31,235,31,74,31,153,31,31,31,123,31,30,31,53,31,175,31,89,31,80,31,101,31,46,31,244,31,244,30,8,31,205,31,148,31,192,31,192,30,192,29,184,31,49,31,253,31,74,31,98,31,196,31,196,30,205,31,17,31,132,31,174,31,60,31,104,31,104,30,209,31,210,31,86,31,86,30,86,29,227,31,206,31,162,31,6,31,96,31,32,31,57,31,57,30,141,31,141,30,116,31,211,31,45,31,45,30,9,31,9,30,25,31,64,31,28,31,208,31,125,31,216,31,60,31,115,31,157,31,157,31,104,31,30,31,30,30,81,31,81,30,90,31,111,31,250,31,250,30,92,31,92,30,206,31,153,31,247,31,50,31,43,31,43,30,185,31,214,31,228,31,214,31,200,31,123,31,114,31,182,31,191,31,74,31,74,30,94,31,162,31,28,31,162,31,253,31,253,30,146,31,146,30,62,31,62,30,188,31,188,30,188,29,91,31,136,31,155,31,129,31,67,31,6,31,58,31,80,31,217,31,137,31,13,31,178,31,178,30,36,31,94,31,211,31,188,31,14,31,172,31,78,31,147,31,148,31,148,30,254,31,134,31,199,31,189,31,123,31,4,31,4,30,4,29,4,28,3,31,189,31,131,31,72,31,235,31,253,31,241,31,208,31,11,31,1,31,1,30,244,31,252,31,12,31,104,31,249,31,37,31,37,30,37,29,126,31,88,31,232,31,232,30,217,31,108,31,22,31,188,31,237,31,190,31,143,31,164,31,189,31,138,31,187,31,77,31,77,30,77,29,226,31,193,31,193,30,224,31,224,30,224,29,224,28,128,31,18,31,204,31,181,31,191,31,62,31,240,31,168,31,64,31,64,30,65,31,152,31,165,31,30,31,67,31,200,31,236,31,232,31,110,31,84,31,44,31,57,31,27,31,169,31,68,31,146,31,146,30,149,31,149,30,86,31,232,31,98,31,200,31,200,30,200,29,33,31,169,31,101,31,23,31,23,30,69,31,183,31,185,31,245,31,245,30,226,31,62,31,90,31,235,31,156,31,29,31,29,31,110,31,32,31,142,31,142,30,188,31,52,31,105,31,106,31,106,30,106,29,188,31,28,31,74,31,210,31,210,30,98,31,112,31,34,31,34,30,34,29,8,31,121,31,157,31,64,31,226,31,175,31,160,31,91,31,91,30,235,31,246,31,187,31,1,31,246,31,128,31,69,31,128,31,251,31,72,31,2,31,152,31,174,31,191,31,109,31,139,31,152,31,152,30,46,31,4,31,101,31,122,31,18,31,151,31,243,31,181,31,234,31,234,30,97,31,97,30,15,31,213,31,213,30,71,31,152,31,138,31,110,31,177,31,14,31,118,31,56,31,163,31,174,31,8,31,224,31,224,30,224,29,16,31,150,31,91,31,62,31,89,31,89,30,94,31,242,31,227,31,100,31,14,31,146,31,49,31,49,30,137,31,137,30,192,31,252,31,117,31,141,31,35,31,251,31,214,31,214,30,233,31,195,31,189,31,154,31,154,30,154,29,6,31,19,31,164,31,46,31,104,31,191,31,191,30,65,31,197,31,109,31,109,30,109,29,3,31,112,31,254,31,52,31,52,30,48,31,218,31,229,31,229,30,229,29,115,31,47,31,208,31,235,31,122,31,30,31,92,31,51,31,106,31,83,31,232,31,158,31,45,31,57,31,211,31,211,30,152,31,152,30,43,31,255,31,98,31,25,31,25,30,200,31,232,31,39,31,142,31,90,31,75,31,123,31,63,31,19,31,92,31,33,31,33,30,135,31,4,31,176,31,132,31,160,31,108,31,104,31,94,31,250,31,218,31,213,31,84,31,36,31,127,31,142,31,142,30,110,31,225,31,117,31,210,31,210,30,131,31,157,31,215,31,208,31,208,30,101,31,126,31,164,31,164,30,78,31,218,31,218,30,218,29,133,31,105,31,105,30,77,31,197,31,223,31,187,31,244,31,250,31,238,31,194,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
