-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_710 is
end project_tb_710;

architecture project_tb_arch_710 of project_tb_710 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 225;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (45,0,61,0,63,0,0,0,109,0,241,0,238,0,32,0,25,0,211,0,143,0,176,0,202,0,102,0,172,0,34,0,248,0,92,0,0,0,190,0,0,0,210,0,194,0,227,0,135,0,253,0,237,0,218,0,0,0,0,0,48,0,63,0,209,0,243,0,60,0,84,0,186,0,253,0,244,0,0,0,68,0,95,0,248,0,102,0,0,0,42,0,79,0,0,0,35,0,62,0,134,0,243,0,204,0,13,0,74,0,32,0,0,0,0,0,199,0,78,0,43,0,76,0,9,0,214,0,0,0,207,0,0,0,211,0,22,0,6,0,225,0,212,0,0,0,97,0,4,0,156,0,51,0,230,0,12,0,140,0,185,0,218,0,0,0,72,0,255,0,80,0,0,0,18,0,193,0,45,0,33,0,3,0,159,0,0,0,124,0,40,0,224,0,58,0,254,0,125,0,3,0,107,0,186,0,247,0,236,0,0,0,0,0,89,0,70,0,98,0,58,0,73,0,0,0,230,0,214,0,0,0,46,0,118,0,146,0,211,0,22,0,142,0,54,0,25,0,128,0,18,0,242,0,113,0,145,0,0,0,229,0,229,0,230,0,0,0,0,0,135,0,0,0,203,0,65,0,223,0,0,0,171,0,101,0,0,0,78,0,218,0,206,0,181,0,125,0,229,0,0,0,72,0,239,0,156,0,246,0,221,0,41,0,136,0,139,0,140,0,90,0,39,0,71,0,40,0,89,0,195,0,182,0,140,0,127,0,181,0,185,0,244,0,28,0,0,0,221,0,14,0,143,0,0,0,13,0,237,0,80,0,72,0,213,0,66,0,234,0,83,0,137,0,90,0,0,0,0,0,153,0,51,0,90,0,94,0,41,0,149,0,243,0,49,0,152,0,52,0,118,0,0,0,0,0,194,0,196,0,59,0,40,0,167,0,179,0,0,0,59,0,63,0,252,0,249,0,123,0,107,0,189,0,242,0,119,0,237,0,154,0,3,0,197,0,173,0,86,0);
signal scenario_full  : scenario_type := (45,31,61,31,63,31,63,30,109,31,241,31,238,31,32,31,25,31,211,31,143,31,176,31,202,31,102,31,172,31,34,31,248,31,92,31,92,30,190,31,190,30,210,31,194,31,227,31,135,31,253,31,237,31,218,31,218,30,218,29,48,31,63,31,209,31,243,31,60,31,84,31,186,31,253,31,244,31,244,30,68,31,95,31,248,31,102,31,102,30,42,31,79,31,79,30,35,31,62,31,134,31,243,31,204,31,13,31,74,31,32,31,32,30,32,29,199,31,78,31,43,31,76,31,9,31,214,31,214,30,207,31,207,30,211,31,22,31,6,31,225,31,212,31,212,30,97,31,4,31,156,31,51,31,230,31,12,31,140,31,185,31,218,31,218,30,72,31,255,31,80,31,80,30,18,31,193,31,45,31,33,31,3,31,159,31,159,30,124,31,40,31,224,31,58,31,254,31,125,31,3,31,107,31,186,31,247,31,236,31,236,30,236,29,89,31,70,31,98,31,58,31,73,31,73,30,230,31,214,31,214,30,46,31,118,31,146,31,211,31,22,31,142,31,54,31,25,31,128,31,18,31,242,31,113,31,145,31,145,30,229,31,229,31,230,31,230,30,230,29,135,31,135,30,203,31,65,31,223,31,223,30,171,31,101,31,101,30,78,31,218,31,206,31,181,31,125,31,229,31,229,30,72,31,239,31,156,31,246,31,221,31,41,31,136,31,139,31,140,31,90,31,39,31,71,31,40,31,89,31,195,31,182,31,140,31,127,31,181,31,185,31,244,31,28,31,28,30,221,31,14,31,143,31,143,30,13,31,237,31,80,31,72,31,213,31,66,31,234,31,83,31,137,31,90,31,90,30,90,29,153,31,51,31,90,31,94,31,41,31,149,31,243,31,49,31,152,31,52,31,118,31,118,30,118,29,194,31,196,31,59,31,40,31,167,31,179,31,179,30,59,31,63,31,252,31,249,31,123,31,107,31,189,31,242,31,119,31,237,31,154,31,3,31,197,31,173,31,86,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
