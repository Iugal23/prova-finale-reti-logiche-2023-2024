-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_713 is
end project_tb_713;

architecture project_tb_arch_713 of project_tb_713 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 421;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (117,0,0,0,173,0,157,0,27,0,110,0,120,0,223,0,86,0,155,0,46,0,0,0,191,0,0,0,0,0,117,0,104,0,0,0,0,0,173,0,55,0,0,0,253,0,166,0,221,0,96,0,254,0,0,0,212,0,0,0,0,0,0,0,41,0,160,0,28,0,86,0,215,0,0,0,243,0,163,0,13,0,167,0,193,0,86,0,255,0,130,0,203,0,16,0,186,0,252,0,205,0,106,0,37,0,210,0,0,0,172,0,136,0,69,0,0,0,181,0,0,0,0,0,153,0,45,0,184,0,110,0,208,0,0,0,0,0,137,0,153,0,2,0,131,0,153,0,0,0,141,0,44,0,61,0,28,0,95,0,105,0,0,0,170,0,0,0,21,0,244,0,74,0,97,0,143,0,238,0,57,0,128,0,71,0,0,0,96,0,66,0,214,0,0,0,108,0,159,0,195,0,187,0,43,0,0,0,0,0,33,0,140,0,0,0,0,0,92,0,142,0,60,0,135,0,215,0,30,0,86,0,114,0,206,0,162,0,251,0,96,0,212,0,180,0,165,0,96,0,0,0,50,0,90,0,42,0,45,0,0,0,141,0,0,0,97,0,0,0,237,0,42,0,70,0,0,0,120,0,107,0,104,0,109,0,25,0,87,0,112,0,86,0,26,0,102,0,247,0,136,0,132,0,151,0,114,0,19,0,254,0,78,0,0,0,0,0,184,0,76,0,214,0,225,0,162,0,234,0,221,0,0,0,133,0,0,0,153,0,1,0,90,0,234,0,0,0,0,0,240,0,222,0,0,0,84,0,203,0,66,0,0,0,150,0,24,0,103,0,0,0,244,0,55,0,99,0,194,0,0,0,0,0,159,0,212,0,248,0,202,0,169,0,32,0,145,0,242,0,195,0,152,0,58,0,121,0,0,0,215,0,13,0,0,0,50,0,0,0,118,0,0,0,26,0,0,0,111,0,163,0,0,0,9,0,53,0,92,0,135,0,207,0,134,0,226,0,239,0,172,0,0,0,67,0,51,0,152,0,125,0,124,0,72,0,111,0,0,0,103,0,98,0,175,0,0,0,172,0,101,0,0,0,34,0,25,0,147,0,0,0,104,0,0,0,0,0,5,0,78,0,0,0,109,0,89,0,69,0,46,0,192,0,35,0,213,0,0,0,244,0,0,0,83,0,0,0,0,0,0,0,4,0,0,0,10,0,104,0,248,0,152,0,86,0,162,0,49,0,27,0,25,0,48,0,92,0,0,0,115,0,244,0,72,0,0,0,9,0,0,0,235,0,18,0,62,0,77,0,193,0,198,0,26,0,81,0,57,0,240,0,0,0,0,0,82,0,201,0,49,0,3,0,0,0,53,0,45,0,89,0,45,0,207,0,235,0,139,0,251,0,62,0,53,0,253,0,0,0,147,0,224,0,50,0,111,0,55,0,178,0,82,0,0,0,194,0,136,0,126,0,46,0,195,0,117,0,102,0,149,0,0,0,0,0,8,0,0,0,159,0,118,0,216,0,59,0,255,0,0,0,37,0,128,0,9,0,239,0,141,0,38,0,74,0,80,0,200,0,0,0,0,0,48,0,49,0,0,0,0,0,225,0,16,0,66,0,29,0,0,0,66,0,191,0,218,0,253,0,107,0,116,0,84,0,251,0,0,0,157,0,231,0,239,0,216,0,51,0,75,0,170,0,9,0,0,0,22,0,30,0,22,0,0,0,129,0,151,0,227,0,208,0,14,0,0,0,176,0,6,0,154,0,206,0,66,0,0,0,118,0,185,0,0,0,36,0,108,0,230,0,229,0,34,0,118,0,243,0,2,0,13,0,190,0,0,0,0,0,193,0,0,0,205,0,208,0,249,0,125,0,0,0,0,0,244,0,31,0,42,0);
signal scenario_full  : scenario_type := (117,31,117,30,173,31,157,31,27,31,110,31,120,31,223,31,86,31,155,31,46,31,46,30,191,31,191,30,191,29,117,31,104,31,104,30,104,29,173,31,55,31,55,30,253,31,166,31,221,31,96,31,254,31,254,30,212,31,212,30,212,29,212,28,41,31,160,31,28,31,86,31,215,31,215,30,243,31,163,31,13,31,167,31,193,31,86,31,255,31,130,31,203,31,16,31,186,31,252,31,205,31,106,31,37,31,210,31,210,30,172,31,136,31,69,31,69,30,181,31,181,30,181,29,153,31,45,31,184,31,110,31,208,31,208,30,208,29,137,31,153,31,2,31,131,31,153,31,153,30,141,31,44,31,61,31,28,31,95,31,105,31,105,30,170,31,170,30,21,31,244,31,74,31,97,31,143,31,238,31,57,31,128,31,71,31,71,30,96,31,66,31,214,31,214,30,108,31,159,31,195,31,187,31,43,31,43,30,43,29,33,31,140,31,140,30,140,29,92,31,142,31,60,31,135,31,215,31,30,31,86,31,114,31,206,31,162,31,251,31,96,31,212,31,180,31,165,31,96,31,96,30,50,31,90,31,42,31,45,31,45,30,141,31,141,30,97,31,97,30,237,31,42,31,70,31,70,30,120,31,107,31,104,31,109,31,25,31,87,31,112,31,86,31,26,31,102,31,247,31,136,31,132,31,151,31,114,31,19,31,254,31,78,31,78,30,78,29,184,31,76,31,214,31,225,31,162,31,234,31,221,31,221,30,133,31,133,30,153,31,1,31,90,31,234,31,234,30,234,29,240,31,222,31,222,30,84,31,203,31,66,31,66,30,150,31,24,31,103,31,103,30,244,31,55,31,99,31,194,31,194,30,194,29,159,31,212,31,248,31,202,31,169,31,32,31,145,31,242,31,195,31,152,31,58,31,121,31,121,30,215,31,13,31,13,30,50,31,50,30,118,31,118,30,26,31,26,30,111,31,163,31,163,30,9,31,53,31,92,31,135,31,207,31,134,31,226,31,239,31,172,31,172,30,67,31,51,31,152,31,125,31,124,31,72,31,111,31,111,30,103,31,98,31,175,31,175,30,172,31,101,31,101,30,34,31,25,31,147,31,147,30,104,31,104,30,104,29,5,31,78,31,78,30,109,31,89,31,69,31,46,31,192,31,35,31,213,31,213,30,244,31,244,30,83,31,83,30,83,29,83,28,4,31,4,30,10,31,104,31,248,31,152,31,86,31,162,31,49,31,27,31,25,31,48,31,92,31,92,30,115,31,244,31,72,31,72,30,9,31,9,30,235,31,18,31,62,31,77,31,193,31,198,31,26,31,81,31,57,31,240,31,240,30,240,29,82,31,201,31,49,31,3,31,3,30,53,31,45,31,89,31,45,31,207,31,235,31,139,31,251,31,62,31,53,31,253,31,253,30,147,31,224,31,50,31,111,31,55,31,178,31,82,31,82,30,194,31,136,31,126,31,46,31,195,31,117,31,102,31,149,31,149,30,149,29,8,31,8,30,159,31,118,31,216,31,59,31,255,31,255,30,37,31,128,31,9,31,239,31,141,31,38,31,74,31,80,31,200,31,200,30,200,29,48,31,49,31,49,30,49,29,225,31,16,31,66,31,29,31,29,30,66,31,191,31,218,31,253,31,107,31,116,31,84,31,251,31,251,30,157,31,231,31,239,31,216,31,51,31,75,31,170,31,9,31,9,30,22,31,30,31,22,31,22,30,129,31,151,31,227,31,208,31,14,31,14,30,176,31,6,31,154,31,206,31,66,31,66,30,118,31,185,31,185,30,36,31,108,31,230,31,229,31,34,31,118,31,243,31,2,31,13,31,190,31,190,30,190,29,193,31,193,30,205,31,208,31,249,31,125,31,125,30,125,29,244,31,31,31,42,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
