-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_706 is
end project_tb_706;

architecture project_tb_arch_706 of project_tb_706 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 200;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (100,0,189,0,32,0,0,0,197,0,0,0,59,0,184,0,148,0,182,0,116,0,0,0,13,0,37,0,74,0,66,0,41,0,0,0,35,0,179,0,193,0,100,0,54,0,78,0,134,0,132,0,0,0,0,0,38,0,13,0,129,0,66,0,0,0,0,0,246,0,213,0,223,0,55,0,174,0,252,0,62,0,0,0,140,0,203,0,189,0,10,0,177,0,0,0,16,0,42,0,23,0,0,0,39,0,0,0,0,0,0,0,248,0,47,0,218,0,20,0,0,0,247,0,193,0,230,0,0,0,13,0,0,0,241,0,90,0,132,0,162,0,91,0,240,0,0,0,63,0,22,0,0,0,28,0,249,0,7,0,185,0,0,0,123,0,198,0,0,0,0,0,221,0,30,0,54,0,79,0,0,0,218,0,254,0,217,0,175,0,78,0,236,0,42,0,0,0,25,0,119,0,149,0,180,0,0,0,142,0,218,0,148,0,19,0,234,0,62,0,124,0,216,0,127,0,0,0,56,0,0,0,83,0,0,0,64,0,2,0,5,0,215,0,245,0,166,0,92,0,2,0,36,0,12,0,144,0,233,0,101,0,241,0,0,0,134,0,19,0,245,0,19,0,0,0,147,0,187,0,125,0,0,0,254,0,181,0,11,0,114,0,206,0,67,0,96,0,29,0,62,0,149,0,76,0,167,0,133,0,0,0,144,0,69,0,165,0,190,0,220,0,52,0,167,0,32,0,144,0,196,0,255,0,34,0,132,0,0,0,82,0,0,0,244,0,176,0,26,0,0,0,238,0,89,0,102,0,109,0,11,0,140,0,0,0,222,0,44,0,163,0,121,0,0,0,102,0,135,0,84,0,204,0,0,0,122,0,0,0,206,0,0,0,116,0,139,0,76,0);
signal scenario_full  : scenario_type := (100,31,189,31,32,31,32,30,197,31,197,30,59,31,184,31,148,31,182,31,116,31,116,30,13,31,37,31,74,31,66,31,41,31,41,30,35,31,179,31,193,31,100,31,54,31,78,31,134,31,132,31,132,30,132,29,38,31,13,31,129,31,66,31,66,30,66,29,246,31,213,31,223,31,55,31,174,31,252,31,62,31,62,30,140,31,203,31,189,31,10,31,177,31,177,30,16,31,42,31,23,31,23,30,39,31,39,30,39,29,39,28,248,31,47,31,218,31,20,31,20,30,247,31,193,31,230,31,230,30,13,31,13,30,241,31,90,31,132,31,162,31,91,31,240,31,240,30,63,31,22,31,22,30,28,31,249,31,7,31,185,31,185,30,123,31,198,31,198,30,198,29,221,31,30,31,54,31,79,31,79,30,218,31,254,31,217,31,175,31,78,31,236,31,42,31,42,30,25,31,119,31,149,31,180,31,180,30,142,31,218,31,148,31,19,31,234,31,62,31,124,31,216,31,127,31,127,30,56,31,56,30,83,31,83,30,64,31,2,31,5,31,215,31,245,31,166,31,92,31,2,31,36,31,12,31,144,31,233,31,101,31,241,31,241,30,134,31,19,31,245,31,19,31,19,30,147,31,187,31,125,31,125,30,254,31,181,31,11,31,114,31,206,31,67,31,96,31,29,31,62,31,149,31,76,31,167,31,133,31,133,30,144,31,69,31,165,31,190,31,220,31,52,31,167,31,32,31,144,31,196,31,255,31,34,31,132,31,132,30,82,31,82,30,244,31,176,31,26,31,26,30,238,31,89,31,102,31,109,31,11,31,140,31,140,30,222,31,44,31,163,31,121,31,121,30,102,31,135,31,84,31,204,31,204,30,122,31,122,30,206,31,206,30,116,31,139,31,76,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
