-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 948;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (3,0,0,0,0,0,90,0,50,0,153,0,152,0,252,0,201,0,15,0,112,0,0,0,250,0,0,0,158,0,0,0,57,0,0,0,252,0,0,0,170,0,188,0,196,0,225,0,192,0,3,0,48,0,0,0,159,0,124,0,35,0,55,0,104,0,150,0,203,0,0,0,0,0,151,0,165,0,247,0,5,0,133,0,11,0,151,0,64,0,3,0,139,0,208,0,0,0,117,0,84,0,136,0,130,0,38,0,146,0,184,0,145,0,55,0,177,0,133,0,108,0,251,0,84,0,54,0,65,0,190,0,32,0,226,0,0,0,83,0,38,0,75,0,0,0,120,0,185,0,69,0,67,0,142,0,17,0,136,0,25,0,0,0,76,0,134,0,0,0,0,0,199,0,245,0,0,0,100,0,120,0,0,0,89,0,0,0,129,0,107,0,19,0,130,0,104,0,133,0,164,0,23,0,229,0,249,0,151,0,0,0,201,0,188,0,46,0,180,0,0,0,230,0,137,0,221,0,209,0,69,0,98,0,123,0,139,0,172,0,1,0,155,0,155,0,59,0,4,0,193,0,0,0,132,0,63,0,10,0,70,0,220,0,103,0,108,0,186,0,54,0,166,0,0,0,27,0,0,0,246,0,201,0,233,0,0,0,51,0,24,0,64,0,238,0,221,0,186,0,191,0,200,0,16,0,0,0,249,0,94,0,21,0,246,0,80,0,94,0,53,0,100,0,11,0,0,0,44,0,148,0,141,0,0,0,203,0,0,0,241,0,108,0,93,0,46,0,4,0,56,0,130,0,79,0,164,0,2,0,231,0,139,0,80,0,89,0,48,0,150,0,219,0,255,0,11,0,116,0,33,0,116,0,3,0,73,0,202,0,58,0,252,0,171,0,89,0,0,0,238,0,163,0,211,0,98,0,130,0,46,0,129,0,255,0,0,0,65,0,44,0,250,0,55,0,249,0,0,0,0,0,205,0,96,0,166,0,196,0,25,0,0,0,41,0,230,0,37,0,181,0,123,0,172,0,246,0,0,0,74,0,160,0,0,0,25,0,0,0,225,0,206,0,123,0,69,0,5,0,130,0,0,0,130,0,137,0,2,0,0,0,224,0,0,0,161,0,83,0,227,0,0,0,215,0,161,0,102,0,76,0,89,0,0,0,162,0,138,0,191,0,14,0,134,0,76,0,0,0,230,0,0,0,0,0,98,0,164,0,152,0,113,0,37,0,29,0,0,0,163,0,173,0,114,0,207,0,57,0,226,0,0,0,72,0,96,0,0,0,55,0,66,0,0,0,184,0,236,0,226,0,248,0,40,0,0,0,41,0,16,0,164,0,193,0,1,0,0,0,255,0,0,0,212,0,238,0,85,0,122,0,128,0,0,0,110,0,119,0,8,0,165,0,0,0,45,0,105,0,36,0,21,0,0,0,24,0,77,0,86,0,0,0,102,0,0,0,81,0,0,0,179,0,127,0,202,0,54,0,16,0,67,0,103,0,86,0,88,0,151,0,30,0,57,0,71,0,56,0,2,0,91,0,0,0,92,0,85,0,0,0,26,0,253,0,6,0,238,0,212,0,208,0,47,0,139,0,155,0,0,0,207,0,48,0,112,0,131,0,202,0,0,0,171,0,147,0,0,0,0,0,246,0,174,0,38,0,230,0,202,0,206,0,137,0,30,0,0,0,177,0,6,0,41,0,42,0,0,0,0,0,0,0,91,0,106,0,100,0,6,0,0,0,69,0,33,0,30,0,106,0,117,0,0,0,162,0,67,0,151,0,152,0,22,0,243,0,0,0,102,0,236,0,211,0,181,0,99,0,37,0,77,0,105,0,217,0,161,0,244,0,93,0,5,0,220,0,164,0,189,0,196,0,159,0,145,0,0,0,146,0,230,0,216,0,124,0,55,0,19,0,84,0,0,0,107,0,0,0,124,0,35,0,0,0,0,0,63,0,206,0,0,0,3,0,0,0,0,0,1,0,171,0,243,0,193,0,88,0,0,0,184,0,127,0,216,0,0,0,0,0,0,0,97,0,42,0,0,0,0,0,23,0,116,0,233,0,245,0,95,0,227,0,204,0,182,0,199,0,78,0,242,0,0,0,0,0,102,0,165,0,201,0,254,0,207,0,0,0,58,0,162,0,60,0,0,0,231,0,0,0,0,0,0,0,0,0,0,0,26,0,49,0,20,0,224,0,179,0,2,0,80,0,57,0,229,0,116,0,4,0,180,0,0,0,0,0,133,0,88,0,198,0,5,0,94,0,84,0,232,0,30,0,148,0,183,0,193,0,15,0,27,0,207,0,115,0,58,0,2,0,168,0,197,0,102,0,149,0,21,0,0,0,184,0,75,0,80,0,210,0,69,0,240,0,89,0,91,0,240,0,191,0,113,0,38,0,34,0,179,0,92,0,157,0,0,0,81,0,110,0,114,0,0,0,213,0,0,0,0,0,26,0,7,0,0,0,127,0,254,0,176,0,0,0,0,0,60,0,231,0,0,0,0,0,140,0,130,0,210,0,69,0,101,0,13,0,29,0,64,0,31,0,120,0,63,0,83,0,181,0,0,0,254,0,127,0,10,0,63,0,228,0,229,0,248,0,104,0,120,0,180,0,56,0,0,0,117,0,154,0,0,0,0,0,223,0,162,0,9,0,140,0,186,0,58,0,28,0,139,0,85,0,212,0,123,0,72,0,163,0,114,0,177,0,166,0,197,0,0,0,79,0,34,0,214,0,98,0,104,0,201,0,96,0,0,0,230,0,0,0,114,0,114,0,114,0,9,0,0,0,0,0,150,0,27,0,0,0,23,0,216,0,122,0,156,0,111,0,91,0,143,0,209,0,93,0,225,0,161,0,228,0,0,0,178,0,66,0,0,0,89,0,45,0,124,0,132,0,54,0,71,0,20,0,57,0,201,0,189,0,95,0,96,0,245,0,0,0,60,0,0,0,242,0,185,0,56,0,0,0,193,0,180,0,65,0,82,0,149,0,171,0,219,0,162,0,12,0,184,0,12,0,93,0,210,0,0,0,206,0,0,0,88,0,81,0,0,0,0,0,0,0,200,0,126,0,0,0,0,0,160,0,153,0,0,0,0,0,71,0,242,0,126,0,77,0,213,0,0,0,66,0,124,0,60,0,0,0,253,0,160,0,131,0,44,0,0,0,213,0,188,0,28,0,101,0,0,0,214,0,55,0,0,0,43,0,43,0,65,0,104,0,0,0,181,0,236,0,78,0,106,0,29,0,207,0,105,0,109,0,0,0,48,0,244,0,163,0,0,0,91,0,58,0,109,0,111,0,243,0,108,0,56,0,233,0,150,0,0,0,82,0,0,0,151,0,176,0,0,0,254,0,0,0,107,0,133,0,4,0,245,0,209,0,177,0,243,0,105,0,234,0,28,0,0,0,87,0,0,0,224,0,153,0,45,0,45,0,161,0,207,0,210,0,191,0,0,0,33,0,48,0,0,0,136,0,143,0,241,0,61,0,175,0,133,0,214,0,253,0,0,0,157,0,218,0,0,0,66,0,119,0,0,0,44,0,14,0,40,0,211,0,187,0,18,0,0,0,56,0,208,0,0,0,208,0,101,0,0,0,132,0,135,0,195,0,82,0,0,0,0,0,18,0,36,0,93,0,0,0,59,0,134,0,147,0,0,0,0,0,168,0,0,0,237,0,0,0,45,0,44,0,0,0,241,0,132,0,0,0,133,0,95,0,190,0,78,0,191,0,0,0,98,0,108,0,181,0,74,0,143,0,24,0,151,0,219,0,58,0,109,0,216,0,0,0,60,0,191,0,104,0,57,0,59,0,103,0,38,0,193,0,66,0,124,0,113,0,5,0,0,0,185,0,241,0,198,0,125,0,19,0,0,0,133,0,157,0,0,0,187,0,107,0,224,0,51,0,0,0,50,0,167,0,21,0,158,0,211,0,0,0,0,0,3,0,246,0,0,0,104,0,240,0,0,0,32,0,5,0,118,0,246,0,237,0,219,0,39,0,56,0,166,0,0,0,239,0,45,0,48,0,180,0,108,0,189,0,143,0,61,0,16,0,178,0,3,0,92,0,39,0,46,0,199,0,0,0,0,0,0,0,30,0,0,0,0,0,208,0,94,0,0,0,214,0,87,0,155,0,177,0,0,0,111,0,215,0,0,0,0,0,137,0,99,0,175,0,55,0,129,0,251,0,94,0,23,0,103,0,147,0,79,0,0,0,190,0,0,0,188,0,114,0,13,0,215,0,104,0,144,0,0,0);
signal scenario_full  : scenario_type := (3,31,3,30,3,29,90,31,50,31,153,31,152,31,252,31,201,31,15,31,112,31,112,30,250,31,250,30,158,31,158,30,57,31,57,30,252,31,252,30,170,31,188,31,196,31,225,31,192,31,3,31,48,31,48,30,159,31,124,31,35,31,55,31,104,31,150,31,203,31,203,30,203,29,151,31,165,31,247,31,5,31,133,31,11,31,151,31,64,31,3,31,139,31,208,31,208,30,117,31,84,31,136,31,130,31,38,31,146,31,184,31,145,31,55,31,177,31,133,31,108,31,251,31,84,31,54,31,65,31,190,31,32,31,226,31,226,30,83,31,38,31,75,31,75,30,120,31,185,31,69,31,67,31,142,31,17,31,136,31,25,31,25,30,76,31,134,31,134,30,134,29,199,31,245,31,245,30,100,31,120,31,120,30,89,31,89,30,129,31,107,31,19,31,130,31,104,31,133,31,164,31,23,31,229,31,249,31,151,31,151,30,201,31,188,31,46,31,180,31,180,30,230,31,137,31,221,31,209,31,69,31,98,31,123,31,139,31,172,31,1,31,155,31,155,31,59,31,4,31,193,31,193,30,132,31,63,31,10,31,70,31,220,31,103,31,108,31,186,31,54,31,166,31,166,30,27,31,27,30,246,31,201,31,233,31,233,30,51,31,24,31,64,31,238,31,221,31,186,31,191,31,200,31,16,31,16,30,249,31,94,31,21,31,246,31,80,31,94,31,53,31,100,31,11,31,11,30,44,31,148,31,141,31,141,30,203,31,203,30,241,31,108,31,93,31,46,31,4,31,56,31,130,31,79,31,164,31,2,31,231,31,139,31,80,31,89,31,48,31,150,31,219,31,255,31,11,31,116,31,33,31,116,31,3,31,73,31,202,31,58,31,252,31,171,31,89,31,89,30,238,31,163,31,211,31,98,31,130,31,46,31,129,31,255,31,255,30,65,31,44,31,250,31,55,31,249,31,249,30,249,29,205,31,96,31,166,31,196,31,25,31,25,30,41,31,230,31,37,31,181,31,123,31,172,31,246,31,246,30,74,31,160,31,160,30,25,31,25,30,225,31,206,31,123,31,69,31,5,31,130,31,130,30,130,31,137,31,2,31,2,30,224,31,224,30,161,31,83,31,227,31,227,30,215,31,161,31,102,31,76,31,89,31,89,30,162,31,138,31,191,31,14,31,134,31,76,31,76,30,230,31,230,30,230,29,98,31,164,31,152,31,113,31,37,31,29,31,29,30,163,31,173,31,114,31,207,31,57,31,226,31,226,30,72,31,96,31,96,30,55,31,66,31,66,30,184,31,236,31,226,31,248,31,40,31,40,30,41,31,16,31,164,31,193,31,1,31,1,30,255,31,255,30,212,31,238,31,85,31,122,31,128,31,128,30,110,31,119,31,8,31,165,31,165,30,45,31,105,31,36,31,21,31,21,30,24,31,77,31,86,31,86,30,102,31,102,30,81,31,81,30,179,31,127,31,202,31,54,31,16,31,67,31,103,31,86,31,88,31,151,31,30,31,57,31,71,31,56,31,2,31,91,31,91,30,92,31,85,31,85,30,26,31,253,31,6,31,238,31,212,31,208,31,47,31,139,31,155,31,155,30,207,31,48,31,112,31,131,31,202,31,202,30,171,31,147,31,147,30,147,29,246,31,174,31,38,31,230,31,202,31,206,31,137,31,30,31,30,30,177,31,6,31,41,31,42,31,42,30,42,29,42,28,91,31,106,31,100,31,6,31,6,30,69,31,33,31,30,31,106,31,117,31,117,30,162,31,67,31,151,31,152,31,22,31,243,31,243,30,102,31,236,31,211,31,181,31,99,31,37,31,77,31,105,31,217,31,161,31,244,31,93,31,5,31,220,31,164,31,189,31,196,31,159,31,145,31,145,30,146,31,230,31,216,31,124,31,55,31,19,31,84,31,84,30,107,31,107,30,124,31,35,31,35,30,35,29,63,31,206,31,206,30,3,31,3,30,3,29,1,31,171,31,243,31,193,31,88,31,88,30,184,31,127,31,216,31,216,30,216,29,216,28,97,31,42,31,42,30,42,29,23,31,116,31,233,31,245,31,95,31,227,31,204,31,182,31,199,31,78,31,242,31,242,30,242,29,102,31,165,31,201,31,254,31,207,31,207,30,58,31,162,31,60,31,60,30,231,31,231,30,231,29,231,28,231,27,231,26,26,31,49,31,20,31,224,31,179,31,2,31,80,31,57,31,229,31,116,31,4,31,180,31,180,30,180,29,133,31,88,31,198,31,5,31,94,31,84,31,232,31,30,31,148,31,183,31,193,31,15,31,27,31,207,31,115,31,58,31,2,31,168,31,197,31,102,31,149,31,21,31,21,30,184,31,75,31,80,31,210,31,69,31,240,31,89,31,91,31,240,31,191,31,113,31,38,31,34,31,179,31,92,31,157,31,157,30,81,31,110,31,114,31,114,30,213,31,213,30,213,29,26,31,7,31,7,30,127,31,254,31,176,31,176,30,176,29,60,31,231,31,231,30,231,29,140,31,130,31,210,31,69,31,101,31,13,31,29,31,64,31,31,31,120,31,63,31,83,31,181,31,181,30,254,31,127,31,10,31,63,31,228,31,229,31,248,31,104,31,120,31,180,31,56,31,56,30,117,31,154,31,154,30,154,29,223,31,162,31,9,31,140,31,186,31,58,31,28,31,139,31,85,31,212,31,123,31,72,31,163,31,114,31,177,31,166,31,197,31,197,30,79,31,34,31,214,31,98,31,104,31,201,31,96,31,96,30,230,31,230,30,114,31,114,31,114,31,9,31,9,30,9,29,150,31,27,31,27,30,23,31,216,31,122,31,156,31,111,31,91,31,143,31,209,31,93,31,225,31,161,31,228,31,228,30,178,31,66,31,66,30,89,31,45,31,124,31,132,31,54,31,71,31,20,31,57,31,201,31,189,31,95,31,96,31,245,31,245,30,60,31,60,30,242,31,185,31,56,31,56,30,193,31,180,31,65,31,82,31,149,31,171,31,219,31,162,31,12,31,184,31,12,31,93,31,210,31,210,30,206,31,206,30,88,31,81,31,81,30,81,29,81,28,200,31,126,31,126,30,126,29,160,31,153,31,153,30,153,29,71,31,242,31,126,31,77,31,213,31,213,30,66,31,124,31,60,31,60,30,253,31,160,31,131,31,44,31,44,30,213,31,188,31,28,31,101,31,101,30,214,31,55,31,55,30,43,31,43,31,65,31,104,31,104,30,181,31,236,31,78,31,106,31,29,31,207,31,105,31,109,31,109,30,48,31,244,31,163,31,163,30,91,31,58,31,109,31,111,31,243,31,108,31,56,31,233,31,150,31,150,30,82,31,82,30,151,31,176,31,176,30,254,31,254,30,107,31,133,31,4,31,245,31,209,31,177,31,243,31,105,31,234,31,28,31,28,30,87,31,87,30,224,31,153,31,45,31,45,31,161,31,207,31,210,31,191,31,191,30,33,31,48,31,48,30,136,31,143,31,241,31,61,31,175,31,133,31,214,31,253,31,253,30,157,31,218,31,218,30,66,31,119,31,119,30,44,31,14,31,40,31,211,31,187,31,18,31,18,30,56,31,208,31,208,30,208,31,101,31,101,30,132,31,135,31,195,31,82,31,82,30,82,29,18,31,36,31,93,31,93,30,59,31,134,31,147,31,147,30,147,29,168,31,168,30,237,31,237,30,45,31,44,31,44,30,241,31,132,31,132,30,133,31,95,31,190,31,78,31,191,31,191,30,98,31,108,31,181,31,74,31,143,31,24,31,151,31,219,31,58,31,109,31,216,31,216,30,60,31,191,31,104,31,57,31,59,31,103,31,38,31,193,31,66,31,124,31,113,31,5,31,5,30,185,31,241,31,198,31,125,31,19,31,19,30,133,31,157,31,157,30,187,31,107,31,224,31,51,31,51,30,50,31,167,31,21,31,158,31,211,31,211,30,211,29,3,31,246,31,246,30,104,31,240,31,240,30,32,31,5,31,118,31,246,31,237,31,219,31,39,31,56,31,166,31,166,30,239,31,45,31,48,31,180,31,108,31,189,31,143,31,61,31,16,31,178,31,3,31,92,31,39,31,46,31,199,31,199,30,199,29,199,28,30,31,30,30,30,29,208,31,94,31,94,30,214,31,87,31,155,31,177,31,177,30,111,31,215,31,215,30,215,29,137,31,99,31,175,31,55,31,129,31,251,31,94,31,23,31,103,31,147,31,79,31,79,30,190,31,190,30,188,31,114,31,13,31,215,31,104,31,144,31,144,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
