-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 865;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (2,0,229,0,193,0,18,0,236,0,31,0,43,0,250,0,18,0,0,0,214,0,237,0,227,0,239,0,194,0,0,0,233,0,38,0,246,0,96,0,12,0,57,0,160,0,0,0,64,0,68,0,23,0,48,0,49,0,156,0,43,0,132,0,111,0,69,0,100,0,240,0,94,0,255,0,189,0,107,0,0,0,197,0,91,0,0,0,193,0,54,0,196,0,0,0,212,0,97,0,207,0,147,0,207,0,195,0,148,0,204,0,233,0,124,0,187,0,235,0,0,0,0,0,172,0,45,0,0,0,113,0,125,0,132,0,137,0,0,0,238,0,41,0,110,0,189,0,0,0,245,0,0,0,173,0,238,0,131,0,18,0,225,0,41,0,216,0,0,0,42,0,78,0,164,0,58,0,0,0,0,0,127,0,84,0,26,0,222,0,14,0,23,0,0,0,216,0,151,0,31,0,234,0,4,0,242,0,244,0,229,0,133,0,70,0,0,0,190,0,0,0,0,0,63,0,95,0,82,0,1,0,0,0,188,0,201,0,0,0,146,0,126,0,253,0,0,0,0,0,0,0,95,0,244,0,240,0,56,0,0,0,171,0,140,0,0,0,213,0,168,0,109,0,140,0,25,0,150,0,0,0,188,0,26,0,14,0,137,0,92,0,216,0,34,0,220,0,0,0,59,0,148,0,92,0,137,0,212,0,95,0,0,0,0,0,247,0,34,0,244,0,0,0,106,0,242,0,30,0,99,0,42,0,122,0,148,0,167,0,190,0,0,0,178,0,233,0,2,0,98,0,0,0,44,0,207,0,133,0,101,0,35,0,109,0,170,0,26,0,175,0,188,0,0,0,115,0,45,0,167,0,0,0,27,0,134,0,54,0,0,0,126,0,244,0,0,0,75,0,0,0,182,0,94,0,40,0,248,0,162,0,0,0,34,0,28,0,112,0,76,0,77,0,217,0,75,0,47,0,251,0,184,0,0,0,221,0,68,0,45,0,41,0,0,0,0,0,94,0,155,0,22,0,249,0,174,0,106,0,254,0,152,0,181,0,220,0,101,0,0,0,21,0,171,0,0,0,58,0,0,0,115,0,2,0,218,0,27,0,36,0,206,0,66,0,203,0,0,0,12,0,0,0,95,0,206,0,106,0,173,0,148,0,228,0,3,0,0,0,67,0,122,0,56,0,0,0,51,0,2,0,0,0,0,0,153,0,138,0,201,0,221,0,182,0,0,0,223,0,51,0,32,0,141,0,244,0,22,0,50,0,0,0,141,0,168,0,93,0,31,0,103,0,130,0,126,0,2,0,158,0,24,0,0,0,70,0,164,0,49,0,197,0,131,0,0,0,93,0,159,0,13,0,0,0,207,0,0,0,222,0,125,0,63,0,79,0,166,0,203,0,164,0,220,0,185,0,99,0,115,0,74,0,240,0,223,0,3,0,0,0,251,0,0,0,8,0,115,0,0,0,44,0,174,0,51,0,217,0,123,0,0,0,177,0,43,0,169,0,73,0,100,0,113,0,0,0,170,0,181,0,0,0,237,0,187,0,221,0,0,0,35,0,220,0,0,0,174,0,141,0,14,0,217,0,10,0,176,0,79,0,3,0,0,0,27,0,0,0,41,0,209,0,84,0,51,0,5,0,21,0,84,0,148,0,183,0,0,0,172,0,204,0,0,0,108,0,225,0,194,0,95,0,0,0,0,0,118,0,207,0,70,0,205,0,0,0,0,0,0,0,0,0,0,0,196,0,78,0,167,0,84,0,0,0,190,0,168,0,0,0,211,0,120,0,0,0,42,0,0,0,238,0,51,0,173,0,0,0,59,0,166,0,83,0,251,0,221,0,47,0,200,0,0,0,107,0,23,0,185,0,138,0,163,0,145,0,12,0,171,0,0,0,198,0,149,0,187,0,0,0,0,0,59,0,10,0,218,0,101,0,0,0,38,0,65,0,212,0,113,0,164,0,0,0,76,0,76,0,103,0,177,0,74,0,192,0,0,0,230,0,80,0,211,0,164,0,204,0,214,0,31,0,186,0,245,0,172,0,182,0,113,0,55,0,245,0,75,0,156,0,176,0,167,0,172,0,5,0,72,0,211,0,125,0,18,0,254,0,121,0,175,0,215,0,199,0,63,0,168,0,231,0,0,0,86,0,107,0,178,0,0,0,63,0,0,0,68,0,175,0,110,0,177,0,104,0,220,0,25,0,85,0,197,0,238,0,0,0,0,0,14,0,0,0,118,0,37,0,119,0,148,0,183,0,197,0,23,0,86,0,137,0,73,0,88,0,120,0,0,0,172,0,21,0,130,0,0,0,175,0,231,0,126,0,150,0,209,0,145,0,204,0,0,0,0,0,117,0,0,0,78,0,0,0,223,0,134,0,58,0,105,0,154,0,216,0,68,0,0,0,57,0,254,0,26,0,91,0,62,0,0,0,0,0,124,0,224,0,127,0,127,0,85,0,71,0,27,0,209,0,0,0,51,0,178,0,40,0,178,0,173,0,120,0,0,0,11,0,101,0,0,0,123,0,152,0,75,0,121,0,0,0,226,0,104,0,183,0,46,0,95,0,228,0,0,0,1,0,0,0,88,0,80,0,6,0,114,0,0,0,192,0,147,0,150,0,80,0,177,0,179,0,99,0,8,0,101,0,0,0,144,0,129,0,101,0,29,0,190,0,0,0,0,0,169,0,139,0,8,0,104,0,199,0,109,0,0,0,136,0,46,0,92,0,10,0,201,0,43,0,19,0,11,0,40,0,0,0,27,0,175,0,139,0,0,0,91,0,7,0,170,0,93,0,147,0,59,0,0,0,198,0,89,0,222,0,42,0,196,0,72,0,0,0,246,0,51,0,0,0,43,0,0,0,0,0,34,0,163,0,215,0,0,0,126,0,138,0,181,0,176,0,0,0,255,0,243,0,156,0,141,0,84,0,122,0,0,0,34,0,0,0,235,0,117,0,98,0,200,0,0,0,0,0,100,0,115,0,0,0,0,0,51,0,66,0,94,0,228,0,0,0,126,0,0,0,27,0,9,0,210,0,74,0,145,0,102,0,188,0,131,0,178,0,0,0,16,0,41,0,213,0,3,0,67,0,3,0,97,0,2,0,206,0,190,0,136,0,105,0,0,0,45,0,117,0,245,0,152,0,211,0,174,0,223,0,20,0,130,0,223,0,249,0,95,0,169,0,233,0,29,0,217,0,137,0,97,0,83,0,0,0,13,0,86,0,117,0,89,0,0,0,127,0,0,0,246,0,0,0,158,0,87,0,0,0,140,0,83,0,0,0,0,0,8,0,18,0,0,0,191,0,227,0,0,0,0,0,35,0,0,0,35,0,6,0,0,0,176,0,216,0,31,0,0,0,0,0,13,0,27,0,148,0,54,0,238,0,236,0,179,0,130,0,226,0,113,0,23,0,108,0,226,0,77,0,168,0,21,0,227,0,219,0,0,0,135,0,120,0,81,0,61,0,0,0,32,0,102,0,125,0,100,0,0,0,18,0,128,0,86,0,165,0,59,0,208,0,98,0,208,0,62,0,23,0,106,0,0,0,128,0,251,0,30,0,220,0,0,0,53,0,164,0,251,0,175,0,201,0,244,0,0,0,12,0,0,0,192,0,81,0,0,0,60,0,252,0,215,0,210,0,0,0,255,0,15,0,88,0,0,0,213,0,16,0,228,0,122,0,114,0,0,0,0,0,167,0,86,0,3,0,176,0,234,0,148,0,241,0,241,0,187,0,0,0,230,0,124,0,13,0,22,0,105,0,148,0,177,0,165,0,19,0,116,0,141,0,174,0,191,0,5,0,0,0,90,0,58,0,54,0,251,0,110,0,211,0,229,0,230,0,0,0,92,0,212,0,173,0,136,0,0,0,0,0,230,0);
signal scenario_full  : scenario_type := (2,31,229,31,193,31,18,31,236,31,31,31,43,31,250,31,18,31,18,30,214,31,237,31,227,31,239,31,194,31,194,30,233,31,38,31,246,31,96,31,12,31,57,31,160,31,160,30,64,31,68,31,23,31,48,31,49,31,156,31,43,31,132,31,111,31,69,31,100,31,240,31,94,31,255,31,189,31,107,31,107,30,197,31,91,31,91,30,193,31,54,31,196,31,196,30,212,31,97,31,207,31,147,31,207,31,195,31,148,31,204,31,233,31,124,31,187,31,235,31,235,30,235,29,172,31,45,31,45,30,113,31,125,31,132,31,137,31,137,30,238,31,41,31,110,31,189,31,189,30,245,31,245,30,173,31,238,31,131,31,18,31,225,31,41,31,216,31,216,30,42,31,78,31,164,31,58,31,58,30,58,29,127,31,84,31,26,31,222,31,14,31,23,31,23,30,216,31,151,31,31,31,234,31,4,31,242,31,244,31,229,31,133,31,70,31,70,30,190,31,190,30,190,29,63,31,95,31,82,31,1,31,1,30,188,31,201,31,201,30,146,31,126,31,253,31,253,30,253,29,253,28,95,31,244,31,240,31,56,31,56,30,171,31,140,31,140,30,213,31,168,31,109,31,140,31,25,31,150,31,150,30,188,31,26,31,14,31,137,31,92,31,216,31,34,31,220,31,220,30,59,31,148,31,92,31,137,31,212,31,95,31,95,30,95,29,247,31,34,31,244,31,244,30,106,31,242,31,30,31,99,31,42,31,122,31,148,31,167,31,190,31,190,30,178,31,233,31,2,31,98,31,98,30,44,31,207,31,133,31,101,31,35,31,109,31,170,31,26,31,175,31,188,31,188,30,115,31,45,31,167,31,167,30,27,31,134,31,54,31,54,30,126,31,244,31,244,30,75,31,75,30,182,31,94,31,40,31,248,31,162,31,162,30,34,31,28,31,112,31,76,31,77,31,217,31,75,31,47,31,251,31,184,31,184,30,221,31,68,31,45,31,41,31,41,30,41,29,94,31,155,31,22,31,249,31,174,31,106,31,254,31,152,31,181,31,220,31,101,31,101,30,21,31,171,31,171,30,58,31,58,30,115,31,2,31,218,31,27,31,36,31,206,31,66,31,203,31,203,30,12,31,12,30,95,31,206,31,106,31,173,31,148,31,228,31,3,31,3,30,67,31,122,31,56,31,56,30,51,31,2,31,2,30,2,29,153,31,138,31,201,31,221,31,182,31,182,30,223,31,51,31,32,31,141,31,244,31,22,31,50,31,50,30,141,31,168,31,93,31,31,31,103,31,130,31,126,31,2,31,158,31,24,31,24,30,70,31,164,31,49,31,197,31,131,31,131,30,93,31,159,31,13,31,13,30,207,31,207,30,222,31,125,31,63,31,79,31,166,31,203,31,164,31,220,31,185,31,99,31,115,31,74,31,240,31,223,31,3,31,3,30,251,31,251,30,8,31,115,31,115,30,44,31,174,31,51,31,217,31,123,31,123,30,177,31,43,31,169,31,73,31,100,31,113,31,113,30,170,31,181,31,181,30,237,31,187,31,221,31,221,30,35,31,220,31,220,30,174,31,141,31,14,31,217,31,10,31,176,31,79,31,3,31,3,30,27,31,27,30,41,31,209,31,84,31,51,31,5,31,21,31,84,31,148,31,183,31,183,30,172,31,204,31,204,30,108,31,225,31,194,31,95,31,95,30,95,29,118,31,207,31,70,31,205,31,205,30,205,29,205,28,205,27,205,26,196,31,78,31,167,31,84,31,84,30,190,31,168,31,168,30,211,31,120,31,120,30,42,31,42,30,238,31,51,31,173,31,173,30,59,31,166,31,83,31,251,31,221,31,47,31,200,31,200,30,107,31,23,31,185,31,138,31,163,31,145,31,12,31,171,31,171,30,198,31,149,31,187,31,187,30,187,29,59,31,10,31,218,31,101,31,101,30,38,31,65,31,212,31,113,31,164,31,164,30,76,31,76,31,103,31,177,31,74,31,192,31,192,30,230,31,80,31,211,31,164,31,204,31,214,31,31,31,186,31,245,31,172,31,182,31,113,31,55,31,245,31,75,31,156,31,176,31,167,31,172,31,5,31,72,31,211,31,125,31,18,31,254,31,121,31,175,31,215,31,199,31,63,31,168,31,231,31,231,30,86,31,107,31,178,31,178,30,63,31,63,30,68,31,175,31,110,31,177,31,104,31,220,31,25,31,85,31,197,31,238,31,238,30,238,29,14,31,14,30,118,31,37,31,119,31,148,31,183,31,197,31,23,31,86,31,137,31,73,31,88,31,120,31,120,30,172,31,21,31,130,31,130,30,175,31,231,31,126,31,150,31,209,31,145,31,204,31,204,30,204,29,117,31,117,30,78,31,78,30,223,31,134,31,58,31,105,31,154,31,216,31,68,31,68,30,57,31,254,31,26,31,91,31,62,31,62,30,62,29,124,31,224,31,127,31,127,31,85,31,71,31,27,31,209,31,209,30,51,31,178,31,40,31,178,31,173,31,120,31,120,30,11,31,101,31,101,30,123,31,152,31,75,31,121,31,121,30,226,31,104,31,183,31,46,31,95,31,228,31,228,30,1,31,1,30,88,31,80,31,6,31,114,31,114,30,192,31,147,31,150,31,80,31,177,31,179,31,99,31,8,31,101,31,101,30,144,31,129,31,101,31,29,31,190,31,190,30,190,29,169,31,139,31,8,31,104,31,199,31,109,31,109,30,136,31,46,31,92,31,10,31,201,31,43,31,19,31,11,31,40,31,40,30,27,31,175,31,139,31,139,30,91,31,7,31,170,31,93,31,147,31,59,31,59,30,198,31,89,31,222,31,42,31,196,31,72,31,72,30,246,31,51,31,51,30,43,31,43,30,43,29,34,31,163,31,215,31,215,30,126,31,138,31,181,31,176,31,176,30,255,31,243,31,156,31,141,31,84,31,122,31,122,30,34,31,34,30,235,31,117,31,98,31,200,31,200,30,200,29,100,31,115,31,115,30,115,29,51,31,66,31,94,31,228,31,228,30,126,31,126,30,27,31,9,31,210,31,74,31,145,31,102,31,188,31,131,31,178,31,178,30,16,31,41,31,213,31,3,31,67,31,3,31,97,31,2,31,206,31,190,31,136,31,105,31,105,30,45,31,117,31,245,31,152,31,211,31,174,31,223,31,20,31,130,31,223,31,249,31,95,31,169,31,233,31,29,31,217,31,137,31,97,31,83,31,83,30,13,31,86,31,117,31,89,31,89,30,127,31,127,30,246,31,246,30,158,31,87,31,87,30,140,31,83,31,83,30,83,29,8,31,18,31,18,30,191,31,227,31,227,30,227,29,35,31,35,30,35,31,6,31,6,30,176,31,216,31,31,31,31,30,31,29,13,31,27,31,148,31,54,31,238,31,236,31,179,31,130,31,226,31,113,31,23,31,108,31,226,31,77,31,168,31,21,31,227,31,219,31,219,30,135,31,120,31,81,31,61,31,61,30,32,31,102,31,125,31,100,31,100,30,18,31,128,31,86,31,165,31,59,31,208,31,98,31,208,31,62,31,23,31,106,31,106,30,128,31,251,31,30,31,220,31,220,30,53,31,164,31,251,31,175,31,201,31,244,31,244,30,12,31,12,30,192,31,81,31,81,30,60,31,252,31,215,31,210,31,210,30,255,31,15,31,88,31,88,30,213,31,16,31,228,31,122,31,114,31,114,30,114,29,167,31,86,31,3,31,176,31,234,31,148,31,241,31,241,31,187,31,187,30,230,31,124,31,13,31,22,31,105,31,148,31,177,31,165,31,19,31,116,31,141,31,174,31,191,31,5,31,5,30,90,31,58,31,54,31,251,31,110,31,211,31,229,31,230,31,230,30,92,31,212,31,173,31,136,31,136,30,136,29,230,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
