-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 700;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (173,0,0,0,82,0,172,0,171,0,0,0,185,0,77,0,135,0,0,0,47,0,183,0,77,0,14,0,80,0,106,0,33,0,0,0,178,0,0,0,0,0,45,0,170,0,239,0,7,0,153,0,0,0,0,0,186,0,96,0,136,0,0,0,225,0,245,0,0,0,61,0,152,0,0,0,1,0,66,0,148,0,119,0,131,0,210,0,0,0,164,0,112,0,237,0,222,0,251,0,146,0,35,0,90,0,247,0,0,0,91,0,107,0,71,0,47,0,223,0,84,0,4,0,0,0,16,0,0,0,42,0,144,0,65,0,170,0,127,0,242,0,194,0,0,0,89,0,77,0,114,0,0,0,18,0,222,0,0,0,184,0,0,0,7,0,0,0,220,0,0,0,132,0,0,0,221,0,140,0,249,0,123,0,25,0,239,0,14,0,189,0,241,0,29,0,0,0,0,0,233,0,90,0,253,0,89,0,101,0,0,0,254,0,0,0,25,0,0,0,184,0,70,0,192,0,239,0,17,0,249,0,124,0,227,0,217,0,0,0,0,0,0,0,194,0,19,0,45,0,181,0,76,0,208,0,104,0,133,0,46,0,0,0,54,0,0,0,56,0,176,0,120,0,37,0,0,0,35,0,154,0,204,0,204,0,70,0,109,0,195,0,220,0,254,0,0,0,236,0,115,0,110,0,0,0,0,0,173,0,209,0,155,0,107,0,0,0,198,0,0,0,3,0,190,0,96,0,107,0,209,0,114,0,225,0,162,0,13,0,200,0,201,0,246,0,252,0,105,0,1,0,185,0,0,0,136,0,168,0,0,0,0,0,29,0,0,0,181,0,223,0,159,0,228,0,0,0,243,0,122,0,66,0,218,0,52,0,50,0,244,0,0,0,0,0,173,0,89,0,0,0,34,0,0,0,0,0,0,0,64,0,55,0,2,0,0,0,149,0,19,0,196,0,184,0,24,0,132,0,0,0,23,0,23,0,255,0,81,0,80,0,29,0,169,0,31,0,103,0,239,0,138,0,0,0,162,0,54,0,72,0,7,0,110,0,0,0,54,0,0,0,1,0,110,0,116,0,152,0,35,0,34,0,0,0,143,0,10,0,150,0,43,0,242,0,27,0,0,0,73,0,0,0,243,0,117,0,254,0,0,0,45,0,136,0,110,0,41,0,108,0,0,0,144,0,114,0,92,0,181,0,187,0,155,0,118,0,51,0,238,0,0,0,160,0,203,0,212,0,0,0,141,0,216,0,0,0,132,0,19,0,51,0,0,0,0,0,229,0,131,0,223,0,53,0,190,0,115,0,0,0,0,0,252,0,58,0,222,0,69,0,240,0,229,0,238,0,0,0,0,0,0,0,220,0,144,0,148,0,0,0,232,0,237,0,112,0,0,0,0,0,145,0,0,0,92,0,0,0,106,0,157,0,0,0,182,0,0,0,0,0,0,0,246,0,172,0,147,0,143,0,73,0,117,0,22,0,158,0,137,0,0,0,187,0,147,0,119,0,77,0,0,0,181,0,89,0,0,0,39,0,194,0,77,0,26,0,159,0,128,0,67,0,107,0,142,0,208,0,232,0,32,0,17,0,48,0,117,0,0,0,229,0,0,0,89,0,95,0,140,0,216,0,160,0,67,0,211,0,6,0,215,0,168,0,131,0,50,0,164,0,88,0,184,0,255,0,38,0,0,0,170,0,10,0,142,0,101,0,11,0,138,0,203,0,159,0,202,0,0,0,0,0,167,0,42,0,1,0,71,0,0,0,232,0,0,0,35,0,96,0,140,0,42,0,8,0,0,0,159,0,0,0,0,0,77,0,255,0,95,0,182,0,46,0,200,0,68,0,0,0,206,0,114,0,41,0,0,0,121,0,138,0,153,0,90,0,0,0,20,0,128,0,0,0,251,0,30,0,1,0,207,0,0,0,0,0,241,0,0,0,188,0,94,0,250,0,186,0,18,0,22,0,224,0,25,0,233,0,74,0,131,0,0,0,202,0,36,0,113,0,248,0,115,0,113,0,28,0,177,0,203,0,31,0,51,0,78,0,10,0,38,0,167,0,64,0,128,0,136,0,0,0,191,0,133,0,217,0,0,0,142,0,0,0,247,0,0,0,49,0,0,0,131,0,254,0,37,0,248,0,32,0,69,0,74,0,57,0,32,0,227,0,228,0,168,0,52,0,0,0,0,0,2,0,80,0,108,0,38,0,0,0,161,0,204,0,184,0,156,0,34,0,115,0,0,0,0,0,214,0,0,0,15,0,0,0,253,0,20,0,254,0,22,0,247,0,0,0,247,0,30,0,74,0,146,0,76,0,170,0,127,0,0,0,217,0,8,0,134,0,0,0,0,0,0,0,44,0,69,0,196,0,39,0,38,0,0,0,234,0,50,0,150,0,3,0,210,0,0,0,17,0,22,0,135,0,253,0,46,0,68,0,66,0,61,0,0,0,222,0,0,0,1,0,238,0,209,0,0,0,188,0,164,0,219,0,215,0,101,0,101,0,0,0,22,0,91,0,55,0,0,0,205,0,41,0,191,0,0,0,130,0,45,0,249,0,0,0,0,0,0,0,176,0,209,0,23,0,186,0,151,0,0,0,0,0,0,0,190,0,43,0,236,0,6,0,128,0,13,0,170,0,122,0,111,0,42,0,0,0,72,0,153,0,244,0,184,0,96,0,79,0,101,0,111,0,16,0,30,0,242,0,17,0,0,0,229,0,0,0,208,0,111,0,98,0,252,0,182,0,0,0,180,0,199,0,0,0,126,0,32,0,12,0,0,0,217,0,0,0,16,0,40,0,215,0,71,0,25,0,71,0,155,0,166,0,180,0,240,0,0,0,194,0,56,0,0,0,146,0,110,0,23,0,129,0,0,0,214,0,8,0,21,0,169,0,0,0,60,0,124,0,0,0,41,0,205,0,152,0,0,0,239,0,50,0,50,0,167,0,150,0,0,0,0,0,0,0,2,0,216,0,138,0,121,0,104,0,37,0,248,0,174,0,38,0,3,0,18,0,0,0,7,0,0,0,250,0,114,0,27,0,77,0,109,0,242,0,0,0,161,0,12,0,0,0,0,0,201,0,148,0,0,0,0,0,219,0,0,0,5,0,130,0,0,0,100,0,198,0,215,0,151,0,240,0,172,0);
signal scenario_full  : scenario_type := (173,31,173,30,82,31,172,31,171,31,171,30,185,31,77,31,135,31,135,30,47,31,183,31,77,31,14,31,80,31,106,31,33,31,33,30,178,31,178,30,178,29,45,31,170,31,239,31,7,31,153,31,153,30,153,29,186,31,96,31,136,31,136,30,225,31,245,31,245,30,61,31,152,31,152,30,1,31,66,31,148,31,119,31,131,31,210,31,210,30,164,31,112,31,237,31,222,31,251,31,146,31,35,31,90,31,247,31,247,30,91,31,107,31,71,31,47,31,223,31,84,31,4,31,4,30,16,31,16,30,42,31,144,31,65,31,170,31,127,31,242,31,194,31,194,30,89,31,77,31,114,31,114,30,18,31,222,31,222,30,184,31,184,30,7,31,7,30,220,31,220,30,132,31,132,30,221,31,140,31,249,31,123,31,25,31,239,31,14,31,189,31,241,31,29,31,29,30,29,29,233,31,90,31,253,31,89,31,101,31,101,30,254,31,254,30,25,31,25,30,184,31,70,31,192,31,239,31,17,31,249,31,124,31,227,31,217,31,217,30,217,29,217,28,194,31,19,31,45,31,181,31,76,31,208,31,104,31,133,31,46,31,46,30,54,31,54,30,56,31,176,31,120,31,37,31,37,30,35,31,154,31,204,31,204,31,70,31,109,31,195,31,220,31,254,31,254,30,236,31,115,31,110,31,110,30,110,29,173,31,209,31,155,31,107,31,107,30,198,31,198,30,3,31,190,31,96,31,107,31,209,31,114,31,225,31,162,31,13,31,200,31,201,31,246,31,252,31,105,31,1,31,185,31,185,30,136,31,168,31,168,30,168,29,29,31,29,30,181,31,223,31,159,31,228,31,228,30,243,31,122,31,66,31,218,31,52,31,50,31,244,31,244,30,244,29,173,31,89,31,89,30,34,31,34,30,34,29,34,28,64,31,55,31,2,31,2,30,149,31,19,31,196,31,184,31,24,31,132,31,132,30,23,31,23,31,255,31,81,31,80,31,29,31,169,31,31,31,103,31,239,31,138,31,138,30,162,31,54,31,72,31,7,31,110,31,110,30,54,31,54,30,1,31,110,31,116,31,152,31,35,31,34,31,34,30,143,31,10,31,150,31,43,31,242,31,27,31,27,30,73,31,73,30,243,31,117,31,254,31,254,30,45,31,136,31,110,31,41,31,108,31,108,30,144,31,114,31,92,31,181,31,187,31,155,31,118,31,51,31,238,31,238,30,160,31,203,31,212,31,212,30,141,31,216,31,216,30,132,31,19,31,51,31,51,30,51,29,229,31,131,31,223,31,53,31,190,31,115,31,115,30,115,29,252,31,58,31,222,31,69,31,240,31,229,31,238,31,238,30,238,29,238,28,220,31,144,31,148,31,148,30,232,31,237,31,112,31,112,30,112,29,145,31,145,30,92,31,92,30,106,31,157,31,157,30,182,31,182,30,182,29,182,28,246,31,172,31,147,31,143,31,73,31,117,31,22,31,158,31,137,31,137,30,187,31,147,31,119,31,77,31,77,30,181,31,89,31,89,30,39,31,194,31,77,31,26,31,159,31,128,31,67,31,107,31,142,31,208,31,232,31,32,31,17,31,48,31,117,31,117,30,229,31,229,30,89,31,95,31,140,31,216,31,160,31,67,31,211,31,6,31,215,31,168,31,131,31,50,31,164,31,88,31,184,31,255,31,38,31,38,30,170,31,10,31,142,31,101,31,11,31,138,31,203,31,159,31,202,31,202,30,202,29,167,31,42,31,1,31,71,31,71,30,232,31,232,30,35,31,96,31,140,31,42,31,8,31,8,30,159,31,159,30,159,29,77,31,255,31,95,31,182,31,46,31,200,31,68,31,68,30,206,31,114,31,41,31,41,30,121,31,138,31,153,31,90,31,90,30,20,31,128,31,128,30,251,31,30,31,1,31,207,31,207,30,207,29,241,31,241,30,188,31,94,31,250,31,186,31,18,31,22,31,224,31,25,31,233,31,74,31,131,31,131,30,202,31,36,31,113,31,248,31,115,31,113,31,28,31,177,31,203,31,31,31,51,31,78,31,10,31,38,31,167,31,64,31,128,31,136,31,136,30,191,31,133,31,217,31,217,30,142,31,142,30,247,31,247,30,49,31,49,30,131,31,254,31,37,31,248,31,32,31,69,31,74,31,57,31,32,31,227,31,228,31,168,31,52,31,52,30,52,29,2,31,80,31,108,31,38,31,38,30,161,31,204,31,184,31,156,31,34,31,115,31,115,30,115,29,214,31,214,30,15,31,15,30,253,31,20,31,254,31,22,31,247,31,247,30,247,31,30,31,74,31,146,31,76,31,170,31,127,31,127,30,217,31,8,31,134,31,134,30,134,29,134,28,44,31,69,31,196,31,39,31,38,31,38,30,234,31,50,31,150,31,3,31,210,31,210,30,17,31,22,31,135,31,253,31,46,31,68,31,66,31,61,31,61,30,222,31,222,30,1,31,238,31,209,31,209,30,188,31,164,31,219,31,215,31,101,31,101,31,101,30,22,31,91,31,55,31,55,30,205,31,41,31,191,31,191,30,130,31,45,31,249,31,249,30,249,29,249,28,176,31,209,31,23,31,186,31,151,31,151,30,151,29,151,28,190,31,43,31,236,31,6,31,128,31,13,31,170,31,122,31,111,31,42,31,42,30,72,31,153,31,244,31,184,31,96,31,79,31,101,31,111,31,16,31,30,31,242,31,17,31,17,30,229,31,229,30,208,31,111,31,98,31,252,31,182,31,182,30,180,31,199,31,199,30,126,31,32,31,12,31,12,30,217,31,217,30,16,31,40,31,215,31,71,31,25,31,71,31,155,31,166,31,180,31,240,31,240,30,194,31,56,31,56,30,146,31,110,31,23,31,129,31,129,30,214,31,8,31,21,31,169,31,169,30,60,31,124,31,124,30,41,31,205,31,152,31,152,30,239,31,50,31,50,31,167,31,150,31,150,30,150,29,150,28,2,31,216,31,138,31,121,31,104,31,37,31,248,31,174,31,38,31,3,31,18,31,18,30,7,31,7,30,250,31,114,31,27,31,77,31,109,31,242,31,242,30,161,31,12,31,12,30,12,29,201,31,148,31,148,30,148,29,219,31,219,30,5,31,130,31,130,30,100,31,198,31,215,31,151,31,240,31,172,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
