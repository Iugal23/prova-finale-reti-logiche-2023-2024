-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 644;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (64,0,107,0,0,0,4,0,0,0,254,0,155,0,212,0,136,0,147,0,155,0,0,0,210,0,107,0,217,0,10,0,0,0,139,0,60,0,11,0,0,0,210,0,192,0,7,0,219,0,89,0,2,0,244,0,0,0,0,0,182,0,178,0,41,0,213,0,237,0,64,0,99,0,58,0,56,0,0,0,152,0,130,0,229,0,214,0,0,0,38,0,93,0,240,0,0,0,0,0,0,0,84,0,0,0,0,0,240,0,45,0,0,0,6,0,221,0,175,0,74,0,107,0,17,0,35,0,114,0,0,0,28,0,3,0,157,0,0,0,198,0,186,0,36,0,232,0,198,0,162,0,78,0,108,0,229,0,247,0,120,0,187,0,76,0,0,0,122,0,102,0,106,0,132,0,3,0,27,0,105,0,81,0,142,0,68,0,41,0,16,0,120,0,200,0,167,0,129,0,0,0,251,0,67,0,43,0,0,0,238,0,0,0,176,0,200,0,0,0,170,0,0,0,21,0,248,0,97,0,185,0,19,0,0,0,157,0,9,0,20,0,83,0,164,0,255,0,96,0,175,0,211,0,84,0,60,0,161,0,12,0,206,0,98,0,233,0,46,0,104,0,11,0,58,0,160,0,0,0,0,0,1,0,0,0,196,0,0,0,211,0,0,0,0,0,0,0,185,0,131,0,61,0,117,0,32,0,110,0,248,0,217,0,0,0,16,0,1,0,0,0,0,0,198,0,1,0,250,0,197,0,243,0,0,0,0,0,104,0,135,0,233,0,75,0,0,0,52,0,65,0,224,0,0,0,34,0,228,0,244,0,90,0,94,0,69,0,20,0,0,0,0,0,226,0,59,0,91,0,181,0,16,0,216,0,161,0,241,0,78,0,0,0,0,0,251,0,178,0,9,0,94,0,4,0,0,0,0,0,117,0,201,0,141,0,110,0,0,0,49,0,60,0,220,0,193,0,36,0,70,0,170,0,171,0,84,0,0,0,0,0,69,0,143,0,76,0,52,0,252,0,130,0,34,0,241,0,0,0,187,0,206,0,0,0,0,0,96,0,253,0,0,0,250,0,199,0,233,0,169,0,252,0,71,0,0,0,0,0,0,0,166,0,5,0,119,0,162,0,108,0,162,0,110,0,157,0,0,0,180,0,212,0,0,0,40,0,251,0,13,0,160,0,130,0,165,0,157,0,0,0,247,0,0,0,237,0,188,0,30,0,115,0,128,0,232,0,216,0,56,0,0,0,69,0,0,0,0,0,156,0,152,0,163,0,110,0,0,0,0,0,178,0,102,0,232,0,231,0,220,0,232,0,148,0,131,0,16,0,4,0,205,0,21,0,227,0,51,0,0,0,15,0,182,0,137,0,108,0,0,0,157,0,225,0,221,0,246,0,0,0,189,0,233,0,90,0,0,0,0,0,157,0,0,0,178,0,243,0,0,0,114,0,0,0,60,0,223,0,246,0,182,0,0,0,113,0,112,0,68,0,0,0,23,0,1,0,232,0,102,0,79,0,141,0,55,0,171,0,208,0,230,0,177,0,235,0,11,0,168,0,119,0,177,0,198,0,209,0,74,0,0,0,0,0,179,0,111,0,0,0,137,0,32,0,22,0,99,0,201,0,0,0,236,0,211,0,3,0,6,0,221,0,121,0,134,0,0,0,176,0,19,0,115,0,246,0,0,0,0,0,222,0,0,0,160,0,0,0,192,0,218,0,52,0,2,0,64,0,27,0,0,0,0,0,0,0,114,0,91,0,129,0,236,0,49,0,67,0,85,0,0,0,196,0,4,0,0,0,41,0,0,0,0,0,228,0,0,0,206,0,228,0,177,0,181,0,35,0,100,0,245,0,0,0,73,0,17,0,0,0,20,0,239,0,251,0,96,0,29,0,0,0,155,0,68,0,63,0,141,0,9,0,7,0,77,0,0,0,75,0,104,0,0,0,205,0,143,0,132,0,0,0,48,0,0,0,54,0,100,0,210,0,37,0,0,0,75,0,49,0,137,0,254,0,132,0,169,0,239,0,247,0,0,0,69,0,26,0,22,0,159,0,236,0,53,0,24,0,220,0,54,0,120,0,139,0,29,0,66,0,0,0,112,0,0,0,213,0,0,0,0,0,39,0,35,0,136,0,0,0,0,0,198,0,0,0,193,0,22,0,208,0,0,0,57,0,188,0,7,0,180,0,81,0,139,0,102,0,0,0,194,0,224,0,53,0,38,0,231,0,194,0,0,0,220,0,0,0,221,0,0,0,152,0,67,0,172,0,6,0,52,0,118,0,79,0,236,0,57,0,244,0,194,0,51,0,135,0,69,0,3,0,0,0,0,0,79,0,214,0,0,0,126,0,118,0,97,0,0,0,30,0,0,0,207,0,80,0,0,0,132,0,199,0,79,0,134,0,5,0,206,0,19,0,245,0,87,0,23,0,226,0,39,0,162,0,81,0,0,0,142,0,109,0,180,0,204,0,101,0,42,0,159,0,26,0,131,0,120,0,0,0,138,0,0,0,140,0,0,0,0,0,98,0,73,0,199,0,245,0,140,0,232,0,26,0,131,0,0,0,0,0,3,0,176,0,0,0,0,0,199,0,92,0,179,0,154,0,252,0,140,0,177,0,0,0,255,0,0,0,161,0,0,0,58,0,0,0,221,0,174,0,203,0,52,0,0,0,217,0,69,0,127,0,233,0,90,0,17,0,248,0,54,0,238,0,122,0,0,0,219,0,0,0,38,0,235,0,229,0,0,0,173,0,252,0,62,0,0,0,210,0,0,0,36,0,125,0,138,0,0,0,70,0,0,0,0,0,129,0,47,0,212,0,12,0,0,0,119,0,96,0,71,0,175,0,190,0,0,0,68,0,32,0,0,0,22,0,221,0,26,0,248,0,235,0);
signal scenario_full  : scenario_type := (64,31,107,31,107,30,4,31,4,30,254,31,155,31,212,31,136,31,147,31,155,31,155,30,210,31,107,31,217,31,10,31,10,30,139,31,60,31,11,31,11,30,210,31,192,31,7,31,219,31,89,31,2,31,244,31,244,30,244,29,182,31,178,31,41,31,213,31,237,31,64,31,99,31,58,31,56,31,56,30,152,31,130,31,229,31,214,31,214,30,38,31,93,31,240,31,240,30,240,29,240,28,84,31,84,30,84,29,240,31,45,31,45,30,6,31,221,31,175,31,74,31,107,31,17,31,35,31,114,31,114,30,28,31,3,31,157,31,157,30,198,31,186,31,36,31,232,31,198,31,162,31,78,31,108,31,229,31,247,31,120,31,187,31,76,31,76,30,122,31,102,31,106,31,132,31,3,31,27,31,105,31,81,31,142,31,68,31,41,31,16,31,120,31,200,31,167,31,129,31,129,30,251,31,67,31,43,31,43,30,238,31,238,30,176,31,200,31,200,30,170,31,170,30,21,31,248,31,97,31,185,31,19,31,19,30,157,31,9,31,20,31,83,31,164,31,255,31,96,31,175,31,211,31,84,31,60,31,161,31,12,31,206,31,98,31,233,31,46,31,104,31,11,31,58,31,160,31,160,30,160,29,1,31,1,30,196,31,196,30,211,31,211,30,211,29,211,28,185,31,131,31,61,31,117,31,32,31,110,31,248,31,217,31,217,30,16,31,1,31,1,30,1,29,198,31,1,31,250,31,197,31,243,31,243,30,243,29,104,31,135,31,233,31,75,31,75,30,52,31,65,31,224,31,224,30,34,31,228,31,244,31,90,31,94,31,69,31,20,31,20,30,20,29,226,31,59,31,91,31,181,31,16,31,216,31,161,31,241,31,78,31,78,30,78,29,251,31,178,31,9,31,94,31,4,31,4,30,4,29,117,31,201,31,141,31,110,31,110,30,49,31,60,31,220,31,193,31,36,31,70,31,170,31,171,31,84,31,84,30,84,29,69,31,143,31,76,31,52,31,252,31,130,31,34,31,241,31,241,30,187,31,206,31,206,30,206,29,96,31,253,31,253,30,250,31,199,31,233,31,169,31,252,31,71,31,71,30,71,29,71,28,166,31,5,31,119,31,162,31,108,31,162,31,110,31,157,31,157,30,180,31,212,31,212,30,40,31,251,31,13,31,160,31,130,31,165,31,157,31,157,30,247,31,247,30,237,31,188,31,30,31,115,31,128,31,232,31,216,31,56,31,56,30,69,31,69,30,69,29,156,31,152,31,163,31,110,31,110,30,110,29,178,31,102,31,232,31,231,31,220,31,232,31,148,31,131,31,16,31,4,31,205,31,21,31,227,31,51,31,51,30,15,31,182,31,137,31,108,31,108,30,157,31,225,31,221,31,246,31,246,30,189,31,233,31,90,31,90,30,90,29,157,31,157,30,178,31,243,31,243,30,114,31,114,30,60,31,223,31,246,31,182,31,182,30,113,31,112,31,68,31,68,30,23,31,1,31,232,31,102,31,79,31,141,31,55,31,171,31,208,31,230,31,177,31,235,31,11,31,168,31,119,31,177,31,198,31,209,31,74,31,74,30,74,29,179,31,111,31,111,30,137,31,32,31,22,31,99,31,201,31,201,30,236,31,211,31,3,31,6,31,221,31,121,31,134,31,134,30,176,31,19,31,115,31,246,31,246,30,246,29,222,31,222,30,160,31,160,30,192,31,218,31,52,31,2,31,64,31,27,31,27,30,27,29,27,28,114,31,91,31,129,31,236,31,49,31,67,31,85,31,85,30,196,31,4,31,4,30,41,31,41,30,41,29,228,31,228,30,206,31,228,31,177,31,181,31,35,31,100,31,245,31,245,30,73,31,17,31,17,30,20,31,239,31,251,31,96,31,29,31,29,30,155,31,68,31,63,31,141,31,9,31,7,31,77,31,77,30,75,31,104,31,104,30,205,31,143,31,132,31,132,30,48,31,48,30,54,31,100,31,210,31,37,31,37,30,75,31,49,31,137,31,254,31,132,31,169,31,239,31,247,31,247,30,69,31,26,31,22,31,159,31,236,31,53,31,24,31,220,31,54,31,120,31,139,31,29,31,66,31,66,30,112,31,112,30,213,31,213,30,213,29,39,31,35,31,136,31,136,30,136,29,198,31,198,30,193,31,22,31,208,31,208,30,57,31,188,31,7,31,180,31,81,31,139,31,102,31,102,30,194,31,224,31,53,31,38,31,231,31,194,31,194,30,220,31,220,30,221,31,221,30,152,31,67,31,172,31,6,31,52,31,118,31,79,31,236,31,57,31,244,31,194,31,51,31,135,31,69,31,3,31,3,30,3,29,79,31,214,31,214,30,126,31,118,31,97,31,97,30,30,31,30,30,207,31,80,31,80,30,132,31,199,31,79,31,134,31,5,31,206,31,19,31,245,31,87,31,23,31,226,31,39,31,162,31,81,31,81,30,142,31,109,31,180,31,204,31,101,31,42,31,159,31,26,31,131,31,120,31,120,30,138,31,138,30,140,31,140,30,140,29,98,31,73,31,199,31,245,31,140,31,232,31,26,31,131,31,131,30,131,29,3,31,176,31,176,30,176,29,199,31,92,31,179,31,154,31,252,31,140,31,177,31,177,30,255,31,255,30,161,31,161,30,58,31,58,30,221,31,174,31,203,31,52,31,52,30,217,31,69,31,127,31,233,31,90,31,17,31,248,31,54,31,238,31,122,31,122,30,219,31,219,30,38,31,235,31,229,31,229,30,173,31,252,31,62,31,62,30,210,31,210,30,36,31,125,31,138,31,138,30,70,31,70,30,70,29,129,31,47,31,212,31,12,31,12,30,119,31,96,31,71,31,175,31,190,31,190,30,68,31,32,31,32,30,22,31,221,31,26,31,248,31,235,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
