-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 882;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,252,0,20,0,52,0,0,0,184,0,194,0,0,0,103,0,64,0,0,0,92,0,3,0,17,0,206,0,197,0,78,0,0,0,79,0,0,0,103,0,47,0,38,0,86,0,135,0,65,0,0,0,115,0,101,0,0,0,0,0,80,0,84,0,226,0,7,0,0,0,122,0,122,0,0,0,0,0,237,0,140,0,172,0,100,0,117,0,0,0,123,0,153,0,197,0,0,0,154,0,72,0,129,0,189,0,149,0,97,0,116,0,199,0,0,0,168,0,178,0,126,0,228,0,231,0,154,0,30,0,240,0,0,0,210,0,34,0,47,0,104,0,164,0,195,0,36,0,139,0,172,0,195,0,124,0,40,0,230,0,185,0,220,0,239,0,69,0,118,0,0,0,2,0,219,0,112,0,57,0,206,0,135,0,252,0,149,0,221,0,20,0,0,0,149,0,5,0,169,0,0,0,189,0,177,0,34,0,72,0,255,0,188,0,217,0,123,0,216,0,237,0,173,0,37,0,207,0,0,0,148,0,204,0,148,0,136,0,23,0,48,0,231,0,248,0,75,0,0,0,153,0,74,0,113,0,0,0,197,0,44,0,209,0,131,0,34,0,0,0,0,0,53,0,79,0,0,0,9,0,153,0,161,0,0,0,144,0,0,0,128,0,47,0,230,0,248,0,0,0,120,0,0,0,16,0,12,0,205,0,0,0,128,0,65,0,180,0,43,0,181,0,63,0,77,0,203,0,0,0,17,0,0,0,228,0,36,0,64,0,0,0,100,0,149,0,121,0,110,0,0,0,104,0,50,0,90,0,102,0,0,0,89,0,249,0,49,0,183,0,46,0,87,0,123,0,99,0,77,0,6,0,235,0,157,0,208,0,0,0,12,0,51,0,43,0,230,0,0,0,120,0,34,0,227,0,149,0,78,0,29,0,214,0,0,0,121,0,196,0,134,0,229,0,105,0,2,0,13,0,99,0,52,0,0,0,120,0,187,0,74,0,65,0,0,0,29,0,189,0,3,0,0,0,249,0,53,0,102,0,30,0,253,0,160,0,169,0,69,0,179,0,77,0,0,0,254,0,81,0,188,0,12,0,101,0,203,0,188,0,0,0,151,0,0,0,169,0,116,0,0,0,0,0,134,0,246,0,202,0,219,0,186,0,0,0,209,0,28,0,31,0,227,0,184,0,121,0,208,0,3,0,41,0,192,0,218,0,143,0,150,0,243,0,0,0,44,0,9,0,159,0,209,0,118,0,218,0,223,0,155,0,154,0,210,0,0,0,0,0,226,0,0,0,117,0,162,0,128,0,212,0,192,0,13,0,244,0,155,0,72,0,223,0,175,0,103,0,226,0,170,0,130,0,61,0,132,0,213,0,174,0,226,0,81,0,173,0,142,0,38,0,101,0,165,0,59,0,226,0,172,0,180,0,53,0,78,0,168,0,0,0,162,0,45,0,213,0,233,0,169,0,212,0,186,0,180,0,7,0,249,0,175,0,201,0,62,0,0,0,65,0,23,0,0,0,146,0,122,0,15,0,0,0,165,0,0,0,2,0,255,0,0,0,190,0,235,0,183,0,55,0,188,0,92,0,3,0,0,0,60,0,148,0,0,0,225,0,31,0,110,0,61,0,100,0,27,0,129,0,192,0,133,0,137,0,153,0,198,0,61,0,146,0,0,0,20,0,22,0,55,0,221,0,20,0,164,0,171,0,119,0,0,0,151,0,180,0,76,0,120,0,131,0,0,0,0,0,202,0,33,0,0,0,158,0,84,0,171,0,213,0,61,0,74,0,213,0,231,0,0,0,208,0,109,0,0,0,47,0,0,0,120,0,105,0,0,0,0,0,241,0,113,0,71,0,181,0,108,0,0,0,247,0,194,0,129,0,0,0,226,0,191,0,91,0,186,0,86,0,0,0,4,0,180,0,0,0,0,0,209,0,0,0,236,0,139,0,138,0,0,0,25,0,126,0,154,0,87,0,211,0,135,0,70,0,181,0,147,0,209,0,135,0,216,0,36,0,0,0,0,0,109,0,123,0,143,0,0,0,0,0,190,0,196,0,89,0,194,0,47,0,34,0,153,0,0,0,78,0,104,0,170,0,96,0,117,0,0,0,0,0,0,0,12,0,0,0,223,0,93,0,62,0,180,0,0,0,90,0,53,0,93,0,0,0,65,0,0,0,105,0,193,0,0,0,181,0,38,0,0,0,221,0,151,0,108,0,67,0,135,0,0,0,205,0,81,0,0,0,128,0,239,0,0,0,115,0,195,0,0,0,131,0,103,0,0,0,0,0,0,0,50,0,0,0,25,0,42,0,32,0,133,0,69,0,101,0,144,0,119,0,227,0,122,0,142,0,0,0,0,0,164,0,23,0,251,0,244,0,255,0,218,0,101,0,237,0,60,0,81,0,59,0,99,0,108,0,219,0,161,0,46,0,62,0,240,0,169,0,159,0,60,0,195,0,232,0,77,0,3,0,236,0,139,0,0,0,201,0,0,0,193,0,70,0,58,0,103,0,0,0,71,0,128,0,201,0,119,0,12,0,19,0,250,0,203,0,242,0,146,0,32,0,137,0,0,0,141,0,223,0,101,0,0,0,172,0,168,0,130,0,0,0,122,0,89,0,60,0,119,0,75,0,35,0,99,0,67,0,188,0,0,0,128,0,85,0,149,0,71,0,188,0,104,0,0,0,202,0,0,0,231,0,16,0,209,0,81,0,61,0,122,0,0,0,157,0,20,0,8,0,8,0,228,0,137,0,236,0,51,0,0,0,199,0,0,0,106,0,115,0,0,0,197,0,0,0,79,0,0,0,145,0,117,0,70,0,194,0,0,0,199,0,91,0,125,0,0,0,57,0,98,0,81,0,28,0,0,0,0,0,0,0,0,0,45,0,17,0,173,0,125,0,233,0,0,0,144,0,69,0,190,0,0,0,121,0,46,0,0,0,43,0,213,0,115,0,169,0,92,0,92,0,15,0,183,0,0,0,81,0,93,0,0,0,68,0,200,0,140,0,157,0,0,0,58,0,39,0,195,0,25,0,75,0,51,0,0,0,211,0,58,0,104,0,79,0,57,0,109,0,0,0,0,0,5,0,0,0,254,0,82,0,13,0,167,0,0,0,201,0,59,0,0,0,84,0,137,0,2,0,95,0,0,0,44,0,163,0,241,0,101,0,0,0,45,0,0,0,83,0,0,0,162,0,240,0,0,0,68,0,12,0,239,0,248,0,22,0,152,0,114,0,0,0,212,0,243,0,0,0,157,0,185,0,6,0,219,0,0,0,40,0,219,0,236,0,66,0,118,0,104,0,70,0,85,0,239,0,164,0,249,0,0,0,169,0,34,0,170,0,254,0,49,0,168,0,47,0,60,0,0,0,61,0,0,0,0,0,0,0,70,0,0,0,221,0,0,0,130,0,243,0,215,0,205,0,89,0,172,0,77,0,0,0,229,0,0,0,169,0,237,0,81,0,9,0,91,0,97,0,5,0,255,0,242,0,0,0,103,0,0,0,0,0,145,0,175,0,241,0,90,0,246,0,65,0,111,0,0,0,118,0,236,0,174,0,49,0,0,0,218,0,0,0,0,0,181,0,85,0,219,0,3,0,214,0,61,0,226,0,1,0,0,0,0,0,204,0,34,0,0,0,236,0,248,0,0,0,16,0,142,0,171,0,124,0,2,0,102,0,225,0,238,0,254,0,206,0,32,0,0,0,156,0,196,0,140,0,42,0,70,0,185,0,62,0,79,0,137,0,235,0,0,0,0,0,0,0,26,0,15,0,139,0,0,0,0,0,0,0,182,0,201,0,216,0,133,0,114,0,0,0,154,0,148,0,97,0,98,0,144,0,0,0,252,0,103,0,0,0,36,0,28,0,149,0,177,0,255,0,106,0,139,0,0,0,148,0,78,0,149,0,38,0,122,0,234,0,154,0,179,0,59,0,49,0,165,0,0,0);
signal scenario_full  : scenario_type := (0,0,252,31,20,31,52,31,52,30,184,31,194,31,194,30,103,31,64,31,64,30,92,31,3,31,17,31,206,31,197,31,78,31,78,30,79,31,79,30,103,31,47,31,38,31,86,31,135,31,65,31,65,30,115,31,101,31,101,30,101,29,80,31,84,31,226,31,7,31,7,30,122,31,122,31,122,30,122,29,237,31,140,31,172,31,100,31,117,31,117,30,123,31,153,31,197,31,197,30,154,31,72,31,129,31,189,31,149,31,97,31,116,31,199,31,199,30,168,31,178,31,126,31,228,31,231,31,154,31,30,31,240,31,240,30,210,31,34,31,47,31,104,31,164,31,195,31,36,31,139,31,172,31,195,31,124,31,40,31,230,31,185,31,220,31,239,31,69,31,118,31,118,30,2,31,219,31,112,31,57,31,206,31,135,31,252,31,149,31,221,31,20,31,20,30,149,31,5,31,169,31,169,30,189,31,177,31,34,31,72,31,255,31,188,31,217,31,123,31,216,31,237,31,173,31,37,31,207,31,207,30,148,31,204,31,148,31,136,31,23,31,48,31,231,31,248,31,75,31,75,30,153,31,74,31,113,31,113,30,197,31,44,31,209,31,131,31,34,31,34,30,34,29,53,31,79,31,79,30,9,31,153,31,161,31,161,30,144,31,144,30,128,31,47,31,230,31,248,31,248,30,120,31,120,30,16,31,12,31,205,31,205,30,128,31,65,31,180,31,43,31,181,31,63,31,77,31,203,31,203,30,17,31,17,30,228,31,36,31,64,31,64,30,100,31,149,31,121,31,110,31,110,30,104,31,50,31,90,31,102,31,102,30,89,31,249,31,49,31,183,31,46,31,87,31,123,31,99,31,77,31,6,31,235,31,157,31,208,31,208,30,12,31,51,31,43,31,230,31,230,30,120,31,34,31,227,31,149,31,78,31,29,31,214,31,214,30,121,31,196,31,134,31,229,31,105,31,2,31,13,31,99,31,52,31,52,30,120,31,187,31,74,31,65,31,65,30,29,31,189,31,3,31,3,30,249,31,53,31,102,31,30,31,253,31,160,31,169,31,69,31,179,31,77,31,77,30,254,31,81,31,188,31,12,31,101,31,203,31,188,31,188,30,151,31,151,30,169,31,116,31,116,30,116,29,134,31,246,31,202,31,219,31,186,31,186,30,209,31,28,31,31,31,227,31,184,31,121,31,208,31,3,31,41,31,192,31,218,31,143,31,150,31,243,31,243,30,44,31,9,31,159,31,209,31,118,31,218,31,223,31,155,31,154,31,210,31,210,30,210,29,226,31,226,30,117,31,162,31,128,31,212,31,192,31,13,31,244,31,155,31,72,31,223,31,175,31,103,31,226,31,170,31,130,31,61,31,132,31,213,31,174,31,226,31,81,31,173,31,142,31,38,31,101,31,165,31,59,31,226,31,172,31,180,31,53,31,78,31,168,31,168,30,162,31,45,31,213,31,233,31,169,31,212,31,186,31,180,31,7,31,249,31,175,31,201,31,62,31,62,30,65,31,23,31,23,30,146,31,122,31,15,31,15,30,165,31,165,30,2,31,255,31,255,30,190,31,235,31,183,31,55,31,188,31,92,31,3,31,3,30,60,31,148,31,148,30,225,31,31,31,110,31,61,31,100,31,27,31,129,31,192,31,133,31,137,31,153,31,198,31,61,31,146,31,146,30,20,31,22,31,55,31,221,31,20,31,164,31,171,31,119,31,119,30,151,31,180,31,76,31,120,31,131,31,131,30,131,29,202,31,33,31,33,30,158,31,84,31,171,31,213,31,61,31,74,31,213,31,231,31,231,30,208,31,109,31,109,30,47,31,47,30,120,31,105,31,105,30,105,29,241,31,113,31,71,31,181,31,108,31,108,30,247,31,194,31,129,31,129,30,226,31,191,31,91,31,186,31,86,31,86,30,4,31,180,31,180,30,180,29,209,31,209,30,236,31,139,31,138,31,138,30,25,31,126,31,154,31,87,31,211,31,135,31,70,31,181,31,147,31,209,31,135,31,216,31,36,31,36,30,36,29,109,31,123,31,143,31,143,30,143,29,190,31,196,31,89,31,194,31,47,31,34,31,153,31,153,30,78,31,104,31,170,31,96,31,117,31,117,30,117,29,117,28,12,31,12,30,223,31,93,31,62,31,180,31,180,30,90,31,53,31,93,31,93,30,65,31,65,30,105,31,193,31,193,30,181,31,38,31,38,30,221,31,151,31,108,31,67,31,135,31,135,30,205,31,81,31,81,30,128,31,239,31,239,30,115,31,195,31,195,30,131,31,103,31,103,30,103,29,103,28,50,31,50,30,25,31,42,31,32,31,133,31,69,31,101,31,144,31,119,31,227,31,122,31,142,31,142,30,142,29,164,31,23,31,251,31,244,31,255,31,218,31,101,31,237,31,60,31,81,31,59,31,99,31,108,31,219,31,161,31,46,31,62,31,240,31,169,31,159,31,60,31,195,31,232,31,77,31,3,31,236,31,139,31,139,30,201,31,201,30,193,31,70,31,58,31,103,31,103,30,71,31,128,31,201,31,119,31,12,31,19,31,250,31,203,31,242,31,146,31,32,31,137,31,137,30,141,31,223,31,101,31,101,30,172,31,168,31,130,31,130,30,122,31,89,31,60,31,119,31,75,31,35,31,99,31,67,31,188,31,188,30,128,31,85,31,149,31,71,31,188,31,104,31,104,30,202,31,202,30,231,31,16,31,209,31,81,31,61,31,122,31,122,30,157,31,20,31,8,31,8,31,228,31,137,31,236,31,51,31,51,30,199,31,199,30,106,31,115,31,115,30,197,31,197,30,79,31,79,30,145,31,117,31,70,31,194,31,194,30,199,31,91,31,125,31,125,30,57,31,98,31,81,31,28,31,28,30,28,29,28,28,28,27,45,31,17,31,173,31,125,31,233,31,233,30,144,31,69,31,190,31,190,30,121,31,46,31,46,30,43,31,213,31,115,31,169,31,92,31,92,31,15,31,183,31,183,30,81,31,93,31,93,30,68,31,200,31,140,31,157,31,157,30,58,31,39,31,195,31,25,31,75,31,51,31,51,30,211,31,58,31,104,31,79,31,57,31,109,31,109,30,109,29,5,31,5,30,254,31,82,31,13,31,167,31,167,30,201,31,59,31,59,30,84,31,137,31,2,31,95,31,95,30,44,31,163,31,241,31,101,31,101,30,45,31,45,30,83,31,83,30,162,31,240,31,240,30,68,31,12,31,239,31,248,31,22,31,152,31,114,31,114,30,212,31,243,31,243,30,157,31,185,31,6,31,219,31,219,30,40,31,219,31,236,31,66,31,118,31,104,31,70,31,85,31,239,31,164,31,249,31,249,30,169,31,34,31,170,31,254,31,49,31,168,31,47,31,60,31,60,30,61,31,61,30,61,29,61,28,70,31,70,30,221,31,221,30,130,31,243,31,215,31,205,31,89,31,172,31,77,31,77,30,229,31,229,30,169,31,237,31,81,31,9,31,91,31,97,31,5,31,255,31,242,31,242,30,103,31,103,30,103,29,145,31,175,31,241,31,90,31,246,31,65,31,111,31,111,30,118,31,236,31,174,31,49,31,49,30,218,31,218,30,218,29,181,31,85,31,219,31,3,31,214,31,61,31,226,31,1,31,1,30,1,29,204,31,34,31,34,30,236,31,248,31,248,30,16,31,142,31,171,31,124,31,2,31,102,31,225,31,238,31,254,31,206,31,32,31,32,30,156,31,196,31,140,31,42,31,70,31,185,31,62,31,79,31,137,31,235,31,235,30,235,29,235,28,26,31,15,31,139,31,139,30,139,29,139,28,182,31,201,31,216,31,133,31,114,31,114,30,154,31,148,31,97,31,98,31,144,31,144,30,252,31,103,31,103,30,36,31,28,31,149,31,177,31,255,31,106,31,139,31,139,30,148,31,78,31,149,31,38,31,122,31,234,31,154,31,179,31,59,31,49,31,165,31,165,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
