-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_199 is
end project_tb_199;

architecture project_tb_arch_199 of project_tb_199 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 823;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (13,0,188,0,244,0,78,0,120,0,65,0,177,0,44,0,147,0,103,0,171,0,30,0,203,0,83,0,28,0,0,0,250,0,112,0,0,0,48,0,50,0,193,0,126,0,0,0,244,0,167,0,199,0,3,0,196,0,96,0,245,0,4,0,113,0,203,0,67,0,0,0,225,0,92,0,0,0,85,0,172,0,119,0,217,0,39,0,213,0,50,0,222,0,184,0,4,0,175,0,48,0,190,0,107,0,199,0,89,0,0,0,222,0,164,0,180,0,0,0,120,0,3,0,43,0,196,0,106,0,0,0,123,0,245,0,231,0,230,0,0,0,0,0,27,0,36,0,110,0,47,0,237,0,177,0,32,0,215,0,38,0,171,0,0,0,0,0,254,0,45,0,0,0,253,0,145,0,43,0,0,0,101,0,209,0,17,0,0,0,201,0,166,0,0,0,224,0,0,0,198,0,24,0,170,0,29,0,0,0,194,0,177,0,0,0,206,0,250,0,112,0,62,0,115,0,53,0,0,0,0,0,0,0,183,0,0,0,199,0,12,0,82,0,188,0,87,0,163,0,198,0,175,0,0,0,185,0,0,0,10,0,85,0,0,0,0,0,180,0,134,0,1,0,0,0,195,0,25,0,180,0,121,0,235,0,0,0,29,0,45,0,246,0,36,0,36,0,0,0,129,0,218,0,20,0,0,0,95,0,61,0,170,0,0,0,0,0,238,0,3,0,160,0,178,0,194,0,103,0,48,0,0,0,0,0,92,0,77,0,192,0,159,0,13,0,197,0,155,0,245,0,182,0,116,0,225,0,96,0,0,0,17,0,206,0,147,0,66,0,187,0,26,0,6,0,106,0,12,0,0,0,133,0,92,0,112,0,74,0,192,0,115,0,183,0,176,0,111,0,145,0,18,0,0,0,106,0,13,0,54,0,10,0,249,0,7,0,0,0,132,0,162,0,150,0,231,0,54,0,186,0,0,0,132,0,40,0,134,0,13,0,140,0,208,0,252,0,192,0,208,0,26,0,37,0,0,0,160,0,202,0,7,0,233,0,196,0,144,0,62,0,49,0,218,0,22,0,0,0,162,0,109,0,244,0,35,0,232,0,0,0,206,0,200,0,88,0,117,0,37,0,0,0,243,0,246,0,38,0,140,0,103,0,241,0,0,0,1,0,0,0,199,0,230,0,47,0,0,0,181,0,48,0,65,0,75,0,157,0,45,0,26,0,224,0,254,0,51,0,94,0,235,0,110,0,0,0,243,0,0,0,201,0,76,0,23,0,239,0,147,0,194,0,238,0,115,0,135,0,0,0,77,0,68,0,4,0,0,0,160,0,249,0,182,0,30,0,69,0,0,0,15,0,0,0,95,0,106,0,0,0,195,0,152,0,89,0,0,0,252,0,164,0,20,0,5,0,208,0,54,0,0,0,0,0,0,0,75,0,0,0,66,0,103,0,0,0,0,0,19,0,201,0,253,0,0,0,178,0,229,0,124,0,165,0,176,0,237,0,50,0,156,0,106,0,153,0,229,0,248,0,0,0,180,0,155,0,161,0,170,0,144,0,88,0,73,0,0,0,198,0,102,0,106,0,11,0,109,0,67,0,186,0,197,0,144,0,129,0,73,0,163,0,194,0,112,0,29,0,0,0,57,0,220,0,126,0,159,0,0,0,110,0,65,0,179,0,196,0,116,0,0,0,149,0,6,0,221,0,71,0,89,0,3,0,165,0,0,0,109,0,0,0,230,0,9,0,241,0,242,0,52,0,0,0,170,0,171,0,209,0,225,0,56,0,0,0,91,0,0,0,0,0,172,0,251,0,30,0,193,0,148,0,189,0,191,0,239,0,207,0,0,0,214,0,154,0,202,0,136,0,150,0,44,0,106,0,200,0,0,0,74,0,82,0,173,0,90,0,0,0,238,0,187,0,228,0,241,0,25,0,56,0,175,0,218,0,227,0,192,0,247,0,160,0,0,0,85,0,0,0,139,0,126,0,157,0,180,0,0,0,190,0,128,0,222,0,234,0,213,0,170,0,221,0,0,0,165,0,249,0,182,0,149,0,69,0,0,0,161,0,31,0,114,0,16,0,97,0,36,0,59,0,193,0,0,0,169,0,0,0,43,0,0,0,0,0,0,0,218,0,43,0,174,0,110,0,0,0,173,0,250,0,218,0,40,0,108,0,0,0,214,0,76,0,136,0,50,0,75,0,251,0,86,0,66,0,121,0,176,0,85,0,216,0,6,0,38,0,61,0,61,0,1,0,148,0,0,0,125,0,77,0,19,0,0,0,111,0,0,0,0,0,246,0,79,0,183,0,15,0,147,0,0,0,166,0,138,0,240,0,247,0,102,0,0,0,7,0,75,0,94,0,0,0,72,0,20,0,75,0,146,0,0,0,0,0,0,0,142,0,254,0,68,0,117,0,0,0,192,0,1,0,0,0,174,0,61,0,180,0,154,0,102,0,60,0,0,0,74,0,10,0,8,0,34,0,229,0,186,0,0,0,148,0,96,0,148,0,40,0,0,0,251,0,171,0,53,0,187,0,123,0,0,0,248,0,75,0,147,0,0,0,157,0,79,0,188,0,0,0,74,0,0,0,220,0,84,0,1,0,81,0,221,0,99,0,49,0,254,0,0,0,107,0,104,0,237,0,209,0,232,0,62,0,0,0,249,0,0,0,254,0,12,0,227,0,0,0,194,0,141,0,221,0,145,0,198,0,126,0,73,0,0,0,94,0,133,0,40,0,0,0,0,0,217,0,182,0,0,0,25,0,233,0,41,0,182,0,154,0,195,0,199,0,93,0,104,0,0,0,196,0,0,0,222,0,211,0,58,0,203,0,105,0,150,0,113,0,94,0,179,0,227,0,73,0,221,0,51,0,22,0,20,0,0,0,207,0,130,0,114,0,123,0,3,0,107,0,30,0,234,0,231,0,111,0,188,0,60,0,147,0,41,0,122,0,166,0,186,0,129,0,77,0,12,0,0,0,16,0,0,0,225,0,233,0,162,0,61,0,243,0,27,0,30,0,2,0,198,0,212,0,177,0,235,0,122,0,240,0,86,0,169,0,0,0,0,0,98,0,52,0,0,0,0,0,110,0,0,0,54,0,63,0,69,0,0,0,0,0,201,0,0,0,127,0,92,0,163,0,21,0,26,0,101,0,0,0,39,0,100,0,89,0,98,0,81,0,81,0,133,0,180,0,3,0,108,0,241,0,0,0,24,0,242,0,211,0,224,0,42,0,133,0,217,0,22,0,64,0,157,0,252,0,52,0,72,0,74,0,220,0,192,0,32,0,217,0,140,0,163,0,0,0,100,0,255,0,155,0,200,0,13,0,202,0,5,0,154,0,174,0,133,0,163,0,241,0,127,0,213,0,234,0,213,0,95,0,117,0,142,0,0,0,9,0,6,0,102,0,155,0,165,0,66,0,182,0,225,0,38,0,86,0,170,0,57,0,0,0,47,0,0,0,82,0,55,0,0,0,0,0,192,0,7,0,80,0,176,0,37,0,68,0,0,0,97,0,209,0,254,0,20,0,0,0,83,0,79,0,94,0,55,0,243,0,48,0,10,0,167,0,144,0,152,0,28,0,40,0,42,0,203,0,135,0,0,0,0,0,51,0,103,0,68,0,151,0,0,0,238,0,46,0,174,0,196,0,82,0,110,0,52,0,88,0,74,0,115,0,96,0,0,0);
signal scenario_full  : scenario_type := (13,31,188,31,244,31,78,31,120,31,65,31,177,31,44,31,147,31,103,31,171,31,30,31,203,31,83,31,28,31,28,30,250,31,112,31,112,30,48,31,50,31,193,31,126,31,126,30,244,31,167,31,199,31,3,31,196,31,96,31,245,31,4,31,113,31,203,31,67,31,67,30,225,31,92,31,92,30,85,31,172,31,119,31,217,31,39,31,213,31,50,31,222,31,184,31,4,31,175,31,48,31,190,31,107,31,199,31,89,31,89,30,222,31,164,31,180,31,180,30,120,31,3,31,43,31,196,31,106,31,106,30,123,31,245,31,231,31,230,31,230,30,230,29,27,31,36,31,110,31,47,31,237,31,177,31,32,31,215,31,38,31,171,31,171,30,171,29,254,31,45,31,45,30,253,31,145,31,43,31,43,30,101,31,209,31,17,31,17,30,201,31,166,31,166,30,224,31,224,30,198,31,24,31,170,31,29,31,29,30,194,31,177,31,177,30,206,31,250,31,112,31,62,31,115,31,53,31,53,30,53,29,53,28,183,31,183,30,199,31,12,31,82,31,188,31,87,31,163,31,198,31,175,31,175,30,185,31,185,30,10,31,85,31,85,30,85,29,180,31,134,31,1,31,1,30,195,31,25,31,180,31,121,31,235,31,235,30,29,31,45,31,246,31,36,31,36,31,36,30,129,31,218,31,20,31,20,30,95,31,61,31,170,31,170,30,170,29,238,31,3,31,160,31,178,31,194,31,103,31,48,31,48,30,48,29,92,31,77,31,192,31,159,31,13,31,197,31,155,31,245,31,182,31,116,31,225,31,96,31,96,30,17,31,206,31,147,31,66,31,187,31,26,31,6,31,106,31,12,31,12,30,133,31,92,31,112,31,74,31,192,31,115,31,183,31,176,31,111,31,145,31,18,31,18,30,106,31,13,31,54,31,10,31,249,31,7,31,7,30,132,31,162,31,150,31,231,31,54,31,186,31,186,30,132,31,40,31,134,31,13,31,140,31,208,31,252,31,192,31,208,31,26,31,37,31,37,30,160,31,202,31,7,31,233,31,196,31,144,31,62,31,49,31,218,31,22,31,22,30,162,31,109,31,244,31,35,31,232,31,232,30,206,31,200,31,88,31,117,31,37,31,37,30,243,31,246,31,38,31,140,31,103,31,241,31,241,30,1,31,1,30,199,31,230,31,47,31,47,30,181,31,48,31,65,31,75,31,157,31,45,31,26,31,224,31,254,31,51,31,94,31,235,31,110,31,110,30,243,31,243,30,201,31,76,31,23,31,239,31,147,31,194,31,238,31,115,31,135,31,135,30,77,31,68,31,4,31,4,30,160,31,249,31,182,31,30,31,69,31,69,30,15,31,15,30,95,31,106,31,106,30,195,31,152,31,89,31,89,30,252,31,164,31,20,31,5,31,208,31,54,31,54,30,54,29,54,28,75,31,75,30,66,31,103,31,103,30,103,29,19,31,201,31,253,31,253,30,178,31,229,31,124,31,165,31,176,31,237,31,50,31,156,31,106,31,153,31,229,31,248,31,248,30,180,31,155,31,161,31,170,31,144,31,88,31,73,31,73,30,198,31,102,31,106,31,11,31,109,31,67,31,186,31,197,31,144,31,129,31,73,31,163,31,194,31,112,31,29,31,29,30,57,31,220,31,126,31,159,31,159,30,110,31,65,31,179,31,196,31,116,31,116,30,149,31,6,31,221,31,71,31,89,31,3,31,165,31,165,30,109,31,109,30,230,31,9,31,241,31,242,31,52,31,52,30,170,31,171,31,209,31,225,31,56,31,56,30,91,31,91,30,91,29,172,31,251,31,30,31,193,31,148,31,189,31,191,31,239,31,207,31,207,30,214,31,154,31,202,31,136,31,150,31,44,31,106,31,200,31,200,30,74,31,82,31,173,31,90,31,90,30,238,31,187,31,228,31,241,31,25,31,56,31,175,31,218,31,227,31,192,31,247,31,160,31,160,30,85,31,85,30,139,31,126,31,157,31,180,31,180,30,190,31,128,31,222,31,234,31,213,31,170,31,221,31,221,30,165,31,249,31,182,31,149,31,69,31,69,30,161,31,31,31,114,31,16,31,97,31,36,31,59,31,193,31,193,30,169,31,169,30,43,31,43,30,43,29,43,28,218,31,43,31,174,31,110,31,110,30,173,31,250,31,218,31,40,31,108,31,108,30,214,31,76,31,136,31,50,31,75,31,251,31,86,31,66,31,121,31,176,31,85,31,216,31,6,31,38,31,61,31,61,31,1,31,148,31,148,30,125,31,77,31,19,31,19,30,111,31,111,30,111,29,246,31,79,31,183,31,15,31,147,31,147,30,166,31,138,31,240,31,247,31,102,31,102,30,7,31,75,31,94,31,94,30,72,31,20,31,75,31,146,31,146,30,146,29,146,28,142,31,254,31,68,31,117,31,117,30,192,31,1,31,1,30,174,31,61,31,180,31,154,31,102,31,60,31,60,30,74,31,10,31,8,31,34,31,229,31,186,31,186,30,148,31,96,31,148,31,40,31,40,30,251,31,171,31,53,31,187,31,123,31,123,30,248,31,75,31,147,31,147,30,157,31,79,31,188,31,188,30,74,31,74,30,220,31,84,31,1,31,81,31,221,31,99,31,49,31,254,31,254,30,107,31,104,31,237,31,209,31,232,31,62,31,62,30,249,31,249,30,254,31,12,31,227,31,227,30,194,31,141,31,221,31,145,31,198,31,126,31,73,31,73,30,94,31,133,31,40,31,40,30,40,29,217,31,182,31,182,30,25,31,233,31,41,31,182,31,154,31,195,31,199,31,93,31,104,31,104,30,196,31,196,30,222,31,211,31,58,31,203,31,105,31,150,31,113,31,94,31,179,31,227,31,73,31,221,31,51,31,22,31,20,31,20,30,207,31,130,31,114,31,123,31,3,31,107,31,30,31,234,31,231,31,111,31,188,31,60,31,147,31,41,31,122,31,166,31,186,31,129,31,77,31,12,31,12,30,16,31,16,30,225,31,233,31,162,31,61,31,243,31,27,31,30,31,2,31,198,31,212,31,177,31,235,31,122,31,240,31,86,31,169,31,169,30,169,29,98,31,52,31,52,30,52,29,110,31,110,30,54,31,63,31,69,31,69,30,69,29,201,31,201,30,127,31,92,31,163,31,21,31,26,31,101,31,101,30,39,31,100,31,89,31,98,31,81,31,81,31,133,31,180,31,3,31,108,31,241,31,241,30,24,31,242,31,211,31,224,31,42,31,133,31,217,31,22,31,64,31,157,31,252,31,52,31,72,31,74,31,220,31,192,31,32,31,217,31,140,31,163,31,163,30,100,31,255,31,155,31,200,31,13,31,202,31,5,31,154,31,174,31,133,31,163,31,241,31,127,31,213,31,234,31,213,31,95,31,117,31,142,31,142,30,9,31,6,31,102,31,155,31,165,31,66,31,182,31,225,31,38,31,86,31,170,31,57,31,57,30,47,31,47,30,82,31,55,31,55,30,55,29,192,31,7,31,80,31,176,31,37,31,68,31,68,30,97,31,209,31,254,31,20,31,20,30,83,31,79,31,94,31,55,31,243,31,48,31,10,31,167,31,144,31,152,31,28,31,40,31,42,31,203,31,135,31,135,30,135,29,51,31,103,31,68,31,151,31,151,30,238,31,46,31,174,31,196,31,82,31,110,31,52,31,88,31,74,31,115,31,96,31,96,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
