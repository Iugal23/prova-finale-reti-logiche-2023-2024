-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_247 is
end project_tb_247;

architecture project_tb_arch_247 of project_tb_247 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 950;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (71,0,7,0,191,0,20,0,121,0,180,0,227,0,48,0,154,0,162,0,39,0,37,0,3,0,218,0,117,0,174,0,190,0,150,0,220,0,133,0,0,0,137,0,251,0,220,0,0,0,0,0,135,0,34,0,177,0,105,0,187,0,25,0,142,0,0,0,203,0,207,0,42,0,14,0,7,0,68,0,151,0,1,0,40,0,0,0,202,0,0,0,0,0,165,0,92,0,41,0,0,0,0,0,16,0,191,0,201,0,178,0,53,0,0,0,67,0,55,0,3,0,191,0,242,0,127,0,228,0,43,0,81,0,0,0,48,0,101,0,212,0,228,0,115,0,116,0,0,0,0,0,146,0,112,0,135,0,51,0,57,0,0,0,248,0,0,0,190,0,165,0,15,0,122,0,201,0,0,0,0,0,29,0,152,0,55,0,229,0,7,0,151,0,20,0,81,0,60,0,0,0,49,0,140,0,11,0,184,0,12,0,107,0,182,0,104,0,252,0,183,0,0,0,11,0,57,0,93,0,69,0,0,0,209,0,61,0,0,0,222,0,164,0,230,0,210,0,46,0,180,0,0,0,111,0,91,0,195,0,229,0,143,0,242,0,46,0,133,0,0,0,130,0,132,0,81,0,80,0,207,0,19,0,0,0,244,0,61,0,57,0,0,0,246,0,0,0,182,0,18,0,0,0,186,0,0,0,150,0,239,0,177,0,0,0,0,0,138,0,61,0,0,0,74,0,15,0,247,0,162,0,194,0,66,0,42,0,81,0,21,0,0,0,237,0,3,0,181,0,109,0,174,0,152,0,8,0,174,0,119,0,0,0,248,0,101,0,200,0,91,0,0,0,19,0,123,0,0,0,252,0,233,0,83,0,9,0,0,0,3,0,58,0,0,0,0,0,0,0,58,0,181,0,147,0,0,0,161,0,94,0,145,0,76,0,176,0,197,0,12,0,68,0,122,0,20,0,209,0,37,0,53,0,240,0,104,0,244,0,224,0,35,0,172,0,122,0,0,0,104,0,0,0,242,0,83,0,46,0,62,0,146,0,193,0,0,0,0,0,149,0,178,0,87,0,250,0,178,0,252,0,172,0,241,0,241,0,99,0,190,0,237,0,177,0,0,0,11,0,26,0,67,0,0,0,0,0,0,0,150,0,124,0,247,0,231,0,150,0,107,0,245,0,229,0,246,0,145,0,232,0,233,0,52,0,194,0,0,0,224,0,155,0,169,0,234,0,102,0,0,0,0,0,29,0,30,0,211,0,124,0,19,0,6,0,0,0,0,0,0,0,8,0,128,0,5,0,0,0,99,0,96,0,93,0,62,0,62,0,130,0,59,0,109,0,254,0,81,0,0,0,163,0,126,0,188,0,20,0,152,0,239,0,0,0,158,0,0,0,165,0,135,0,145,0,154,0,168,0,147,0,234,0,49,0,135,0,0,0,211,0,0,0,222,0,175,0,208,0,223,0,108,0,206,0,75,0,135,0,120,0,98,0,242,0,149,0,240,0,0,0,13,0,24,0,220,0,108,0,0,0,168,0,0,0,170,0,214,0,0,0,0,0,234,0,225,0,129,0,38,0,129,0,10,0,174,0,189,0,0,0,0,0,32,0,165,0,0,0,74,0,146,0,175,0,10,0,0,0,47,0,0,0,0,0,59,0,1,0,244,0,77,0,0,0,0,0,208,0,51,0,189,0,161,0,74,0,0,0,158,0,103,0,243,0,0,0,139,0,216,0,249,0,162,0,187,0,240,0,39,0,197,0,69,0,0,0,248,0,0,0,38,0,141,0,0,0,187,0,208,0,134,0,76,0,171,0,219,0,242,0,46,0,206,0,22,0,11,0,17,0,67,0,44,0,202,0,0,0,212,0,104,0,214,0,215,0,110,0,246,0,36,0,16,0,229,0,37,0,198,0,70,0,48,0,176,0,177,0,62,0,88,0,103,0,17,0,87,0,223,0,204,0,78,0,201,0,200,0,129,0,19,0,30,0,49,0,0,0,192,0,17,0,64,0,51,0,119,0,224,0,14,0,137,0,92,0,0,0,6,0,223,0,0,0,46,0,195,0,89,0,168,0,203,0,31,0,187,0,195,0,147,0,66,0,56,0,43,0,177,0,253,0,0,0,0,0,176,0,196,0,206,0,0,0,95,0,103,0,0,0,146,0,14,0,203,0,95,0,16,0,0,0,1,0,140,0,245,0,73,0,228,0,0,0,201,0,198,0,123,0,166,0,71,0,161,0,0,0,158,0,110,0,0,0,80,0,0,0,220,0,142,0,244,0,89,0,150,0,214,0,130,0,0,0,95,0,12,0,128,0,194,0,109,0,15,0,74,0,5,0,133,0,0,0,26,0,0,0,0,0,0,0,13,0,135,0,0,0,180,0,116,0,32,0,183,0,88,0,211,0,20,0,69,0,144,0,122,0,15,0,113,0,254,0,69,0,215,0,0,0,0,0,165,0,107,0,0,0,143,0,90,0,0,0,0,0,83,0,107,0,0,0,136,0,20,0,0,0,60,0,165,0,194,0,0,0,102,0,244,0,17,0,0,0,245,0,175,0,204,0,100,0,77,0,0,0,0,0,165,0,59,0,163,0,141,0,216,0,174,0,251,0,248,0,141,0,141,0,78,0,83,0,243,0,0,0,0,0,28,0,66,0,18,0,146,0,83,0,203,0,0,0,248,0,137,0,0,0,0,0,0,0,140,0,0,0,240,0,0,0,0,0,105,0,0,0,37,0,214,0,38,0,23,0,13,0,0,0,169,0,12,0,124,0,79,0,197,0,50,0,172,0,206,0,248,0,140,0,201,0,250,0,172,0,164,0,164,0,237,0,101,0,151,0,110,0,26,0,224,0,179,0,0,0,155,0,189,0,194,0,255,0,15,0,218,0,200,0,230,0,30,0,146,0,154,0,154,0,205,0,9,0,220,0,153,0,64,0,154,0,115,0,139,0,212,0,63,0,205,0,173,0,3,0,0,0,223,0,207,0,46,0,63,0,127,0,132,0,0,0,54,0,232,0,0,0,12,0,30,0,183,0,196,0,207,0,212,0,88,0,59,0,77,0,65,0,74,0,215,0,116,0,161,0,247,0,158,0,169,0,0,0,8,0,73,0,97,0,0,0,157,0,126,0,217,0,0,0,0,0,0,0,123,0,0,0,15,0,255,0,52,0,121,0,252,0,0,0,120,0,110,0,151,0,141,0,179,0,50,0,238,0,184,0,81,0,213,0,18,0,0,0,238,0,10,0,167,0,139,0,0,0,0,0,92,0,226,0,13,0,68,0,95,0,200,0,0,0,0,0,62,0,0,0,204,0,178,0,22,0,143,0,0,0,216,0,107,0,0,0,89,0,0,0,0,0,216,0,27,0,44,0,56,0,59,0,91,0,28,0,247,0,9,0,0,0,14,0,131,0,116,0,72,0,252,0,253,0,187,0,138,0,179,0,62,0,167,0,217,0,101,0,0,0,54,0,191,0,0,0,0,0,230,0,133,0,0,0,54,0,130,0,180,0,41,0,41,0,198,0,247,0,142,0,153,0,181,0,149,0,80,0,53,0,236,0,0,0,245,0,0,0,0,0,0,0,39,0,240,0,0,0,28,0,174,0,231,0,115,0,65,0,0,0,208,0,64,0,78,0,0,0,20,0,69,0,210,0,224,0,0,0,223,0,78,0,33,0,0,0,63,0,169,0,221,0,184,0,255,0,127,0,13,0,90,0,0,0,41,0,4,0,203,0,0,0,244,0,250,0,142,0,207,0,39,0,113,0,7,0,26,0,234,0,139,0,78,0,178,0,159,0,100,0,164,0,0,0,0,0,205,0,101,0,209,0,0,0,140,0,12,0,8,0,47,0,0,0,66,0,245,0,0,0,16,0,208,0,52,0,170,0,80,0,61,0,250,0,34,0,0,0,43,0,37,0,0,0,27,0,192,0,68,0,240,0,104,0,210,0,173,0,0,0,0,0,239,0,131,0,88,0,130,0,55,0,22,0,0,0,57,0,178,0,80,0,160,0,121,0,96,0,227,0,173,0,175,0,2,0,233,0,72,0,217,0,0,0,11,0,0,0,217,0,148,0,0,0,0,0,7,0,125,0,56,0,253,0,0,0,57,0,205,0,0,0,39,0,255,0,222,0,54,0,24,0,32,0,0,0,0,0,178,0,51,0,223,0,188,0,0,0,218,0,133,0,232,0,254,0,135,0,29,0,145,0,141,0,204,0,137,0,194,0,0,0,65,0,120,0,146,0,0,0,210,0,0,0);
signal scenario_full  : scenario_type := (71,31,7,31,191,31,20,31,121,31,180,31,227,31,48,31,154,31,162,31,39,31,37,31,3,31,218,31,117,31,174,31,190,31,150,31,220,31,133,31,133,30,137,31,251,31,220,31,220,30,220,29,135,31,34,31,177,31,105,31,187,31,25,31,142,31,142,30,203,31,207,31,42,31,14,31,7,31,68,31,151,31,1,31,40,31,40,30,202,31,202,30,202,29,165,31,92,31,41,31,41,30,41,29,16,31,191,31,201,31,178,31,53,31,53,30,67,31,55,31,3,31,191,31,242,31,127,31,228,31,43,31,81,31,81,30,48,31,101,31,212,31,228,31,115,31,116,31,116,30,116,29,146,31,112,31,135,31,51,31,57,31,57,30,248,31,248,30,190,31,165,31,15,31,122,31,201,31,201,30,201,29,29,31,152,31,55,31,229,31,7,31,151,31,20,31,81,31,60,31,60,30,49,31,140,31,11,31,184,31,12,31,107,31,182,31,104,31,252,31,183,31,183,30,11,31,57,31,93,31,69,31,69,30,209,31,61,31,61,30,222,31,164,31,230,31,210,31,46,31,180,31,180,30,111,31,91,31,195,31,229,31,143,31,242,31,46,31,133,31,133,30,130,31,132,31,81,31,80,31,207,31,19,31,19,30,244,31,61,31,57,31,57,30,246,31,246,30,182,31,18,31,18,30,186,31,186,30,150,31,239,31,177,31,177,30,177,29,138,31,61,31,61,30,74,31,15,31,247,31,162,31,194,31,66,31,42,31,81,31,21,31,21,30,237,31,3,31,181,31,109,31,174,31,152,31,8,31,174,31,119,31,119,30,248,31,101,31,200,31,91,31,91,30,19,31,123,31,123,30,252,31,233,31,83,31,9,31,9,30,3,31,58,31,58,30,58,29,58,28,58,31,181,31,147,31,147,30,161,31,94,31,145,31,76,31,176,31,197,31,12,31,68,31,122,31,20,31,209,31,37,31,53,31,240,31,104,31,244,31,224,31,35,31,172,31,122,31,122,30,104,31,104,30,242,31,83,31,46,31,62,31,146,31,193,31,193,30,193,29,149,31,178,31,87,31,250,31,178,31,252,31,172,31,241,31,241,31,99,31,190,31,237,31,177,31,177,30,11,31,26,31,67,31,67,30,67,29,67,28,150,31,124,31,247,31,231,31,150,31,107,31,245,31,229,31,246,31,145,31,232,31,233,31,52,31,194,31,194,30,224,31,155,31,169,31,234,31,102,31,102,30,102,29,29,31,30,31,211,31,124,31,19,31,6,31,6,30,6,29,6,28,8,31,128,31,5,31,5,30,99,31,96,31,93,31,62,31,62,31,130,31,59,31,109,31,254,31,81,31,81,30,163,31,126,31,188,31,20,31,152,31,239,31,239,30,158,31,158,30,165,31,135,31,145,31,154,31,168,31,147,31,234,31,49,31,135,31,135,30,211,31,211,30,222,31,175,31,208,31,223,31,108,31,206,31,75,31,135,31,120,31,98,31,242,31,149,31,240,31,240,30,13,31,24,31,220,31,108,31,108,30,168,31,168,30,170,31,214,31,214,30,214,29,234,31,225,31,129,31,38,31,129,31,10,31,174,31,189,31,189,30,189,29,32,31,165,31,165,30,74,31,146,31,175,31,10,31,10,30,47,31,47,30,47,29,59,31,1,31,244,31,77,31,77,30,77,29,208,31,51,31,189,31,161,31,74,31,74,30,158,31,103,31,243,31,243,30,139,31,216,31,249,31,162,31,187,31,240,31,39,31,197,31,69,31,69,30,248,31,248,30,38,31,141,31,141,30,187,31,208,31,134,31,76,31,171,31,219,31,242,31,46,31,206,31,22,31,11,31,17,31,67,31,44,31,202,31,202,30,212,31,104,31,214,31,215,31,110,31,246,31,36,31,16,31,229,31,37,31,198,31,70,31,48,31,176,31,177,31,62,31,88,31,103,31,17,31,87,31,223,31,204,31,78,31,201,31,200,31,129,31,19,31,30,31,49,31,49,30,192,31,17,31,64,31,51,31,119,31,224,31,14,31,137,31,92,31,92,30,6,31,223,31,223,30,46,31,195,31,89,31,168,31,203,31,31,31,187,31,195,31,147,31,66,31,56,31,43,31,177,31,253,31,253,30,253,29,176,31,196,31,206,31,206,30,95,31,103,31,103,30,146,31,14,31,203,31,95,31,16,31,16,30,1,31,140,31,245,31,73,31,228,31,228,30,201,31,198,31,123,31,166,31,71,31,161,31,161,30,158,31,110,31,110,30,80,31,80,30,220,31,142,31,244,31,89,31,150,31,214,31,130,31,130,30,95,31,12,31,128,31,194,31,109,31,15,31,74,31,5,31,133,31,133,30,26,31,26,30,26,29,26,28,13,31,135,31,135,30,180,31,116,31,32,31,183,31,88,31,211,31,20,31,69,31,144,31,122,31,15,31,113,31,254,31,69,31,215,31,215,30,215,29,165,31,107,31,107,30,143,31,90,31,90,30,90,29,83,31,107,31,107,30,136,31,20,31,20,30,60,31,165,31,194,31,194,30,102,31,244,31,17,31,17,30,245,31,175,31,204,31,100,31,77,31,77,30,77,29,165,31,59,31,163,31,141,31,216,31,174,31,251,31,248,31,141,31,141,31,78,31,83,31,243,31,243,30,243,29,28,31,66,31,18,31,146,31,83,31,203,31,203,30,248,31,137,31,137,30,137,29,137,28,140,31,140,30,240,31,240,30,240,29,105,31,105,30,37,31,214,31,38,31,23,31,13,31,13,30,169,31,12,31,124,31,79,31,197,31,50,31,172,31,206,31,248,31,140,31,201,31,250,31,172,31,164,31,164,31,237,31,101,31,151,31,110,31,26,31,224,31,179,31,179,30,155,31,189,31,194,31,255,31,15,31,218,31,200,31,230,31,30,31,146,31,154,31,154,31,205,31,9,31,220,31,153,31,64,31,154,31,115,31,139,31,212,31,63,31,205,31,173,31,3,31,3,30,223,31,207,31,46,31,63,31,127,31,132,31,132,30,54,31,232,31,232,30,12,31,30,31,183,31,196,31,207,31,212,31,88,31,59,31,77,31,65,31,74,31,215,31,116,31,161,31,247,31,158,31,169,31,169,30,8,31,73,31,97,31,97,30,157,31,126,31,217,31,217,30,217,29,217,28,123,31,123,30,15,31,255,31,52,31,121,31,252,31,252,30,120,31,110,31,151,31,141,31,179,31,50,31,238,31,184,31,81,31,213,31,18,31,18,30,238,31,10,31,167,31,139,31,139,30,139,29,92,31,226,31,13,31,68,31,95,31,200,31,200,30,200,29,62,31,62,30,204,31,178,31,22,31,143,31,143,30,216,31,107,31,107,30,89,31,89,30,89,29,216,31,27,31,44,31,56,31,59,31,91,31,28,31,247,31,9,31,9,30,14,31,131,31,116,31,72,31,252,31,253,31,187,31,138,31,179,31,62,31,167,31,217,31,101,31,101,30,54,31,191,31,191,30,191,29,230,31,133,31,133,30,54,31,130,31,180,31,41,31,41,31,198,31,247,31,142,31,153,31,181,31,149,31,80,31,53,31,236,31,236,30,245,31,245,30,245,29,245,28,39,31,240,31,240,30,28,31,174,31,231,31,115,31,65,31,65,30,208,31,64,31,78,31,78,30,20,31,69,31,210,31,224,31,224,30,223,31,78,31,33,31,33,30,63,31,169,31,221,31,184,31,255,31,127,31,13,31,90,31,90,30,41,31,4,31,203,31,203,30,244,31,250,31,142,31,207,31,39,31,113,31,7,31,26,31,234,31,139,31,78,31,178,31,159,31,100,31,164,31,164,30,164,29,205,31,101,31,209,31,209,30,140,31,12,31,8,31,47,31,47,30,66,31,245,31,245,30,16,31,208,31,52,31,170,31,80,31,61,31,250,31,34,31,34,30,43,31,37,31,37,30,27,31,192,31,68,31,240,31,104,31,210,31,173,31,173,30,173,29,239,31,131,31,88,31,130,31,55,31,22,31,22,30,57,31,178,31,80,31,160,31,121,31,96,31,227,31,173,31,175,31,2,31,233,31,72,31,217,31,217,30,11,31,11,30,217,31,148,31,148,30,148,29,7,31,125,31,56,31,253,31,253,30,57,31,205,31,205,30,39,31,255,31,222,31,54,31,24,31,32,31,32,30,32,29,178,31,51,31,223,31,188,31,188,30,218,31,133,31,232,31,254,31,135,31,29,31,145,31,141,31,204,31,137,31,194,31,194,30,65,31,120,31,146,31,146,30,210,31,210,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
