-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 508;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (223,0,48,0,0,0,89,0,73,0,89,0,80,0,188,0,47,0,121,0,114,0,0,0,245,0,207,0,186,0,22,0,4,0,0,0,103,0,202,0,109,0,60,0,32,0,78,0,129,0,14,0,76,0,184,0,230,0,243,0,0,0,76,0,62,0,135,0,103,0,0,0,203,0,178,0,136,0,169,0,0,0,94,0,17,0,0,0,9,0,56,0,0,0,199,0,196,0,0,0,0,0,32,0,90,0,107,0,112,0,26,0,113,0,0,0,230,0,0,0,179,0,12,0,249,0,25,0,146,0,69,0,39,0,83,0,196,0,36,0,0,0,151,0,129,0,0,0,157,0,246,0,0,0,0,0,23,0,54,0,238,0,154,0,198,0,48,0,10,0,254,0,158,0,0,0,0,0,147,0,150,0,0,0,151,0,115,0,132,0,0,0,153,0,111,0,133,0,216,0,229,0,43,0,102,0,107,0,0,0,110,0,202,0,157,0,47,0,178,0,107,0,169,0,94,0,173,0,34,0,0,0,0,0,126,0,168,0,176,0,0,0,10,0,48,0,0,0,0,0,98,0,100,0,27,0,123,0,99,0,89,0,143,0,129,0,221,0,90,0,68,0,130,0,122,0,0,0,196,0,139,0,235,0,91,0,33,0,88,0,0,0,201,0,149,0,125,0,9,0,0,0,0,0,0,0,132,0,157,0,75,0,92,0,143,0,51,0,117,0,237,0,0,0,0,0,133,0,0,0,10,0,109,0,241,0,228,0,255,0,245,0,52,0,37,0,145,0,151,0,0,0,20,0,0,0,117,0,253,0,58,0,151,0,71,0,0,0,220,0,124,0,0,0,61,0,90,0,78,0,0,0,0,0,191,0,62,0,0,0,93,0,30,0,199,0,200,0,241,0,79,0,121,0,138,0,62,0,0,0,0,0,0,0,15,0,232,0,26,0,97,0,205,0,2,0,100,0,248,0,0,0,28,0,66,0,146,0,204,0,0,0,67,0,145,0,32,0,125,0,88,0,173,0,43,0,252,0,38,0,168,0,125,0,41,0,0,0,0,0,0,0,15,0,148,0,125,0,112,0,129,0,235,0,155,0,63,0,249,0,160,0,0,0,0,0,0,0,0,0,0,0,120,0,0,0,0,0,0,0,30,0,0,0,175,0,139,0,161,0,179,0,106,0,134,0,205,0,232,0,58,0,226,0,90,0,0,0,108,0,0,0,157,0,0,0,79,0,136,0,242,0,68,0,124,0,0,0,0,0,18,0,239,0,52,0,166,0,105,0,67,0,122,0,0,0,63,0,214,0,31,0,64,0,0,0,0,0,81,0,136,0,15,0,234,0,119,0,6,0,29,0,42,0,71,0,198,0,248,0,0,0,0,0,31,0,71,0,0,0,128,0,125,0,0,0,229,0,2,0,150,0,201,0,176,0,244,0,16,0,117,0,252,0,157,0,181,0,210,0,155,0,161,0,31,0,204,0,109,0,175,0,226,0,216,0,193,0,0,0,81,0,0,0,0,0,27,0,66,0,151,0,53,0,224,0,140,0,8,0,214,0,245,0,188,0,136,0,9,0,138,0,186,0,210,0,22,0,164,0,210,0,152,0,77,0,255,0,180,0,5,0,160,0,191,0,0,0,59,0,233,0,88,0,221,0,26,0,90,0,0,0,0,0,108,0,248,0,51,0,120,0,188,0,0,0,188,0,0,0,33,0,206,0,188,0,240,0,163,0,184,0,37,0,240,0,144,0,108,0,0,0,17,0,141,0,31,0,138,0,202,0,44,0,0,0,0,0,10,0,128,0,250,0,60,0,185,0,0,0,156,0,230,0,174,0,172,0,0,0,227,0,95,0,114,0,3,0,0,0,121,0,162,0,0,0,0,0,123,0,0,0,57,0,0,0,0,0,114,0,146,0,0,0,114,0,221,0,0,0,222,0,161,0,20,0,0,0,204,0,0,0,111,0,240,0,0,0,176,0,200,0,140,0,140,0,132,0,0,0,65,0,77,0,109,0,102,0,0,0,182,0,202,0,124,0,21,0,0,0,47,0,20,0,104,0,2,0,160,0,175,0,168,0,162,0,140,0,235,0,55,0,34,0,9,0,181,0,204,0,0,0,214,0,198,0,61,0,183,0,138,0,0,0,0,0,213,0,167,0,199,0,0,0,144,0,240,0,0,0,0,0,124,0,77,0,85,0,206,0,246,0,242,0,213,0,0,0,22,0,101,0,37,0,110,0,20,0,102,0,123,0,0,0,38,0,249,0,200,0,0,0,0,0,139,0);
signal scenario_full  : scenario_type := (223,31,48,31,48,30,89,31,73,31,89,31,80,31,188,31,47,31,121,31,114,31,114,30,245,31,207,31,186,31,22,31,4,31,4,30,103,31,202,31,109,31,60,31,32,31,78,31,129,31,14,31,76,31,184,31,230,31,243,31,243,30,76,31,62,31,135,31,103,31,103,30,203,31,178,31,136,31,169,31,169,30,94,31,17,31,17,30,9,31,56,31,56,30,199,31,196,31,196,30,196,29,32,31,90,31,107,31,112,31,26,31,113,31,113,30,230,31,230,30,179,31,12,31,249,31,25,31,146,31,69,31,39,31,83,31,196,31,36,31,36,30,151,31,129,31,129,30,157,31,246,31,246,30,246,29,23,31,54,31,238,31,154,31,198,31,48,31,10,31,254,31,158,31,158,30,158,29,147,31,150,31,150,30,151,31,115,31,132,31,132,30,153,31,111,31,133,31,216,31,229,31,43,31,102,31,107,31,107,30,110,31,202,31,157,31,47,31,178,31,107,31,169,31,94,31,173,31,34,31,34,30,34,29,126,31,168,31,176,31,176,30,10,31,48,31,48,30,48,29,98,31,100,31,27,31,123,31,99,31,89,31,143,31,129,31,221,31,90,31,68,31,130,31,122,31,122,30,196,31,139,31,235,31,91,31,33,31,88,31,88,30,201,31,149,31,125,31,9,31,9,30,9,29,9,28,132,31,157,31,75,31,92,31,143,31,51,31,117,31,237,31,237,30,237,29,133,31,133,30,10,31,109,31,241,31,228,31,255,31,245,31,52,31,37,31,145,31,151,31,151,30,20,31,20,30,117,31,253,31,58,31,151,31,71,31,71,30,220,31,124,31,124,30,61,31,90,31,78,31,78,30,78,29,191,31,62,31,62,30,93,31,30,31,199,31,200,31,241,31,79,31,121,31,138,31,62,31,62,30,62,29,62,28,15,31,232,31,26,31,97,31,205,31,2,31,100,31,248,31,248,30,28,31,66,31,146,31,204,31,204,30,67,31,145,31,32,31,125,31,88,31,173,31,43,31,252,31,38,31,168,31,125,31,41,31,41,30,41,29,41,28,15,31,148,31,125,31,112,31,129,31,235,31,155,31,63,31,249,31,160,31,160,30,160,29,160,28,160,27,160,26,120,31,120,30,120,29,120,28,30,31,30,30,175,31,139,31,161,31,179,31,106,31,134,31,205,31,232,31,58,31,226,31,90,31,90,30,108,31,108,30,157,31,157,30,79,31,136,31,242,31,68,31,124,31,124,30,124,29,18,31,239,31,52,31,166,31,105,31,67,31,122,31,122,30,63,31,214,31,31,31,64,31,64,30,64,29,81,31,136,31,15,31,234,31,119,31,6,31,29,31,42,31,71,31,198,31,248,31,248,30,248,29,31,31,71,31,71,30,128,31,125,31,125,30,229,31,2,31,150,31,201,31,176,31,244,31,16,31,117,31,252,31,157,31,181,31,210,31,155,31,161,31,31,31,204,31,109,31,175,31,226,31,216,31,193,31,193,30,81,31,81,30,81,29,27,31,66,31,151,31,53,31,224,31,140,31,8,31,214,31,245,31,188,31,136,31,9,31,138,31,186,31,210,31,22,31,164,31,210,31,152,31,77,31,255,31,180,31,5,31,160,31,191,31,191,30,59,31,233,31,88,31,221,31,26,31,90,31,90,30,90,29,108,31,248,31,51,31,120,31,188,31,188,30,188,31,188,30,33,31,206,31,188,31,240,31,163,31,184,31,37,31,240,31,144,31,108,31,108,30,17,31,141,31,31,31,138,31,202,31,44,31,44,30,44,29,10,31,128,31,250,31,60,31,185,31,185,30,156,31,230,31,174,31,172,31,172,30,227,31,95,31,114,31,3,31,3,30,121,31,162,31,162,30,162,29,123,31,123,30,57,31,57,30,57,29,114,31,146,31,146,30,114,31,221,31,221,30,222,31,161,31,20,31,20,30,204,31,204,30,111,31,240,31,240,30,176,31,200,31,140,31,140,31,132,31,132,30,65,31,77,31,109,31,102,31,102,30,182,31,202,31,124,31,21,31,21,30,47,31,20,31,104,31,2,31,160,31,175,31,168,31,162,31,140,31,235,31,55,31,34,31,9,31,181,31,204,31,204,30,214,31,198,31,61,31,183,31,138,31,138,30,138,29,213,31,167,31,199,31,199,30,144,31,240,31,240,30,240,29,124,31,77,31,85,31,206,31,246,31,242,31,213,31,213,30,22,31,101,31,37,31,110,31,20,31,102,31,123,31,123,30,38,31,249,31,200,31,200,30,200,29,139,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
