-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 745;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (135,0,0,0,0,0,55,0,36,0,210,0,6,0,206,0,0,0,35,0,102,0,156,0,124,0,167,0,253,0,251,0,195,0,95,0,0,0,0,0,25,0,137,0,159,0,80,0,88,0,163,0,138,0,102,0,69,0,91,0,89,0,79,0,0,0,18,0,120,0,128,0,79,0,0,0,137,0,220,0,0,0,88,0,89,0,56,0,186,0,181,0,0,0,0,0,250,0,0,0,0,0,0,0,13,0,210,0,226,0,196,0,85,0,100,0,248,0,146,0,58,0,240,0,202,0,84,0,86,0,85,0,0,0,125,0,88,0,0,0,57,0,144,0,70,0,159,0,255,0,0,0,2,0,25,0,181,0,139,0,0,0,0,0,106,0,38,0,47,0,95,0,233,0,145,0,0,0,142,0,229,0,110,0,162,0,61,0,0,0,0,0,0,0,181,0,79,0,156,0,0,0,0,0,86,0,193,0,43,0,0,0,195,0,61,0,147,0,0,0,252,0,0,0,249,0,0,0,0,0,239,0,0,0,222,0,172,0,116,0,0,0,34,0,161,0,0,0,27,0,18,0,0,0,1,0,0,0,0,0,190,0,178,0,97,0,163,0,0,0,36,0,129,0,162,0,105,0,108,0,157,0,0,0,42,0,251,0,114,0,163,0,97,0,36,0,0,0,235,0,144,0,213,0,130,0,89,0,54,0,200,0,234,0,0,0,236,0,0,0,64,0,0,0,0,0,230,0,0,0,0,0,160,0,221,0,144,0,0,0,106,0,0,0,37,0,75,0,77,0,212,0,192,0,247,0,0,0,184,0,117,0,44,0,223,0,112,0,195,0,142,0,0,0,162,0,43,0,181,0,0,0,202,0,76,0,4,0,39,0,20,0,60,0,183,0,180,0,17,0,37,0,143,0,52,0,155,0,250,0,239,0,190,0,229,0,179,0,244,0,0,0,0,0,44,0,160,0,169,0,158,0,0,0,252,0,176,0,49,0,94,0,116,0,244,0,38,0,183,0,66,0,92,0,0,0,227,0,180,0,108,0,207,0,152,0,159,0,13,0,95,0,188,0,175,0,81,0,103,0,250,0,107,0,4,0,193,0,0,0,54,0,219,0,0,0,191,0,18,0,247,0,0,0,0,0,166,0,155,0,0,0,102,0,52,0,130,0,0,0,39,0,115,0,208,0,124,0,114,0,0,0,0,0,75,0,0,0,212,0,67,0,116,0,14,0,0,0,0,0,99,0,82,0,248,0,158,0,178,0,115,0,117,0,89,0,141,0,238,0,19,0,179,0,248,0,0,0,121,0,23,0,184,0,0,0,215,0,70,0,254,0,17,0,0,0,214,0,221,0,0,0,206,0,0,0,0,0,224,0,0,0,51,0,7,0,3,0,118,0,235,0,229,0,196,0,85,0,193,0,77,0,153,0,184,0,240,0,156,0,221,0,209,0,204,0,231,0,92,0,0,0,79,0,110,0,0,0,246,0,107,0,208,0,151,0,0,0,206,0,148,0,124,0,58,0,105,0,185,0,163,0,158,0,0,0,215,0,0,0,169,0,34,0,0,0,106,0,111,0,49,0,205,0,57,0,69,0,188,0,0,0,237,0,156,0,111,0,0,0,146,0,183,0,78,0,184,0,186,0,92,0,0,0,16,0,214,0,0,0,0,0,249,0,0,0,199,0,228,0,168,0,0,0,197,0,0,0,203,0,22,0,154,0,222,0,39,0,0,0,217,0,237,0,0,0,26,0,41,0,33,0,17,0,238,0,0,0,173,0,82,0,141,0,64,0,164,0,42,0,223,0,217,0,0,0,0,0,81,0,0,0,89,0,0,0,119,0,45,0,116,0,78,0,135,0,0,0,0,0,154,0,0,0,145,0,0,0,223,0,0,0,92,0,231,0,239,0,202,0,71,0,21,0,82,0,165,0,210,0,244,0,0,0,1,0,0,0,198,0,230,0,96,0,0,0,0,0,245,0,84,0,29,0,0,0,176,0,193,0,106,0,232,0,249,0,127,0,184,0,0,0,0,0,118,0,61,0,235,0,245,0,29,0,199,0,33,0,16,0,0,0,146,0,0,0,101,0,245,0,56,0,226,0,1,0,30,0,243,0,164,0,198,0,11,0,130,0,8,0,192,0,206,0,133,0,247,0,35,0,0,0,79,0,113,0,186,0,85,0,169,0,169,0,231,0,60,0,251,0,82,0,142,0,155,0,0,0,63,0,115,0,46,0,0,0,162,0,148,0,29,0,203,0,147,0,234,0,83,0,108,0,0,0,0,0,177,0,251,0,171,0,120,0,0,0,231,0,147,0,0,0,120,0,65,0,101,0,0,0,0,0,5,0,14,0,0,0,4,0,139,0,231,0,112,0,0,0,0,0,38,0,171,0,44,0,0,0,253,0,184,0,126,0,60,0,0,0,198,0,120,0,60,0,130,0,41,0,49,0,61,0,247,0,68,0,0,0,0,0,51,0,150,0,133,0,156,0,117,0,116,0,67,0,164,0,139,0,39,0,218,0,134,0,149,0,24,0,239,0,24,0,0,0,21,0,40,0,0,0,191,0,99,0,0,0,13,0,0,0,183,0,220,0,0,0,225,0,0,0,2,0,210,0,176,0,0,0,236,0,106,0,87,0,108,0,172,0,65,0,88,0,3,0,90,0,171,0,1,0,61,0,59,0,11,0,57,0,0,0,81,0,0,0,0,0,90,0,0,0,74,0,0,0,17,0,51,0,137,0,234,0,219,0,0,0,0,0,31,0,61,0,214,0,37,0,202,0,216,0,0,0,0,0,237,0,96,0,0,0,125,0,0,0,45,0,0,0,156,0,210,0,41,0,12,0,98,0,59,0,145,0,197,0,230,0,234,0,116,0,95,0,8,0,88,0,52,0,247,0,0,0,15,0,97,0,145,0,85,0,0,0,90,0,0,0,133,0,116,0,179,0,122,0,120,0,243,0,15,0,51,0,0,0,23,0,201,0,249,0,103,0,51,0,157,0,0,0,179,0,147,0,31,0,84,0,216,0,93,0,153,0,0,0,0,0,241,0,157,0,23,0,128,0,0,0,44,0,63,0,30,0,83,0,162,0,0,0,48,0,101,0,189,0,0,0,231,0,212,0,100,0,0,0,100,0,205,0,136,0,219,0,57,0,252,0,108,0,0,0,0,0,0,0,65,0,153,0,26,0,105,0,0,0,114,0,39,0,0,0,143,0,21,0,10,0,52,0,217,0,180,0,169,0,190,0,207,0,165,0,141,0,105,0,25,0,12,0,142,0,27,0,176,0,135,0,120,0,17,0,142,0,39,0,0,0,12,0,120,0,0,0,143,0,114,0,37,0,0,0);
signal scenario_full  : scenario_type := (135,31,135,30,135,29,55,31,36,31,210,31,6,31,206,31,206,30,35,31,102,31,156,31,124,31,167,31,253,31,251,31,195,31,95,31,95,30,95,29,25,31,137,31,159,31,80,31,88,31,163,31,138,31,102,31,69,31,91,31,89,31,79,31,79,30,18,31,120,31,128,31,79,31,79,30,137,31,220,31,220,30,88,31,89,31,56,31,186,31,181,31,181,30,181,29,250,31,250,30,250,29,250,28,13,31,210,31,226,31,196,31,85,31,100,31,248,31,146,31,58,31,240,31,202,31,84,31,86,31,85,31,85,30,125,31,88,31,88,30,57,31,144,31,70,31,159,31,255,31,255,30,2,31,25,31,181,31,139,31,139,30,139,29,106,31,38,31,47,31,95,31,233,31,145,31,145,30,142,31,229,31,110,31,162,31,61,31,61,30,61,29,61,28,181,31,79,31,156,31,156,30,156,29,86,31,193,31,43,31,43,30,195,31,61,31,147,31,147,30,252,31,252,30,249,31,249,30,249,29,239,31,239,30,222,31,172,31,116,31,116,30,34,31,161,31,161,30,27,31,18,31,18,30,1,31,1,30,1,29,190,31,178,31,97,31,163,31,163,30,36,31,129,31,162,31,105,31,108,31,157,31,157,30,42,31,251,31,114,31,163,31,97,31,36,31,36,30,235,31,144,31,213,31,130,31,89,31,54,31,200,31,234,31,234,30,236,31,236,30,64,31,64,30,64,29,230,31,230,30,230,29,160,31,221,31,144,31,144,30,106,31,106,30,37,31,75,31,77,31,212,31,192,31,247,31,247,30,184,31,117,31,44,31,223,31,112,31,195,31,142,31,142,30,162,31,43,31,181,31,181,30,202,31,76,31,4,31,39,31,20,31,60,31,183,31,180,31,17,31,37,31,143,31,52,31,155,31,250,31,239,31,190,31,229,31,179,31,244,31,244,30,244,29,44,31,160,31,169,31,158,31,158,30,252,31,176,31,49,31,94,31,116,31,244,31,38,31,183,31,66,31,92,31,92,30,227,31,180,31,108,31,207,31,152,31,159,31,13,31,95,31,188,31,175,31,81,31,103,31,250,31,107,31,4,31,193,31,193,30,54,31,219,31,219,30,191,31,18,31,247,31,247,30,247,29,166,31,155,31,155,30,102,31,52,31,130,31,130,30,39,31,115,31,208,31,124,31,114,31,114,30,114,29,75,31,75,30,212,31,67,31,116,31,14,31,14,30,14,29,99,31,82,31,248,31,158,31,178,31,115,31,117,31,89,31,141,31,238,31,19,31,179,31,248,31,248,30,121,31,23,31,184,31,184,30,215,31,70,31,254,31,17,31,17,30,214,31,221,31,221,30,206,31,206,30,206,29,224,31,224,30,51,31,7,31,3,31,118,31,235,31,229,31,196,31,85,31,193,31,77,31,153,31,184,31,240,31,156,31,221,31,209,31,204,31,231,31,92,31,92,30,79,31,110,31,110,30,246,31,107,31,208,31,151,31,151,30,206,31,148,31,124,31,58,31,105,31,185,31,163,31,158,31,158,30,215,31,215,30,169,31,34,31,34,30,106,31,111,31,49,31,205,31,57,31,69,31,188,31,188,30,237,31,156,31,111,31,111,30,146,31,183,31,78,31,184,31,186,31,92,31,92,30,16,31,214,31,214,30,214,29,249,31,249,30,199,31,228,31,168,31,168,30,197,31,197,30,203,31,22,31,154,31,222,31,39,31,39,30,217,31,237,31,237,30,26,31,41,31,33,31,17,31,238,31,238,30,173,31,82,31,141,31,64,31,164,31,42,31,223,31,217,31,217,30,217,29,81,31,81,30,89,31,89,30,119,31,45,31,116,31,78,31,135,31,135,30,135,29,154,31,154,30,145,31,145,30,223,31,223,30,92,31,231,31,239,31,202,31,71,31,21,31,82,31,165,31,210,31,244,31,244,30,1,31,1,30,198,31,230,31,96,31,96,30,96,29,245,31,84,31,29,31,29,30,176,31,193,31,106,31,232,31,249,31,127,31,184,31,184,30,184,29,118,31,61,31,235,31,245,31,29,31,199,31,33,31,16,31,16,30,146,31,146,30,101,31,245,31,56,31,226,31,1,31,30,31,243,31,164,31,198,31,11,31,130,31,8,31,192,31,206,31,133,31,247,31,35,31,35,30,79,31,113,31,186,31,85,31,169,31,169,31,231,31,60,31,251,31,82,31,142,31,155,31,155,30,63,31,115,31,46,31,46,30,162,31,148,31,29,31,203,31,147,31,234,31,83,31,108,31,108,30,108,29,177,31,251,31,171,31,120,31,120,30,231,31,147,31,147,30,120,31,65,31,101,31,101,30,101,29,5,31,14,31,14,30,4,31,139,31,231,31,112,31,112,30,112,29,38,31,171,31,44,31,44,30,253,31,184,31,126,31,60,31,60,30,198,31,120,31,60,31,130,31,41,31,49,31,61,31,247,31,68,31,68,30,68,29,51,31,150,31,133,31,156,31,117,31,116,31,67,31,164,31,139,31,39,31,218,31,134,31,149,31,24,31,239,31,24,31,24,30,21,31,40,31,40,30,191,31,99,31,99,30,13,31,13,30,183,31,220,31,220,30,225,31,225,30,2,31,210,31,176,31,176,30,236,31,106,31,87,31,108,31,172,31,65,31,88,31,3,31,90,31,171,31,1,31,61,31,59,31,11,31,57,31,57,30,81,31,81,30,81,29,90,31,90,30,74,31,74,30,17,31,51,31,137,31,234,31,219,31,219,30,219,29,31,31,61,31,214,31,37,31,202,31,216,31,216,30,216,29,237,31,96,31,96,30,125,31,125,30,45,31,45,30,156,31,210,31,41,31,12,31,98,31,59,31,145,31,197,31,230,31,234,31,116,31,95,31,8,31,88,31,52,31,247,31,247,30,15,31,97,31,145,31,85,31,85,30,90,31,90,30,133,31,116,31,179,31,122,31,120,31,243,31,15,31,51,31,51,30,23,31,201,31,249,31,103,31,51,31,157,31,157,30,179,31,147,31,31,31,84,31,216,31,93,31,153,31,153,30,153,29,241,31,157,31,23,31,128,31,128,30,44,31,63,31,30,31,83,31,162,31,162,30,48,31,101,31,189,31,189,30,231,31,212,31,100,31,100,30,100,31,205,31,136,31,219,31,57,31,252,31,108,31,108,30,108,29,108,28,65,31,153,31,26,31,105,31,105,30,114,31,39,31,39,30,143,31,21,31,10,31,52,31,217,31,180,31,169,31,190,31,207,31,165,31,141,31,105,31,25,31,12,31,142,31,27,31,176,31,135,31,120,31,17,31,142,31,39,31,39,30,12,31,120,31,120,30,143,31,114,31,37,31,37,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
