-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 765;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (120,0,0,0,191,0,0,0,159,0,183,0,241,0,0,0,0,0,0,0,18,0,209,0,32,0,30,0,245,0,48,0,217,0,0,0,0,0,118,0,252,0,213,0,92,0,237,0,113,0,204,0,42,0,254,0,0,0,0,0,59,0,130,0,2,0,147,0,0,0,91,0,0,0,0,0,200,0,190,0,168,0,0,0,182,0,0,0,123,0,55,0,0,0,157,0,49,0,246,0,224,0,61,0,254,0,77,0,101,0,0,0,137,0,87,0,252,0,20,0,30,0,73,0,131,0,154,0,0,0,110,0,87,0,221,0,253,0,238,0,0,0,0,0,108,0,214,0,217,0,48,0,0,0,3,0,175,0,116,0,211,0,204,0,10,0,32,0,0,0,0,0,0,0,118,0,0,0,0,0,66,0,35,0,190,0,96,0,151,0,96,0,49,0,182,0,53,0,46,0,250,0,200,0,179,0,0,0,187,0,96,0,0,0,164,0,0,0,70,0,199,0,23,0,111,0,208,0,161,0,131,0,0,0,11,0,180,0,55,0,0,0,112,0,0,0,154,0,8,0,237,0,211,0,107,0,143,0,13,0,0,0,130,0,0,0,2,0,58,0,4,0,110,0,27,0,91,0,134,0,196,0,158,0,67,0,45,0,28,0,211,0,128,0,126,0,63,0,232,0,241,0,4,0,59,0,105,0,215,0,119,0,139,0,32,0,168,0,1,0,103,0,0,0,93,0,241,0,189,0,27,0,255,0,101,0,182,0,0,0,53,0,6,0,85,0,24,0,159,0,50,0,17,0,238,0,40,0,0,0,0,0,145,0,133,0,64,0,206,0,0,0,35,0,163,0,150,0,31,0,21,0,0,0,0,0,82,0,218,0,146,0,103,0,242,0,196,0,242,0,0,0,109,0,28,0,68,0,129,0,16,0,0,0,216,0,4,0,211,0,88,0,242,0,251,0,206,0,36,0,77,0,0,0,112,0,0,0,64,0,231,0,36,0,151,0,32,0,10,0,157,0,251,0,136,0,0,0,245,0,123,0,80,0,211,0,64,0,0,0,103,0,89,0,228,0,211,0,71,0,222,0,0,0,142,0,0,0,188,0,0,0,81,0,0,0,175,0,189,0,195,0,0,0,0,0,135,0,40,0,0,0,29,0,9,0,58,0,5,0,219,0,143,0,102,0,15,0,220,0,250,0,246,0,0,0,125,0,0,0,102,0,235,0,91,0,89,0,111,0,0,0,122,0,0,0,222,0,108,0,85,0,0,0,0,0,38,0,57,0,87,0,204,0,36,0,139,0,166,0,24,0,0,0,118,0,238,0,0,0,248,0,242,0,68,0,32,0,0,0,0,0,169,0,52,0,6,0,252,0,80,0,100,0,210,0,111,0,59,0,3,0,0,0,109,0,0,0,116,0,112,0,0,0,160,0,215,0,0,0,190,0,255,0,184,0,232,0,193,0,199,0,236,0,44,0,29,0,64,0,101,0,24,0,234,0,0,0,192,0,163,0,87,0,88,0,0,0,196,0,227,0,174,0,133,0,86,0,194,0,0,0,203,0,10,0,41,0,0,0,200,0,86,0,14,0,117,0,228,0,0,0,24,0,40,0,16,0,255,0,128,0,112,0,218,0,0,0,95,0,124,0,0,0,214,0,0,0,63,0,136,0,91,0,156,0,185,0,29,0,0,0,181,0,105,0,150,0,235,0,33,0,68,0,85,0,203,0,103,0,147,0,0,0,152,0,107,0,0,0,55,0,49,0,31,0,71,0,176,0,0,0,238,0,95,0,81,0,195,0,0,0,99,0,0,0,0,0,131,0,0,0,138,0,163,0,245,0,241,0,12,0,0,0,127,0,80,0,177,0,129,0,96,0,76,0,0,0,84,0,0,0,125,0,158,0,0,0,202,0,137,0,231,0,243,0,119,0,0,0,212,0,0,0,224,0,158,0,228,0,181,0,83,0,240,0,86,0,119,0,44,0,175,0,249,0,69,0,133,0,197,0,5,0,0,0,77,0,0,0,98,0,182,0,204,0,0,0,0,0,0,0,164,0,167,0,24,0,183,0,134,0,69,0,162,0,34,0,188,0,40,0,0,0,25,0,105,0,0,0,0,0,9,0,45,0,50,0,215,0,165,0,228,0,230,0,112,0,21,0,187,0,0,0,66,0,15,0,0,0,156,0,31,0,79,0,0,0,218,0,0,0,145,0,153,0,21,0,118,0,109,0,30,0,174,0,147,0,28,0,197,0,0,0,232,0,172,0,166,0,245,0,119,0,87,0,175,0,100,0,78,0,0,0,110,0,0,0,249,0,243,0,0,0,201,0,150,0,235,0,65,0,228,0,80,0,101,0,226,0,0,0,214,0,141,0,205,0,66,0,211,0,24,0,126,0,62,0,10,0,0,0,57,0,0,0,0,0,107,0,0,0,246,0,86,0,209,0,142,0,218,0,251,0,254,0,189,0,253,0,114,0,157,0,0,0,146,0,133,0,0,0,0,0,149,0,74,0,25,0,0,0,175,0,54,0,156,0,0,0,0,0,131,0,79,0,0,0,149,0,49,0,217,0,95,0,21,0,87,0,236,0,214,0,72,0,0,0,36,0,78,0,177,0,184,0,0,0,159,0,248,0,0,0,0,0,205,0,19,0,219,0,0,0,42,0,0,0,254,0,90,0,32,0,72,0,40,0,45,0,216,0,162,0,53,0,73,0,45,0,0,0,147,0,101,0,143,0,88,0,155,0,162,0,86,0,134,0,36,0,0,0,0,0,13,0,144,0,83,0,8,0,8,0,0,0,179,0,226,0,165,0,91,0,0,0,195,0,120,0,53,0,41,0,118,0,214,0,191,0,160,0,229,0,0,0,13,0,0,0,230,0,0,0,0,0,194,0,1,0,116,0,137,0,157,0,129,0,66,0,191,0,254,0,0,0,62,0,86,0,205,0,127,0,147,0,21,0,238,0,139,0,241,0,77,0,43,0,48,0,46,0,18,0,108,0,116,0,199,0,170,0,220,0,129,0,78,0,0,0,0,0,47,0,185,0,238,0,10,0,86,0,0,0,83,0,238,0,155,0,0,0,195,0,109,0,236,0,93,0,4,0,25,0,202,0,134,0,0,0,121,0,105,0,240,0,0,0,153,0,64,0,44,0,0,0,1,0,198,0,198,0,34,0,163,0,154,0,25,0,44,0,156,0,108,0,0,0,144,0,72,0,167,0,59,0,0,0,48,0,66,0,196,0,50,0,241,0,91,0,177,0,0,0,189,0,49,0,106,0,133,0,156,0,174,0,229,0,63,0,0,0,0,0,239,0,152,0,91,0,0,0,175,0,24,0,82,0,114,0,230,0,0,0,64,0,91,0,110,0,111,0,66,0,9,0,215,0,204,0,203,0,0,0,131,0,212,0,225,0,0,0,197,0,168,0,120,0,219,0);
signal scenario_full  : scenario_type := (120,31,120,30,191,31,191,30,159,31,183,31,241,31,241,30,241,29,241,28,18,31,209,31,32,31,30,31,245,31,48,31,217,31,217,30,217,29,118,31,252,31,213,31,92,31,237,31,113,31,204,31,42,31,254,31,254,30,254,29,59,31,130,31,2,31,147,31,147,30,91,31,91,30,91,29,200,31,190,31,168,31,168,30,182,31,182,30,123,31,55,31,55,30,157,31,49,31,246,31,224,31,61,31,254,31,77,31,101,31,101,30,137,31,87,31,252,31,20,31,30,31,73,31,131,31,154,31,154,30,110,31,87,31,221,31,253,31,238,31,238,30,238,29,108,31,214,31,217,31,48,31,48,30,3,31,175,31,116,31,211,31,204,31,10,31,32,31,32,30,32,29,32,28,118,31,118,30,118,29,66,31,35,31,190,31,96,31,151,31,96,31,49,31,182,31,53,31,46,31,250,31,200,31,179,31,179,30,187,31,96,31,96,30,164,31,164,30,70,31,199,31,23,31,111,31,208,31,161,31,131,31,131,30,11,31,180,31,55,31,55,30,112,31,112,30,154,31,8,31,237,31,211,31,107,31,143,31,13,31,13,30,130,31,130,30,2,31,58,31,4,31,110,31,27,31,91,31,134,31,196,31,158,31,67,31,45,31,28,31,211,31,128,31,126,31,63,31,232,31,241,31,4,31,59,31,105,31,215,31,119,31,139,31,32,31,168,31,1,31,103,31,103,30,93,31,241,31,189,31,27,31,255,31,101,31,182,31,182,30,53,31,6,31,85,31,24,31,159,31,50,31,17,31,238,31,40,31,40,30,40,29,145,31,133,31,64,31,206,31,206,30,35,31,163,31,150,31,31,31,21,31,21,30,21,29,82,31,218,31,146,31,103,31,242,31,196,31,242,31,242,30,109,31,28,31,68,31,129,31,16,31,16,30,216,31,4,31,211,31,88,31,242,31,251,31,206,31,36,31,77,31,77,30,112,31,112,30,64,31,231,31,36,31,151,31,32,31,10,31,157,31,251,31,136,31,136,30,245,31,123,31,80,31,211,31,64,31,64,30,103,31,89,31,228,31,211,31,71,31,222,31,222,30,142,31,142,30,188,31,188,30,81,31,81,30,175,31,189,31,195,31,195,30,195,29,135,31,40,31,40,30,29,31,9,31,58,31,5,31,219,31,143,31,102,31,15,31,220,31,250,31,246,31,246,30,125,31,125,30,102,31,235,31,91,31,89,31,111,31,111,30,122,31,122,30,222,31,108,31,85,31,85,30,85,29,38,31,57,31,87,31,204,31,36,31,139,31,166,31,24,31,24,30,118,31,238,31,238,30,248,31,242,31,68,31,32,31,32,30,32,29,169,31,52,31,6,31,252,31,80,31,100,31,210,31,111,31,59,31,3,31,3,30,109,31,109,30,116,31,112,31,112,30,160,31,215,31,215,30,190,31,255,31,184,31,232,31,193,31,199,31,236,31,44,31,29,31,64,31,101,31,24,31,234,31,234,30,192,31,163,31,87,31,88,31,88,30,196,31,227,31,174,31,133,31,86,31,194,31,194,30,203,31,10,31,41,31,41,30,200,31,86,31,14,31,117,31,228,31,228,30,24,31,40,31,16,31,255,31,128,31,112,31,218,31,218,30,95,31,124,31,124,30,214,31,214,30,63,31,136,31,91,31,156,31,185,31,29,31,29,30,181,31,105,31,150,31,235,31,33,31,68,31,85,31,203,31,103,31,147,31,147,30,152,31,107,31,107,30,55,31,49,31,31,31,71,31,176,31,176,30,238,31,95,31,81,31,195,31,195,30,99,31,99,30,99,29,131,31,131,30,138,31,163,31,245,31,241,31,12,31,12,30,127,31,80,31,177,31,129,31,96,31,76,31,76,30,84,31,84,30,125,31,158,31,158,30,202,31,137,31,231,31,243,31,119,31,119,30,212,31,212,30,224,31,158,31,228,31,181,31,83,31,240,31,86,31,119,31,44,31,175,31,249,31,69,31,133,31,197,31,5,31,5,30,77,31,77,30,98,31,182,31,204,31,204,30,204,29,204,28,164,31,167,31,24,31,183,31,134,31,69,31,162,31,34,31,188,31,40,31,40,30,25,31,105,31,105,30,105,29,9,31,45,31,50,31,215,31,165,31,228,31,230,31,112,31,21,31,187,31,187,30,66,31,15,31,15,30,156,31,31,31,79,31,79,30,218,31,218,30,145,31,153,31,21,31,118,31,109,31,30,31,174,31,147,31,28,31,197,31,197,30,232,31,172,31,166,31,245,31,119,31,87,31,175,31,100,31,78,31,78,30,110,31,110,30,249,31,243,31,243,30,201,31,150,31,235,31,65,31,228,31,80,31,101,31,226,31,226,30,214,31,141,31,205,31,66,31,211,31,24,31,126,31,62,31,10,31,10,30,57,31,57,30,57,29,107,31,107,30,246,31,86,31,209,31,142,31,218,31,251,31,254,31,189,31,253,31,114,31,157,31,157,30,146,31,133,31,133,30,133,29,149,31,74,31,25,31,25,30,175,31,54,31,156,31,156,30,156,29,131,31,79,31,79,30,149,31,49,31,217,31,95,31,21,31,87,31,236,31,214,31,72,31,72,30,36,31,78,31,177,31,184,31,184,30,159,31,248,31,248,30,248,29,205,31,19,31,219,31,219,30,42,31,42,30,254,31,90,31,32,31,72,31,40,31,45,31,216,31,162,31,53,31,73,31,45,31,45,30,147,31,101,31,143,31,88,31,155,31,162,31,86,31,134,31,36,31,36,30,36,29,13,31,144,31,83,31,8,31,8,31,8,30,179,31,226,31,165,31,91,31,91,30,195,31,120,31,53,31,41,31,118,31,214,31,191,31,160,31,229,31,229,30,13,31,13,30,230,31,230,30,230,29,194,31,1,31,116,31,137,31,157,31,129,31,66,31,191,31,254,31,254,30,62,31,86,31,205,31,127,31,147,31,21,31,238,31,139,31,241,31,77,31,43,31,48,31,46,31,18,31,108,31,116,31,199,31,170,31,220,31,129,31,78,31,78,30,78,29,47,31,185,31,238,31,10,31,86,31,86,30,83,31,238,31,155,31,155,30,195,31,109,31,236,31,93,31,4,31,25,31,202,31,134,31,134,30,121,31,105,31,240,31,240,30,153,31,64,31,44,31,44,30,1,31,198,31,198,31,34,31,163,31,154,31,25,31,44,31,156,31,108,31,108,30,144,31,72,31,167,31,59,31,59,30,48,31,66,31,196,31,50,31,241,31,91,31,177,31,177,30,189,31,49,31,106,31,133,31,156,31,174,31,229,31,63,31,63,30,63,29,239,31,152,31,91,31,91,30,175,31,24,31,82,31,114,31,230,31,230,30,64,31,91,31,110,31,111,31,66,31,9,31,215,31,204,31,203,31,203,30,131,31,212,31,225,31,225,30,197,31,168,31,120,31,219,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
