-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 325;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (109,0,125,0,199,0,0,0,118,0,63,0,225,0,242,0,160,0,67,0,199,0,0,0,37,0,0,0,123,0,34,0,95,0,142,0,146,0,157,0,208,0,121,0,187,0,68,0,95,0,0,0,211,0,223,0,135,0,143,0,113,0,0,0,217,0,0,0,139,0,236,0,227,0,121,0,211,0,181,0,1,0,158,0,187,0,91,0,126,0,0,0,242,0,10,0,97,0,171,0,0,0,165,0,0,0,86,0,120,0,142,0,153,0,30,0,0,0,28,0,126,0,161,0,96,0,0,0,0,0,16,0,59,0,137,0,191,0,108,0,18,0,96,0,0,0,126,0,109,0,0,0,0,0,0,0,98,0,195,0,215,0,240,0,199,0,78,0,130,0,0,0,42,0,133,0,12,0,196,0,228,0,112,0,71,0,72,0,119,0,0,0,120,0,145,0,141,0,0,0,94,0,121,0,0,0,0,0,79,0,96,0,0,0,97,0,125,0,249,0,148,0,156,0,41,0,42,0,152,0,95,0,167,0,71,0,123,0,195,0,227,0,7,0,180,0,97,0,210,0,132,0,156,0,102,0,40,0,109,0,0,0,52,0,0,0,46,0,31,0,49,0,0,0,39,0,11,0,0,0,102,0,188,0,0,0,0,0,0,0,100,0,193,0,0,0,70,0,0,0,0,0,113,0,221,0,0,0,162,0,131,0,0,0,79,0,198,0,218,0,86,0,156,0,0,0,0,0,21,0,3,0,81,0,4,0,88,0,166,0,35,0,152,0,0,0,3,0,91,0,0,0,241,0,241,0,0,0,0,0,37,0,0,0,132,0,205,0,0,0,0,0,165,0,176,0,75,0,64,0,40,0,119,0,0,0,116,0,238,0,0,0,149,0,227,0,32,0,232,0,87,0,0,0,26,0,0,0,210,0,192,0,156,0,155,0,185,0,0,0,0,0,0,0,95,0,201,0,29,0,219,0,0,0,12,0,245,0,0,0,0,0,209,0,224,0,43,0,69,0,143,0,0,0,34,0,90,0,137,0,106,0,217,0,3,0,52,0,130,0,0,0,85,0,227,0,61,0,205,0,40,0,59,0,132,0,224,0,0,0,135,0,111,0,41,0,0,0,78,0,2,0,208,0,170,0,87,0,203,0,180,0,89,0,140,0,0,0,0,0,164,0,131,0,14,0,205,0,60,0,126,0,84,0,0,0,22,0,0,0,75,0,200,0,128,0,206,0,155,0,251,0,143,0,1,0,5,0,128,0,0,0,239,0,0,0,186,0,27,0,252,0,77,0,0,0,122,0,200,0,8,0,177,0,166,0,190,0,195,0,136,0,217,0,158,0,76,0,105,0,102,0,0,0,83,0,34,0,0,0,0,0,80,0,9,0,140,0,0,0,100,0,21,0,214,0,70,0,75,0,228,0,0,0,203,0,141,0,187,0,198,0,242,0,129,0,51,0,35,0);
signal scenario_full  : scenario_type := (109,31,125,31,199,31,199,30,118,31,63,31,225,31,242,31,160,31,67,31,199,31,199,30,37,31,37,30,123,31,34,31,95,31,142,31,146,31,157,31,208,31,121,31,187,31,68,31,95,31,95,30,211,31,223,31,135,31,143,31,113,31,113,30,217,31,217,30,139,31,236,31,227,31,121,31,211,31,181,31,1,31,158,31,187,31,91,31,126,31,126,30,242,31,10,31,97,31,171,31,171,30,165,31,165,30,86,31,120,31,142,31,153,31,30,31,30,30,28,31,126,31,161,31,96,31,96,30,96,29,16,31,59,31,137,31,191,31,108,31,18,31,96,31,96,30,126,31,109,31,109,30,109,29,109,28,98,31,195,31,215,31,240,31,199,31,78,31,130,31,130,30,42,31,133,31,12,31,196,31,228,31,112,31,71,31,72,31,119,31,119,30,120,31,145,31,141,31,141,30,94,31,121,31,121,30,121,29,79,31,96,31,96,30,97,31,125,31,249,31,148,31,156,31,41,31,42,31,152,31,95,31,167,31,71,31,123,31,195,31,227,31,7,31,180,31,97,31,210,31,132,31,156,31,102,31,40,31,109,31,109,30,52,31,52,30,46,31,31,31,49,31,49,30,39,31,11,31,11,30,102,31,188,31,188,30,188,29,188,28,100,31,193,31,193,30,70,31,70,30,70,29,113,31,221,31,221,30,162,31,131,31,131,30,79,31,198,31,218,31,86,31,156,31,156,30,156,29,21,31,3,31,81,31,4,31,88,31,166,31,35,31,152,31,152,30,3,31,91,31,91,30,241,31,241,31,241,30,241,29,37,31,37,30,132,31,205,31,205,30,205,29,165,31,176,31,75,31,64,31,40,31,119,31,119,30,116,31,238,31,238,30,149,31,227,31,32,31,232,31,87,31,87,30,26,31,26,30,210,31,192,31,156,31,155,31,185,31,185,30,185,29,185,28,95,31,201,31,29,31,219,31,219,30,12,31,245,31,245,30,245,29,209,31,224,31,43,31,69,31,143,31,143,30,34,31,90,31,137,31,106,31,217,31,3,31,52,31,130,31,130,30,85,31,227,31,61,31,205,31,40,31,59,31,132,31,224,31,224,30,135,31,111,31,41,31,41,30,78,31,2,31,208,31,170,31,87,31,203,31,180,31,89,31,140,31,140,30,140,29,164,31,131,31,14,31,205,31,60,31,126,31,84,31,84,30,22,31,22,30,75,31,200,31,128,31,206,31,155,31,251,31,143,31,1,31,5,31,128,31,128,30,239,31,239,30,186,31,27,31,252,31,77,31,77,30,122,31,200,31,8,31,177,31,166,31,190,31,195,31,136,31,217,31,158,31,76,31,105,31,102,31,102,30,83,31,34,31,34,30,34,29,80,31,9,31,140,31,140,30,100,31,21,31,214,31,70,31,75,31,228,31,228,30,203,31,141,31,187,31,198,31,242,31,129,31,51,31,35,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
