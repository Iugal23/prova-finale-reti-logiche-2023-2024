-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 866;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (134,0,158,0,54,0,176,0,154,0,71,0,163,0,141,0,178,0,156,0,8,0,0,0,9,0,181,0,247,0,9,0,142,0,152,0,114,0,166,0,238,0,179,0,0,0,16,0,245,0,18,0,0,0,38,0,114,0,180,0,243,0,0,0,0,0,13,0,234,0,126,0,165,0,139,0,119,0,178,0,238,0,165,0,0,0,0,0,228,0,20,0,245,0,186,0,151,0,241,0,242,0,122,0,217,0,214,0,170,0,0,0,202,0,219,0,0,0,190,0,246,0,196,0,0,0,176,0,158,0,175,0,182,0,171,0,0,0,100,0,6,0,166,0,0,0,5,0,199,0,0,0,92,0,40,0,107,0,90,0,35,0,206,0,6,0,135,0,96,0,119,0,0,0,96,0,60,0,151,0,153,0,226,0,247,0,234,0,31,0,187,0,0,0,157,0,75,0,95,0,133,0,8,0,103,0,129,0,239,0,0,0,0,0,0,0,0,0,76,0,83,0,0,0,246,0,249,0,124,0,5,0,0,0,141,0,136,0,98,0,76,0,193,0,62,0,221,0,69,0,187,0,63,0,0,0,15,0,204,0,136,0,24,0,0,0,214,0,3,0,120,0,159,0,238,0,139,0,171,0,39,0,154,0,186,0,228,0,38,0,214,0,13,0,51,0,78,0,64,0,251,0,217,0,182,0,124,0,17,0,121,0,236,0,22,0,63,0,40,0,0,0,201,0,231,0,58,0,0,0,99,0,163,0,23,0,249,0,27,0,0,0,216,0,254,0,21,0,135,0,143,0,139,0,0,0,31,0,23,0,0,0,134,0,63,0,53,0,118,0,90,0,11,0,238,0,76,0,191,0,109,0,0,0,254,0,205,0,181,0,97,0,0,0,32,0,181,0,0,0,18,0,193,0,128,0,34,0,0,0,23,0,82,0,19,0,144,0,64,0,250,0,0,0,181,0,0,0,139,0,185,0,39,0,105,0,0,0,78,0,0,0,119,0,151,0,82,0,157,0,11,0,200,0,0,0,1,0,29,0,167,0,235,0,70,0,105,0,0,0,219,0,19,0,179,0,120,0,230,0,246,0,2,0,0,0,96,0,82,0,252,0,0,0,0,0,228,0,245,0,250,0,177,0,3,0,85,0,81,0,160,0,165,0,213,0,27,0,191,0,86,0,102,0,0,0,198,0,0,0,111,0,0,0,86,0,0,0,47,0,131,0,173,0,229,0,198,0,71,0,27,0,141,0,76,0,205,0,197,0,145,0,122,0,227,0,161,0,208,0,14,0,143,0,229,0,12,0,0,0,164,0,193,0,228,0,87,0,227,0,101,0,113,0,74,0,236,0,48,0,0,0,191,0,51,0,0,0,75,0,0,0,189,0,138,0,182,0,179,0,195,0,127,0,0,0,15,0,0,0,20,0,0,0,185,0,0,0,242,0,0,0,207,0,229,0,134,0,82,0,151,0,0,0,80,0,250,0,0,0,81,0,181,0,146,0,224,0,21,0,19,0,239,0,0,0,190,0,54,0,14,0,133,0,135,0,0,0,69,0,0,0,0,0,30,0,72,0,113,0,31,0,133,0,33,0,168,0,0,0,175,0,83,0,0,0,51,0,46,0,95,0,132,0,223,0,200,0,156,0,150,0,0,0,211,0,252,0,234,0,198,0,246,0,89,0,32,0,92,0,220,0,255,0,133,0,174,0,82,0,170,0,29,0,43,0,183,0,0,0,0,0,222,0,67,0,113,0,254,0,187,0,254,0,221,0,0,0,168,0,0,0,0,0,38,0,162,0,232,0,97,0,208,0,24,0,83,0,11,0,67,0,159,0,0,0,117,0,198,0,119,0,215,0,206,0,0,0,179,0,0,0,0,0,66,0,103,0,187,0,9,0,157,0,217,0,0,0,189,0,32,0,0,0,1,0,127,0,93,0,165,0,161,0,231,0,0,0,0,0,13,0,0,0,30,0,188,0,80,0,37,0,202,0,243,0,0,0,0,0,7,0,138,0,47,0,73,0,241,0,8,0,209,0,242,0,185,0,149,0,142,0,151,0,24,0,140,0,196,0,213,0,243,0,131,0,142,0,149,0,20,0,28,0,221,0,190,0,0,0,222,0,8,0,198,0,0,0,109,0,250,0,209,0,61,0,80,0,176,0,84,0,160,0,165,0,36,0,4,0,71,0,253,0,27,0,0,0,225,0,85,0,192,0,104,0,0,0,3,0,63,0,45,0,65,0,31,0,7,0,178,0,199,0,238,0,23,0,0,0,0,0,87,0,42,0,37,0,138,0,0,0,109,0,60,0,173,0,158,0,180,0,111,0,226,0,0,0,104,0,246,0,130,0,129,0,0,0,0,0,124,0,158,0,155,0,25,0,164,0,119,0,115,0,0,0,165,0,162,0,52,0,96,0,164,0,0,0,0,0,244,0,0,0,20,0,200,0,76,0,42,0,0,0,159,0,75,0,0,0,117,0,121,0,16,0,172,0,0,0,29,0,61,0,92,0,100,0,76,0,43,0,218,0,82,0,18,0,14,0,0,0,16,0,135,0,208,0,108,0,227,0,0,0,119,0,201,0,62,0,25,0,143,0,198,0,58,0,0,0,0,0,207,0,32,0,87,0,203,0,53,0,147,0,204,0,83,0,0,0,160,0,145,0,216,0,22,0,39,0,54,0,19,0,16,0,29,0,225,0,136,0,210,0,99,0,19,0,227,0,226,0,0,0,0,0,0,0,29,0,184,0,0,0,0,0,201,0,192,0,177,0,0,0,18,0,41,0,0,0,0,0,208,0,11,0,0,0,148,0,103,0,93,0,93,0,0,0,44,0,105,0,75,0,79,0,82,0,193,0,137,0,225,0,144,0,101,0,21,0,221,0,70,0,0,0,109,0,0,0,0,0,184,0,228,0,217,0,112,0,81,0,62,0,212,0,130,0,254,0,59,0,235,0,80,0,143,0,29,0,47,0,172,0,200,0,0,0,196,0,182,0,90,0,12,0,165,0,11,0,0,0,171,0,51,0,142,0,0,0,106,0,169,0,25,0,156,0,0,0,102,0,2,0,0,0,0,0,237,0,40,0,252,0,122,0,70,0,20,0,0,0,42,0,133,0,0,0,105,0,195,0,114,0,124,0,41,0,174,0,178,0,90,0,65,0,210,0,22,0,153,0,67,0,38,0,227,0,189,0,122,0,0,0,209,0,19,0,39,0,119,0,138,0,42,0,73,0,242,0,23,0,65,0,49,0,181,0,125,0,0,0,136,0,66,0,0,0,77,0,4,0,28,0,112,0,129,0,72,0,0,0,0,0,77,0,32,0,236,0,46,0,0,0,21,0,141,0,41,0,0,0,147,0,98,0,169,0,0,0,19,0,157,0,34,0,47,0,229,0,0,0,133,0,124,0,0,0,43,0,141,0,247,0,97,0,196,0,40,0,81,0,39,0,166,0,42,0,135,0,196,0,16,0,116,0,164,0,127,0,133,0,145,0,142,0,0,0,22,0,0,0,180,0,29,0,14,0,149,0,212,0,234,0,190,0,0,0,0,0,42,0,0,0,129,0,111,0,247,0,4,0,0,0,0,0,20,0,233,0,240,0,98,0,51,0,81,0,89,0,0,0,178,0,227,0,178,0,248,0,0,0,56,0,7,0,241,0,129,0,77,0,5,0,0,0,68,0,103,0,55,0,171,0,214,0,110,0,96,0,3,0,169,0,0,0,165,0,56,0,80,0,146,0,114,0,150,0,250,0,170,0,123,0,0,0,244,0,80,0,47,0,120,0,60,0,33,0,100,0,66,0,49,0,53,0,91,0,184,0,210,0,191,0,32,0,247,0,76,0,0,0,22,0,88,0,124,0,119,0,0,0,30,0,136,0,86,0,92,0,158,0);
signal scenario_full  : scenario_type := (134,31,158,31,54,31,176,31,154,31,71,31,163,31,141,31,178,31,156,31,8,31,8,30,9,31,181,31,247,31,9,31,142,31,152,31,114,31,166,31,238,31,179,31,179,30,16,31,245,31,18,31,18,30,38,31,114,31,180,31,243,31,243,30,243,29,13,31,234,31,126,31,165,31,139,31,119,31,178,31,238,31,165,31,165,30,165,29,228,31,20,31,245,31,186,31,151,31,241,31,242,31,122,31,217,31,214,31,170,31,170,30,202,31,219,31,219,30,190,31,246,31,196,31,196,30,176,31,158,31,175,31,182,31,171,31,171,30,100,31,6,31,166,31,166,30,5,31,199,31,199,30,92,31,40,31,107,31,90,31,35,31,206,31,6,31,135,31,96,31,119,31,119,30,96,31,60,31,151,31,153,31,226,31,247,31,234,31,31,31,187,31,187,30,157,31,75,31,95,31,133,31,8,31,103,31,129,31,239,31,239,30,239,29,239,28,239,27,76,31,83,31,83,30,246,31,249,31,124,31,5,31,5,30,141,31,136,31,98,31,76,31,193,31,62,31,221,31,69,31,187,31,63,31,63,30,15,31,204,31,136,31,24,31,24,30,214,31,3,31,120,31,159,31,238,31,139,31,171,31,39,31,154,31,186,31,228,31,38,31,214,31,13,31,51,31,78,31,64,31,251,31,217,31,182,31,124,31,17,31,121,31,236,31,22,31,63,31,40,31,40,30,201,31,231,31,58,31,58,30,99,31,163,31,23,31,249,31,27,31,27,30,216,31,254,31,21,31,135,31,143,31,139,31,139,30,31,31,23,31,23,30,134,31,63,31,53,31,118,31,90,31,11,31,238,31,76,31,191,31,109,31,109,30,254,31,205,31,181,31,97,31,97,30,32,31,181,31,181,30,18,31,193,31,128,31,34,31,34,30,23,31,82,31,19,31,144,31,64,31,250,31,250,30,181,31,181,30,139,31,185,31,39,31,105,31,105,30,78,31,78,30,119,31,151,31,82,31,157,31,11,31,200,31,200,30,1,31,29,31,167,31,235,31,70,31,105,31,105,30,219,31,19,31,179,31,120,31,230,31,246,31,2,31,2,30,96,31,82,31,252,31,252,30,252,29,228,31,245,31,250,31,177,31,3,31,85,31,81,31,160,31,165,31,213,31,27,31,191,31,86,31,102,31,102,30,198,31,198,30,111,31,111,30,86,31,86,30,47,31,131,31,173,31,229,31,198,31,71,31,27,31,141,31,76,31,205,31,197,31,145,31,122,31,227,31,161,31,208,31,14,31,143,31,229,31,12,31,12,30,164,31,193,31,228,31,87,31,227,31,101,31,113,31,74,31,236,31,48,31,48,30,191,31,51,31,51,30,75,31,75,30,189,31,138,31,182,31,179,31,195,31,127,31,127,30,15,31,15,30,20,31,20,30,185,31,185,30,242,31,242,30,207,31,229,31,134,31,82,31,151,31,151,30,80,31,250,31,250,30,81,31,181,31,146,31,224,31,21,31,19,31,239,31,239,30,190,31,54,31,14,31,133,31,135,31,135,30,69,31,69,30,69,29,30,31,72,31,113,31,31,31,133,31,33,31,168,31,168,30,175,31,83,31,83,30,51,31,46,31,95,31,132,31,223,31,200,31,156,31,150,31,150,30,211,31,252,31,234,31,198,31,246,31,89,31,32,31,92,31,220,31,255,31,133,31,174,31,82,31,170,31,29,31,43,31,183,31,183,30,183,29,222,31,67,31,113,31,254,31,187,31,254,31,221,31,221,30,168,31,168,30,168,29,38,31,162,31,232,31,97,31,208,31,24,31,83,31,11,31,67,31,159,31,159,30,117,31,198,31,119,31,215,31,206,31,206,30,179,31,179,30,179,29,66,31,103,31,187,31,9,31,157,31,217,31,217,30,189,31,32,31,32,30,1,31,127,31,93,31,165,31,161,31,231,31,231,30,231,29,13,31,13,30,30,31,188,31,80,31,37,31,202,31,243,31,243,30,243,29,7,31,138,31,47,31,73,31,241,31,8,31,209,31,242,31,185,31,149,31,142,31,151,31,24,31,140,31,196,31,213,31,243,31,131,31,142,31,149,31,20,31,28,31,221,31,190,31,190,30,222,31,8,31,198,31,198,30,109,31,250,31,209,31,61,31,80,31,176,31,84,31,160,31,165,31,36,31,4,31,71,31,253,31,27,31,27,30,225,31,85,31,192,31,104,31,104,30,3,31,63,31,45,31,65,31,31,31,7,31,178,31,199,31,238,31,23,31,23,30,23,29,87,31,42,31,37,31,138,31,138,30,109,31,60,31,173,31,158,31,180,31,111,31,226,31,226,30,104,31,246,31,130,31,129,31,129,30,129,29,124,31,158,31,155,31,25,31,164,31,119,31,115,31,115,30,165,31,162,31,52,31,96,31,164,31,164,30,164,29,244,31,244,30,20,31,200,31,76,31,42,31,42,30,159,31,75,31,75,30,117,31,121,31,16,31,172,31,172,30,29,31,61,31,92,31,100,31,76,31,43,31,218,31,82,31,18,31,14,31,14,30,16,31,135,31,208,31,108,31,227,31,227,30,119,31,201,31,62,31,25,31,143,31,198,31,58,31,58,30,58,29,207,31,32,31,87,31,203,31,53,31,147,31,204,31,83,31,83,30,160,31,145,31,216,31,22,31,39,31,54,31,19,31,16,31,29,31,225,31,136,31,210,31,99,31,19,31,227,31,226,31,226,30,226,29,226,28,29,31,184,31,184,30,184,29,201,31,192,31,177,31,177,30,18,31,41,31,41,30,41,29,208,31,11,31,11,30,148,31,103,31,93,31,93,31,93,30,44,31,105,31,75,31,79,31,82,31,193,31,137,31,225,31,144,31,101,31,21,31,221,31,70,31,70,30,109,31,109,30,109,29,184,31,228,31,217,31,112,31,81,31,62,31,212,31,130,31,254,31,59,31,235,31,80,31,143,31,29,31,47,31,172,31,200,31,200,30,196,31,182,31,90,31,12,31,165,31,11,31,11,30,171,31,51,31,142,31,142,30,106,31,169,31,25,31,156,31,156,30,102,31,2,31,2,30,2,29,237,31,40,31,252,31,122,31,70,31,20,31,20,30,42,31,133,31,133,30,105,31,195,31,114,31,124,31,41,31,174,31,178,31,90,31,65,31,210,31,22,31,153,31,67,31,38,31,227,31,189,31,122,31,122,30,209,31,19,31,39,31,119,31,138,31,42,31,73,31,242,31,23,31,65,31,49,31,181,31,125,31,125,30,136,31,66,31,66,30,77,31,4,31,28,31,112,31,129,31,72,31,72,30,72,29,77,31,32,31,236,31,46,31,46,30,21,31,141,31,41,31,41,30,147,31,98,31,169,31,169,30,19,31,157,31,34,31,47,31,229,31,229,30,133,31,124,31,124,30,43,31,141,31,247,31,97,31,196,31,40,31,81,31,39,31,166,31,42,31,135,31,196,31,16,31,116,31,164,31,127,31,133,31,145,31,142,31,142,30,22,31,22,30,180,31,29,31,14,31,149,31,212,31,234,31,190,31,190,30,190,29,42,31,42,30,129,31,111,31,247,31,4,31,4,30,4,29,20,31,233,31,240,31,98,31,51,31,81,31,89,31,89,30,178,31,227,31,178,31,248,31,248,30,56,31,7,31,241,31,129,31,77,31,5,31,5,30,68,31,103,31,55,31,171,31,214,31,110,31,96,31,3,31,169,31,169,30,165,31,56,31,80,31,146,31,114,31,150,31,250,31,170,31,123,31,123,30,244,31,80,31,47,31,120,31,60,31,33,31,100,31,66,31,49,31,53,31,91,31,184,31,210,31,191,31,32,31,247,31,76,31,76,30,22,31,88,31,124,31,119,31,119,30,30,31,136,31,86,31,92,31,158,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
