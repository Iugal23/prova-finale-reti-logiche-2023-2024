-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_212 is
end project_tb_212;

architecture project_tb_arch_212 of project_tb_212 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 404;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (133,0,114,0,43,0,116,0,221,0,241,0,200,0,215,0,115,0,22,0,24,0,214,0,0,0,17,0,234,0,48,0,244,0,22,0,0,0,0,0,40,0,187,0,77,0,107,0,70,0,117,0,52,0,131,0,0,0,213,0,34,0,86,0,187,0,229,0,148,0,131,0,0,0,17,0,0,0,239,0,0,0,210,0,206,0,209,0,0,0,85,0,42,0,0,0,204,0,62,0,5,0,0,0,112,0,0,0,137,0,18,0,193,0,203,0,107,0,0,0,232,0,217,0,244,0,38,0,246,0,206,0,106,0,185,0,0,0,196,0,116,0,122,0,94,0,108,0,0,0,0,0,148,0,253,0,49,0,119,0,178,0,63,0,0,0,228,0,214,0,94,0,93,0,55,0,0,0,18,0,80,0,0,0,166,0,194,0,61,0,88,0,191,0,133,0,74,0,0,0,235,0,131,0,0,0,161,0,220,0,0,0,0,0,160,0,132,0,87,0,242,0,63,0,0,0,36,0,193,0,0,0,210,0,39,0,73,0,39,0,0,0,153,0,25,0,122,0,15,0,145,0,193,0,60,0,72,0,0,0,247,0,174,0,155,0,201,0,106,0,0,0,34,0,232,0,50,0,11,0,45,0,174,0,90,0,81,0,0,0,189,0,228,0,139,0,23,0,87,0,31,0,0,0,31,0,200,0,86,0,23,0,254,0,42,0,166,0,178,0,95,0,72,0,28,0,0,0,0,0,118,0,226,0,99,0,191,0,161,0,100,0,138,0,234,0,18,0,0,0,17,0,59,0,2,0,237,0,5,0,249,0,33,0,0,0,204,0,65,0,60,0,17,0,220,0,53,0,136,0,67,0,85,0,0,0,102,0,254,0,208,0,73,0,0,0,164,0,117,0,132,0,190,0,0,0,149,0,0,0,0,0,129,0,109,0,125,0,20,0,0,0,228,0,124,0,0,0,149,0,19,0,84,0,115,0,166,0,34,0,157,0,0,0,228,0,218,0,62,0,169,0,125,0,173,0,0,0,165,0,142,0,199,0,36,0,0,0,112,0,68,0,0,0,204,0,28,0,0,0,187,0,0,0,248,0,159,0,206,0,73,0,230,0,0,0,159,0,133,0,0,0,109,0,178,0,95,0,194,0,78,0,225,0,100,0,170,0,123,0,106,0,0,0,0,0,198,0,37,0,38,0,86,0,52,0,160,0,0,0,110,0,185,0,248,0,101,0,248,0,214,0,49,0,108,0,181,0,0,0,120,0,16,0,58,0,64,0,0,0,174,0,33,0,155,0,185,0,106,0,99,0,147,0,158,0,0,0,175,0,0,0,114,0,0,0,179,0,146,0,26,0,127,0,6,0,14,0,154,0,130,0,166,0,189,0,72,0,174,0,134,0,0,0,20,0,201,0,249,0,49,0,67,0,183,0,50,0,41,0,73,0,126,0,80,0,190,0,60,0,115,0,233,0,13,0,0,0,0,0,149,0,162,0,45,0,71,0,1,0,105,0,148,0,133,0,35,0,166,0,158,0,20,0,143,0,105,0,0,0,0,0,24,0,207,0,203,0,121,0,0,0,75,0,233,0,62,0,93,0,83,0,233,0,199,0,123,0,16,0,99,0,3,0,119,0,233,0,20,0,202,0,83,0,72,0,34,0,67,0,249,0,51,0,252,0,0,0,225,0,0,0,166,0,127,0,202,0,0,0,236,0,18,0,82,0,189,0,251,0,0,0,197,0,14,0,0,0,245,0,0,0,166,0,95,0,108,0,226,0,0,0,247,0,93,0,0,0,148,0,32,0,73,0,218,0,41,0);
signal scenario_full  : scenario_type := (133,31,114,31,43,31,116,31,221,31,241,31,200,31,215,31,115,31,22,31,24,31,214,31,214,30,17,31,234,31,48,31,244,31,22,31,22,30,22,29,40,31,187,31,77,31,107,31,70,31,117,31,52,31,131,31,131,30,213,31,34,31,86,31,187,31,229,31,148,31,131,31,131,30,17,31,17,30,239,31,239,30,210,31,206,31,209,31,209,30,85,31,42,31,42,30,204,31,62,31,5,31,5,30,112,31,112,30,137,31,18,31,193,31,203,31,107,31,107,30,232,31,217,31,244,31,38,31,246,31,206,31,106,31,185,31,185,30,196,31,116,31,122,31,94,31,108,31,108,30,108,29,148,31,253,31,49,31,119,31,178,31,63,31,63,30,228,31,214,31,94,31,93,31,55,31,55,30,18,31,80,31,80,30,166,31,194,31,61,31,88,31,191,31,133,31,74,31,74,30,235,31,131,31,131,30,161,31,220,31,220,30,220,29,160,31,132,31,87,31,242,31,63,31,63,30,36,31,193,31,193,30,210,31,39,31,73,31,39,31,39,30,153,31,25,31,122,31,15,31,145,31,193,31,60,31,72,31,72,30,247,31,174,31,155,31,201,31,106,31,106,30,34,31,232,31,50,31,11,31,45,31,174,31,90,31,81,31,81,30,189,31,228,31,139,31,23,31,87,31,31,31,31,30,31,31,200,31,86,31,23,31,254,31,42,31,166,31,178,31,95,31,72,31,28,31,28,30,28,29,118,31,226,31,99,31,191,31,161,31,100,31,138,31,234,31,18,31,18,30,17,31,59,31,2,31,237,31,5,31,249,31,33,31,33,30,204,31,65,31,60,31,17,31,220,31,53,31,136,31,67,31,85,31,85,30,102,31,254,31,208,31,73,31,73,30,164,31,117,31,132,31,190,31,190,30,149,31,149,30,149,29,129,31,109,31,125,31,20,31,20,30,228,31,124,31,124,30,149,31,19,31,84,31,115,31,166,31,34,31,157,31,157,30,228,31,218,31,62,31,169,31,125,31,173,31,173,30,165,31,142,31,199,31,36,31,36,30,112,31,68,31,68,30,204,31,28,31,28,30,187,31,187,30,248,31,159,31,206,31,73,31,230,31,230,30,159,31,133,31,133,30,109,31,178,31,95,31,194,31,78,31,225,31,100,31,170,31,123,31,106,31,106,30,106,29,198,31,37,31,38,31,86,31,52,31,160,31,160,30,110,31,185,31,248,31,101,31,248,31,214,31,49,31,108,31,181,31,181,30,120,31,16,31,58,31,64,31,64,30,174,31,33,31,155,31,185,31,106,31,99,31,147,31,158,31,158,30,175,31,175,30,114,31,114,30,179,31,146,31,26,31,127,31,6,31,14,31,154,31,130,31,166,31,189,31,72,31,174,31,134,31,134,30,20,31,201,31,249,31,49,31,67,31,183,31,50,31,41,31,73,31,126,31,80,31,190,31,60,31,115,31,233,31,13,31,13,30,13,29,149,31,162,31,45,31,71,31,1,31,105,31,148,31,133,31,35,31,166,31,158,31,20,31,143,31,105,31,105,30,105,29,24,31,207,31,203,31,121,31,121,30,75,31,233,31,62,31,93,31,83,31,233,31,199,31,123,31,16,31,99,31,3,31,119,31,233,31,20,31,202,31,83,31,72,31,34,31,67,31,249,31,51,31,252,31,252,30,225,31,225,30,166,31,127,31,202,31,202,30,236,31,18,31,82,31,189,31,251,31,251,30,197,31,14,31,14,30,245,31,245,30,166,31,95,31,108,31,226,31,226,30,247,31,93,31,93,30,148,31,32,31,73,31,218,31,41,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
