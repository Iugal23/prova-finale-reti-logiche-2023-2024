-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 375;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (149,0,216,0,113,0,250,0,198,0,176,0,41,0,0,0,232,0,180,0,173,0,206,0,28,0,0,0,127,0,163,0,128,0,166,0,93,0,146,0,225,0,206,0,195,0,200,0,112,0,227,0,0,0,61,0,94,0,177,0,37,0,76,0,172,0,36,0,55,0,3,0,0,0,80,0,160,0,0,0,141,0,63,0,174,0,97,0,137,0,190,0,200,0,149,0,150,0,217,0,41,0,72,0,146,0,149,0,74,0,251,0,0,0,221,0,96,0,0,0,140,0,30,0,58,0,239,0,59,0,146,0,0,0,204,0,106,0,186,0,48,0,13,0,82,0,0,0,128,0,190,0,144,0,205,0,77,0,209,0,69,0,65,0,136,0,0,0,222,0,224,0,0,0,0,0,86,0,0,0,115,0,4,0,0,0,147,0,38,0,70,0,49,0,153,0,12,0,39,0,0,0,0,0,199,0,128,0,12,0,201,0,243,0,224,0,91,0,219,0,2,0,163,0,158,0,28,0,66,0,161,0,0,0,247,0,85,0,147,0,90,0,0,0,222,0,161,0,203,0,215,0,49,0,140,0,190,0,22,0,125,0,240,0,134,0,175,0,190,0,122,0,0,0,0,0,95,0,111,0,37,0,81,0,215,0,30,0,0,0,247,0,20,0,34,0,199,0,156,0,9,0,0,0,140,0,41,0,126,0,253,0,28,0,243,0,175,0,156,0,27,0,0,0,0,0,0,0,0,0,71,0,198,0,95,0,182,0,0,0,237,0,139,0,168,0,145,0,26,0,0,0,114,0,20,0,21,0,174,0,185,0,87,0,248,0,5,0,0,0,9,0,21,0,237,0,0,0,0,0,6,0,0,0,199,0,0,0,0,0,0,0,14,0,66,0,201,0,50,0,2,0,152,0,0,0,0,0,200,0,107,0,220,0,68,0,232,0,235,0,0,0,0,0,181,0,220,0,0,0,0,0,56,0,99,0,78,0,119,0,78,0,0,0,247,0,226,0,0,0,84,0,0,0,77,0,192,0,149,0,26,0,238,0,164,0,0,0,12,0,178,0,236,0,0,0,79,0,241,0,61,0,178,0,0,0,0,0,181,0,26,0,0,0,0,0,44,0,87,0,160,0,159,0,0,0,201,0,79,0,5,0,153,0,132,0,122,0,0,0,255,0,15,0,172,0,74,0,0,0,76,0,85,0,91,0,147,0,0,0,41,0,180,0,130,0,126,0,55,0,170,0,0,0,0,0,222,0,175,0,183,0,69,0,147,0,95,0,14,0,0,0,7,0,70,0,112,0,236,0,49,0,222,0,48,0,196,0,242,0,219,0,190,0,175,0,237,0,82,0,35,0,49,0,0,0,117,0,17,0,61,0,166,0,30,0,0,0,0,0,107,0,108,0,97,0,171,0,0,0,147,0,194,0,0,0,111,0,105,0,25,0,44,0,202,0,250,0,0,0,5,0,0,0,0,0,0,0,149,0,141,0,0,0,133,0,129,0,20,0,189,0,81,0,0,0,32,0,178,0,140,0,173,0,130,0,75,0,14,0,202,0,167,0,222,0,33,0,0,0,143,0,156,0,213,0,0,0,0,0,0,0,45,0,144,0,0,0,133,0,51,0,255,0,0,0,0,0,10,0,238,0,4,0,73,0,47,0,81,0,247,0,0,0,134,0,55,0,214,0);
signal scenario_full  : scenario_type := (149,31,216,31,113,31,250,31,198,31,176,31,41,31,41,30,232,31,180,31,173,31,206,31,28,31,28,30,127,31,163,31,128,31,166,31,93,31,146,31,225,31,206,31,195,31,200,31,112,31,227,31,227,30,61,31,94,31,177,31,37,31,76,31,172,31,36,31,55,31,3,31,3,30,80,31,160,31,160,30,141,31,63,31,174,31,97,31,137,31,190,31,200,31,149,31,150,31,217,31,41,31,72,31,146,31,149,31,74,31,251,31,251,30,221,31,96,31,96,30,140,31,30,31,58,31,239,31,59,31,146,31,146,30,204,31,106,31,186,31,48,31,13,31,82,31,82,30,128,31,190,31,144,31,205,31,77,31,209,31,69,31,65,31,136,31,136,30,222,31,224,31,224,30,224,29,86,31,86,30,115,31,4,31,4,30,147,31,38,31,70,31,49,31,153,31,12,31,39,31,39,30,39,29,199,31,128,31,12,31,201,31,243,31,224,31,91,31,219,31,2,31,163,31,158,31,28,31,66,31,161,31,161,30,247,31,85,31,147,31,90,31,90,30,222,31,161,31,203,31,215,31,49,31,140,31,190,31,22,31,125,31,240,31,134,31,175,31,190,31,122,31,122,30,122,29,95,31,111,31,37,31,81,31,215,31,30,31,30,30,247,31,20,31,34,31,199,31,156,31,9,31,9,30,140,31,41,31,126,31,253,31,28,31,243,31,175,31,156,31,27,31,27,30,27,29,27,28,27,27,71,31,198,31,95,31,182,31,182,30,237,31,139,31,168,31,145,31,26,31,26,30,114,31,20,31,21,31,174,31,185,31,87,31,248,31,5,31,5,30,9,31,21,31,237,31,237,30,237,29,6,31,6,30,199,31,199,30,199,29,199,28,14,31,66,31,201,31,50,31,2,31,152,31,152,30,152,29,200,31,107,31,220,31,68,31,232,31,235,31,235,30,235,29,181,31,220,31,220,30,220,29,56,31,99,31,78,31,119,31,78,31,78,30,247,31,226,31,226,30,84,31,84,30,77,31,192,31,149,31,26,31,238,31,164,31,164,30,12,31,178,31,236,31,236,30,79,31,241,31,61,31,178,31,178,30,178,29,181,31,26,31,26,30,26,29,44,31,87,31,160,31,159,31,159,30,201,31,79,31,5,31,153,31,132,31,122,31,122,30,255,31,15,31,172,31,74,31,74,30,76,31,85,31,91,31,147,31,147,30,41,31,180,31,130,31,126,31,55,31,170,31,170,30,170,29,222,31,175,31,183,31,69,31,147,31,95,31,14,31,14,30,7,31,70,31,112,31,236,31,49,31,222,31,48,31,196,31,242,31,219,31,190,31,175,31,237,31,82,31,35,31,49,31,49,30,117,31,17,31,61,31,166,31,30,31,30,30,30,29,107,31,108,31,97,31,171,31,171,30,147,31,194,31,194,30,111,31,105,31,25,31,44,31,202,31,250,31,250,30,5,31,5,30,5,29,5,28,149,31,141,31,141,30,133,31,129,31,20,31,189,31,81,31,81,30,32,31,178,31,140,31,173,31,130,31,75,31,14,31,202,31,167,31,222,31,33,31,33,30,143,31,156,31,213,31,213,30,213,29,213,28,45,31,144,31,144,30,133,31,51,31,255,31,255,30,255,29,10,31,238,31,4,31,73,31,47,31,81,31,247,31,247,30,134,31,55,31,214,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
