-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 986;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,156,0,0,0,0,0,216,0,147,0,199,0,0,0,0,0,135,0,0,0,185,0,138,0,0,0,159,0,178,0,78,0,97,0,33,0,0,0,3,0,248,0,143,0,112,0,173,0,192,0,238,0,32,0,116,0,188,0,8,0,132,0,143,0,0,0,70,0,41,0,0,0,61,0,82,0,23,0,141,0,149,0,223,0,77,0,0,0,0,0,75,0,155,0,111,0,97,0,0,0,0,0,75,0,121,0,188,0,193,0,0,0,0,0,123,0,64,0,0,0,104,0,244,0,118,0,227,0,0,0,183,0,7,0,45,0,210,0,49,0,116,0,5,0,198,0,0,0,223,0,144,0,178,0,0,0,115,0,222,0,0,0,9,0,0,0,87,0,0,0,23,0,136,0,141,0,145,0,149,0,0,0,0,0,94,0,153,0,0,0,0,0,26,0,139,0,0,0,9,0,0,0,248,0,0,0,200,0,198,0,165,0,146,0,0,0,194,0,0,0,0,0,40,0,150,0,143,0,47,0,0,0,140,0,137,0,250,0,182,0,96,0,132,0,175,0,131,0,39,0,54,0,0,0,0,0,179,0,36,0,0,0,129,0,86,0,27,0,242,0,140,0,6,0,0,0,176,0,184,0,19,0,0,0,251,0,0,0,243,0,190,0,195,0,0,0,0,0,16,0,128,0,0,0,20,0,7,0,109,0,0,0,10,0,0,0,22,0,128,0,91,0,0,0,16,0,45,0,86,0,0,0,92,0,243,0,125,0,0,0,45,0,60,0,235,0,171,0,0,0,66,0,204,0,0,0,120,0,152,0,159,0,252,0,159,0,0,0,104,0,193,0,119,0,101,0,246,0,123,0,0,0,204,0,82,0,4,0,213,0,254,0,199,0,141,0,245,0,0,0,15,0,228,0,81,0,124,0,0,0,0,0,197,0,194,0,231,0,0,0,254,0,28,0,0,0,230,0,184,0,227,0,252,0,185,0,194,0,144,0,194,0,245,0,20,0,207,0,229,0,7,0,0,0,128,0,72,0,188,0,4,0,30,0,126,0,13,0,21,0,150,0,18,0,107,0,112,0,142,0,130,0,176,0,80,0,45,0,104,0,0,0,168,0,106,0,247,0,181,0,206,0,197,0,0,0,0,0,106,0,0,0,242,0,149,0,147,0,0,0,0,0,204,0,0,0,86,0,0,0,55,0,77,0,0,0,116,0,0,0,0,0,9,0,206,0,237,0,195,0,0,0,0,0,198,0,0,0,130,0,198,0,24,0,0,0,0,0,253,0,138,0,187,0,226,0,58,0,0,0,83,0,0,0,0,0,104,0,75,0,158,0,117,0,4,0,245,0,203,0,0,0,129,0,34,0,179,0,20,0,241,0,178,0,0,0,29,0,233,0,170,0,198,0,72,0,0,0,252,0,39,0,163,0,205,0,77,0,152,0,179,0,255,0,169,0,112,0,22,0,111,0,142,0,146,0,174,0,20,0,28,0,136,0,0,0,174,0,164,0,174,0,0,0,4,0,242,0,243,0,21,0,214,0,214,0,0,0,0,0,0,0,129,0,52,0,0,0,160,0,233,0,0,0,140,0,253,0,0,0,124,0,107,0,220,0,0,0,0,0,93,0,0,0,160,0,98,0,107,0,0,0,55,0,146,0,92,0,70,0,112,0,173,0,42,0,20,0,76,0,0,0,170,0,7,0,249,0,8,0,175,0,0,0,0,0,225,0,0,0,224,0,0,0,75,0,203,0,155,0,168,0,0,0,242,0,102,0,113,0,142,0,80,0,64,0,196,0,193,0,213,0,0,0,67,0,184,0,81,0,60,0,58,0,245,0,0,0,180,0,13,0,27,0,114,0,207,0,69,0,0,0,0,0,0,0,51,0,118,0,70,0,109,0,176,0,180,0,145,0,0,0,0,0,223,0,16,0,0,0,125,0,0,0,208,0,180,0,209,0,224,0,92,0,0,0,153,0,57,0,75,0,0,0,108,0,0,0,20,0,2,0,0,0,150,0,199,0,0,0,210,0,92,0,251,0,173,0,181,0,0,0,0,0,176,0,6,0,34,0,21,0,253,0,18,0,156,0,62,0,62,0,0,0,4,0,57,0,132,0,113,0,100,0,226,0,224,0,142,0,166,0,101,0,0,0,110,0,255,0,0,0,187,0,253,0,21,0,0,0,168,0,111,0,34,0,19,0,14,0,36,0,41,0,133,0,224,0,99,0,13,0,87,0,129,0,28,0,78,0,179,0,238,0,158,0,10,0,139,0,53,0,79,0,0,0,83,0,218,0,0,0,7,0,146,0,57,0,16,0,241,0,129,0,112,0,121,0,103,0,66,0,144,0,119,0,21,0,4,0,0,0,0,0,217,0,146,0,58,0,135,0,117,0,50,0,59,0,166,0,175,0,212,0,193,0,165,0,178,0,0,0,162,0,182,0,0,0,0,0,172,0,92,0,43,0,110,0,163,0,0,0,19,0,253,0,79,0,49,0,131,0,34,0,122,0,172,0,117,0,97,0,44,0,0,0,0,0,79,0,79,0,250,0,239,0,6,0,118,0,155,0,13,0,31,0,23,0,145,0,0,0,34,0,241,0,150,0,24,0,198,0,0,0,11,0,148,0,131,0,209,0,63,0,145,0,159,0,134,0,145,0,239,0,192,0,176,0,40,0,114,0,200,0,131,0,197,0,0,0,0,0,44,0,122,0,107,0,209,0,0,0,230,0,139,0,86,0,253,0,39,0,98,0,0,0,0,0,244,0,38,0,0,0,59,0,97,0,57,0,250,0,64,0,207,0,16,0,100,0,203,0,138,0,189,0,59,0,0,0,56,0,69,0,129,0,211,0,153,0,233,0,160,0,56,0,0,0,111,0,87,0,87,0,184,0,238,0,42,0,195,0,0,0,120,0,0,0,0,0,124,0,53,0,103,0,230,0,31,0,0,0,93,0,44,0,85,0,140,0,79,0,0,0,7,0,175,0,190,0,174,0,94,0,78,0,15,0,0,0,192,0,37,0,0,0,180,0,0,0,245,0,142,0,225,0,230,0,61,0,111,0,232,0,238,0,0,0,159,0,0,0,239,0,253,0,127,0,29,0,1,0,213,0,0,0,0,0,45,0,140,0,168,0,190,0,241,0,68,0,82,0,113,0,70,0,77,0,94,0,0,0,232,0,237,0,104,0,16,0,200,0,132,0,134,0,0,0,16,0,138,0,31,0,24,0,158,0,61,0,94,0,0,0,39,0,19,0,0,0,0,0,37,0,148,0,122,0,53,0,147,0,83,0,1,0,0,0,157,0,59,0,143,0,59,0,0,0,41,0,22,0,0,0,170,0,236,0,32,0,91,0,0,0,196,0,54,0,17,0,97,0,179,0,0,0,5,0,0,0,1,0,202,0,62,0,195,0,247,0,134,0,87,0,0,0,145,0,158,0,90,0,251,0,127,0,215,0,33,0,131,0,70,0,0,0,0,0,171,0,34,0,221,0,225,0,67,0,112,0,252,0,68,0,6,0,22,0,215,0,202,0,128,0,65,0,246,0,80,0,0,0,246,0,101,0,0,0,75,0,89,0,0,0,0,0,0,0,238,0,0,0,161,0,251,0,252,0,17,0,158,0,142,0,66,0,114,0,253,0,233,0,156,0,0,0,93,0,0,0,95,0,87,0,13,0,179,0,12,0,0,0,163,0,0,0,187,0,188,0,194,0,67,0,0,0,238,0,200,0,82,0,5,0,0,0,253,0,76,0,150,0,37,0,30,0,157,0,0,0,186,0,39,0,47,0,143,0,42,0,26,0,120,0,183,0,138,0,182,0,0,0,148,0,52,0,189,0,198,0,165,0,147,0,0,0,0,0,225,0,0,0,95,0,58,0,110,0,252,0,201,0,170,0,69,0,117,0,174,0,28,0,139,0,66,0,185,0,8,0,0,0,183,0,175,0,0,0,178,0,71,0,115,0,36,0,20,0,235,0,181,0,16,0,116,0,166,0,167,0,135,0,181,0,49,0,215,0,194,0,228,0,186,0,227,0,108,0,229,0,101,0,0,0,139,0,72,0,0,0,0,0,45,0,0,0,180,0,250,0,0,0,205,0,0,0,173,0,185,0,0,0,2,0,0,0,59,0,0,0,135,0,235,0,200,0,68,0,0,0,117,0,251,0,253,0,63,0,91,0,164,0,155,0,0,0,86,0,93,0,121,0,231,0,243,0,4,0,146,0,137,0,0,0,0,0,147,0,109,0,0,0,14,0,53,0,30,0,0,0,0,0,0,0,202,0,225,0,0,0,104,0,219,0,3,0,13,0,9,0,240,0,244,0,247,0,0,0,65,0,0,0,0,0,246,0,0,0,31,0,200,0,0,0,0,0,0,0,3,0,175,0,0,0,230,0,219,0,234,0,160,0,0,0,78,0,173,0,242,0);
signal scenario_full  : scenario_type := (0,0,156,31,156,30,156,29,216,31,147,31,199,31,199,30,199,29,135,31,135,30,185,31,138,31,138,30,159,31,178,31,78,31,97,31,33,31,33,30,3,31,248,31,143,31,112,31,173,31,192,31,238,31,32,31,116,31,188,31,8,31,132,31,143,31,143,30,70,31,41,31,41,30,61,31,82,31,23,31,141,31,149,31,223,31,77,31,77,30,77,29,75,31,155,31,111,31,97,31,97,30,97,29,75,31,121,31,188,31,193,31,193,30,193,29,123,31,64,31,64,30,104,31,244,31,118,31,227,31,227,30,183,31,7,31,45,31,210,31,49,31,116,31,5,31,198,31,198,30,223,31,144,31,178,31,178,30,115,31,222,31,222,30,9,31,9,30,87,31,87,30,23,31,136,31,141,31,145,31,149,31,149,30,149,29,94,31,153,31,153,30,153,29,26,31,139,31,139,30,9,31,9,30,248,31,248,30,200,31,198,31,165,31,146,31,146,30,194,31,194,30,194,29,40,31,150,31,143,31,47,31,47,30,140,31,137,31,250,31,182,31,96,31,132,31,175,31,131,31,39,31,54,31,54,30,54,29,179,31,36,31,36,30,129,31,86,31,27,31,242,31,140,31,6,31,6,30,176,31,184,31,19,31,19,30,251,31,251,30,243,31,190,31,195,31,195,30,195,29,16,31,128,31,128,30,20,31,7,31,109,31,109,30,10,31,10,30,22,31,128,31,91,31,91,30,16,31,45,31,86,31,86,30,92,31,243,31,125,31,125,30,45,31,60,31,235,31,171,31,171,30,66,31,204,31,204,30,120,31,152,31,159,31,252,31,159,31,159,30,104,31,193,31,119,31,101,31,246,31,123,31,123,30,204,31,82,31,4,31,213,31,254,31,199,31,141,31,245,31,245,30,15,31,228,31,81,31,124,31,124,30,124,29,197,31,194,31,231,31,231,30,254,31,28,31,28,30,230,31,184,31,227,31,252,31,185,31,194,31,144,31,194,31,245,31,20,31,207,31,229,31,7,31,7,30,128,31,72,31,188,31,4,31,30,31,126,31,13,31,21,31,150,31,18,31,107,31,112,31,142,31,130,31,176,31,80,31,45,31,104,31,104,30,168,31,106,31,247,31,181,31,206,31,197,31,197,30,197,29,106,31,106,30,242,31,149,31,147,31,147,30,147,29,204,31,204,30,86,31,86,30,55,31,77,31,77,30,116,31,116,30,116,29,9,31,206,31,237,31,195,31,195,30,195,29,198,31,198,30,130,31,198,31,24,31,24,30,24,29,253,31,138,31,187,31,226,31,58,31,58,30,83,31,83,30,83,29,104,31,75,31,158,31,117,31,4,31,245,31,203,31,203,30,129,31,34,31,179,31,20,31,241,31,178,31,178,30,29,31,233,31,170,31,198,31,72,31,72,30,252,31,39,31,163,31,205,31,77,31,152,31,179,31,255,31,169,31,112,31,22,31,111,31,142,31,146,31,174,31,20,31,28,31,136,31,136,30,174,31,164,31,174,31,174,30,4,31,242,31,243,31,21,31,214,31,214,31,214,30,214,29,214,28,129,31,52,31,52,30,160,31,233,31,233,30,140,31,253,31,253,30,124,31,107,31,220,31,220,30,220,29,93,31,93,30,160,31,98,31,107,31,107,30,55,31,146,31,92,31,70,31,112,31,173,31,42,31,20,31,76,31,76,30,170,31,7,31,249,31,8,31,175,31,175,30,175,29,225,31,225,30,224,31,224,30,75,31,203,31,155,31,168,31,168,30,242,31,102,31,113,31,142,31,80,31,64,31,196,31,193,31,213,31,213,30,67,31,184,31,81,31,60,31,58,31,245,31,245,30,180,31,13,31,27,31,114,31,207,31,69,31,69,30,69,29,69,28,51,31,118,31,70,31,109,31,176,31,180,31,145,31,145,30,145,29,223,31,16,31,16,30,125,31,125,30,208,31,180,31,209,31,224,31,92,31,92,30,153,31,57,31,75,31,75,30,108,31,108,30,20,31,2,31,2,30,150,31,199,31,199,30,210,31,92,31,251,31,173,31,181,31,181,30,181,29,176,31,6,31,34,31,21,31,253,31,18,31,156,31,62,31,62,31,62,30,4,31,57,31,132,31,113,31,100,31,226,31,224,31,142,31,166,31,101,31,101,30,110,31,255,31,255,30,187,31,253,31,21,31,21,30,168,31,111,31,34,31,19,31,14,31,36,31,41,31,133,31,224,31,99,31,13,31,87,31,129,31,28,31,78,31,179,31,238,31,158,31,10,31,139,31,53,31,79,31,79,30,83,31,218,31,218,30,7,31,146,31,57,31,16,31,241,31,129,31,112,31,121,31,103,31,66,31,144,31,119,31,21,31,4,31,4,30,4,29,217,31,146,31,58,31,135,31,117,31,50,31,59,31,166,31,175,31,212,31,193,31,165,31,178,31,178,30,162,31,182,31,182,30,182,29,172,31,92,31,43,31,110,31,163,31,163,30,19,31,253,31,79,31,49,31,131,31,34,31,122,31,172,31,117,31,97,31,44,31,44,30,44,29,79,31,79,31,250,31,239,31,6,31,118,31,155,31,13,31,31,31,23,31,145,31,145,30,34,31,241,31,150,31,24,31,198,31,198,30,11,31,148,31,131,31,209,31,63,31,145,31,159,31,134,31,145,31,239,31,192,31,176,31,40,31,114,31,200,31,131,31,197,31,197,30,197,29,44,31,122,31,107,31,209,31,209,30,230,31,139,31,86,31,253,31,39,31,98,31,98,30,98,29,244,31,38,31,38,30,59,31,97,31,57,31,250,31,64,31,207,31,16,31,100,31,203,31,138,31,189,31,59,31,59,30,56,31,69,31,129,31,211,31,153,31,233,31,160,31,56,31,56,30,111,31,87,31,87,31,184,31,238,31,42,31,195,31,195,30,120,31,120,30,120,29,124,31,53,31,103,31,230,31,31,31,31,30,93,31,44,31,85,31,140,31,79,31,79,30,7,31,175,31,190,31,174,31,94,31,78,31,15,31,15,30,192,31,37,31,37,30,180,31,180,30,245,31,142,31,225,31,230,31,61,31,111,31,232,31,238,31,238,30,159,31,159,30,239,31,253,31,127,31,29,31,1,31,213,31,213,30,213,29,45,31,140,31,168,31,190,31,241,31,68,31,82,31,113,31,70,31,77,31,94,31,94,30,232,31,237,31,104,31,16,31,200,31,132,31,134,31,134,30,16,31,138,31,31,31,24,31,158,31,61,31,94,31,94,30,39,31,19,31,19,30,19,29,37,31,148,31,122,31,53,31,147,31,83,31,1,31,1,30,157,31,59,31,143,31,59,31,59,30,41,31,22,31,22,30,170,31,236,31,32,31,91,31,91,30,196,31,54,31,17,31,97,31,179,31,179,30,5,31,5,30,1,31,202,31,62,31,195,31,247,31,134,31,87,31,87,30,145,31,158,31,90,31,251,31,127,31,215,31,33,31,131,31,70,31,70,30,70,29,171,31,34,31,221,31,225,31,67,31,112,31,252,31,68,31,6,31,22,31,215,31,202,31,128,31,65,31,246,31,80,31,80,30,246,31,101,31,101,30,75,31,89,31,89,30,89,29,89,28,238,31,238,30,161,31,251,31,252,31,17,31,158,31,142,31,66,31,114,31,253,31,233,31,156,31,156,30,93,31,93,30,95,31,87,31,13,31,179,31,12,31,12,30,163,31,163,30,187,31,188,31,194,31,67,31,67,30,238,31,200,31,82,31,5,31,5,30,253,31,76,31,150,31,37,31,30,31,157,31,157,30,186,31,39,31,47,31,143,31,42,31,26,31,120,31,183,31,138,31,182,31,182,30,148,31,52,31,189,31,198,31,165,31,147,31,147,30,147,29,225,31,225,30,95,31,58,31,110,31,252,31,201,31,170,31,69,31,117,31,174,31,28,31,139,31,66,31,185,31,8,31,8,30,183,31,175,31,175,30,178,31,71,31,115,31,36,31,20,31,235,31,181,31,16,31,116,31,166,31,167,31,135,31,181,31,49,31,215,31,194,31,228,31,186,31,227,31,108,31,229,31,101,31,101,30,139,31,72,31,72,30,72,29,45,31,45,30,180,31,250,31,250,30,205,31,205,30,173,31,185,31,185,30,2,31,2,30,59,31,59,30,135,31,235,31,200,31,68,31,68,30,117,31,251,31,253,31,63,31,91,31,164,31,155,31,155,30,86,31,93,31,121,31,231,31,243,31,4,31,146,31,137,31,137,30,137,29,147,31,109,31,109,30,14,31,53,31,30,31,30,30,30,29,30,28,202,31,225,31,225,30,104,31,219,31,3,31,13,31,9,31,240,31,244,31,247,31,247,30,65,31,65,30,65,29,246,31,246,30,31,31,200,31,200,30,200,29,200,28,3,31,175,31,175,30,230,31,219,31,234,31,160,31,160,30,78,31,173,31,242,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
