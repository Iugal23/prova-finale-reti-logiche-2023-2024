-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 899;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,197,0,232,0,0,0,36,0,0,0,0,0,158,0,27,0,242,0,0,0,188,0,185,0,52,0,144,0,192,0,9,0,170,0,96,0,173,0,194,0,11,0,119,0,0,0,0,0,0,0,20,0,49,0,67,0,71,0,73,0,91,0,123,0,189,0,77,0,0,0,159,0,51,0,0,0,60,0,44,0,142,0,230,0,123,0,125,0,195,0,71,0,253,0,0,0,0,0,145,0,243,0,150,0,30,0,0,0,13,0,38,0,0,0,0,0,135,0,228,0,117,0,43,0,0,0,18,0,0,0,77,0,0,0,201,0,0,0,0,0,87,0,0,0,0,0,154,0,159,0,56,0,0,0,220,0,16,0,116,0,37,0,148,0,88,0,248,0,131,0,0,0,86,0,246,0,38,0,76,0,102,0,43,0,173,0,78,0,141,0,101,0,0,0,0,0,106,0,8,0,16,0,154,0,0,0,1,0,0,0,95,0,0,0,112,0,17,0,41,0,0,0,135,0,56,0,246,0,204,0,237,0,0,0,90,0,245,0,171,0,0,0,134,0,150,0,0,0,118,0,143,0,188,0,217,0,234,0,120,0,46,0,174,0,83,0,0,0,0,0,95,0,0,0,0,0,54,0,0,0,0,0,0,0,222,0,115,0,9,0,239,0,0,0,250,0,19,0,23,0,154,0,87,0,10,0,0,0,225,0,0,0,0,0,79,0,128,0,230,0,135,0,139,0,180,0,146,0,83,0,103,0,151,0,135,0,27,0,212,0,2,0,7,0,242,0,53,0,65,0,76,0,134,0,247,0,138,0,205,0,85,0,144,0,0,0,228,0,51,0,133,0,222,0,126,0,161,0,223,0,0,0,153,0,139,0,0,0,0,0,157,0,38,0,14,0,108,0,255,0,89,0,0,0,234,0,116,0,88,0,174,0,0,0,50,0,20,0,101,0,175,0,196,0,87,0,73,0,186,0,0,0,0,0,197,0,18,0,0,0,0,0,104,0,185,0,85,0,23,0,37,0,31,0,254,0,241,0,114,0,130,0,149,0,208,0,98,0,60,0,0,0,128,0,250,0,82,0,177,0,197,0,0,0,129,0,65,0,0,0,77,0,88,0,0,0,10,0,147,0,0,0,127,0,49,0,0,0,254,0,209,0,8,0,18,0,145,0,208,0,116,0,171,0,0,0,100,0,106,0,119,0,101,0,204,0,170,0,206,0,96,0,178,0,0,0,88,0,0,0,117,0,173,0,217,0,0,0,17,0,162,0,0,0,76,0,0,0,6,0,0,0,0,0,0,0,96,0,95,0,231,0,203,0,18,0,0,0,111,0,221,0,211,0,175,0,0,0,151,0,0,0,62,0,190,0,28,0,123,0,102,0,0,0,186,0,42,0,43,0,55,0,156,0,0,0,62,0,218,0,102,0,102,0,0,0,0,0,150,0,222,0,49,0,74,0,218,0,152,0,184,0,237,0,0,0,109,0,253,0,197,0,235,0,225,0,0,0,5,0,162,0,0,0,181,0,85,0,14,0,0,0,0,0,0,0,59,0,201,0,62,0,165,0,8,0,160,0,37,0,0,0,54,0,165,0,53,0,149,0,87,0,91,0,162,0,192,0,173,0,35,0,128,0,124,0,0,0,138,0,215,0,0,0,171,0,199,0,63,0,30,0,72,0,4,0,191,0,0,0,210,0,190,0,208,0,0,0,227,0,111,0,179,0,113,0,235,0,37,0,164,0,212,0,169,0,180,0,0,0,44,0,23,0,98,0,36,0,79,0,205,0,144,0,170,0,243,0,147,0,141,0,96,0,17,0,155,0,7,0,117,0,185,0,236,0,145,0,37,0,252,0,0,0,93,0,0,0,0,0,155,0,228,0,174,0,239,0,0,0,89,0,201,0,0,0,0,0,0,0,0,0,44,0,250,0,0,0,134,0,0,0,0,0,0,0,0,0,156,0,44,0,0,0,62,0,156,0,214,0,7,0,140,0,236,0,0,0,0,0,47,0,209,0,181,0,172,0,43,0,101,0,230,0,0,0,15,0,85,0,239,0,219,0,0,0,183,0,93,0,75,0,186,0,250,0,0,0,137,0,109,0,163,0,81,0,141,0,0,0,99,0,0,0,211,0,0,0,194,0,238,0,221,0,68,0,0,0,225,0,182,0,217,0,68,0,0,0,0,0,141,0,119,0,46,0,111,0,10,0,93,0,0,0,186,0,237,0,141,0,204,0,7,0,160,0,151,0,0,0,0,0,0,0,78,0,192,0,154,0,251,0,181,0,66,0,232,0,177,0,0,0,148,0,244,0,73,0,100,0,57,0,143,0,194,0,0,0,68,0,133,0,2,0,0,0,225,0,83,0,102,0,53,0,98,0,99,0,228,0,8,0,0,0,0,0,0,0,128,0,0,0,104,0,0,0,0,0,47,0,0,0,121,0,10,0,208,0,94,0,10,0,210,0,0,0,145,0,140,0,18,0,0,0,0,0,0,0,0,0,187,0,0,0,100,0,229,0,239,0,8,0,116,0,248,0,0,0,69,0,42,0,89,0,186,0,5,0,0,0,77,0,245,0,238,0,0,0,16,0,216,0,0,0,235,0,235,0,0,0,75,0,0,0,151,0,0,0,69,0,167,0,89,0,186,0,0,0,186,0,94,0,208,0,217,0,49,0,180,0,24,0,0,0,0,0,51,0,63,0,194,0,177,0,71,0,25,0,9,0,0,0,0,0,65,0,239,0,0,0,247,0,83,0,44,0,0,0,206,0,0,0,241,0,194,0,248,0,113,0,247,0,0,0,57,0,127,0,119,0,0,0,218,0,154,0,160,0,211,0,60,0,93,0,23,0,0,0,48,0,0,0,0,0,69,0,0,0,116,0,198,0,0,0,220,0,136,0,232,0,0,0,75,0,127,0,91,0,0,0,123,0,253,0,206,0,237,0,50,0,151,0,125,0,0,0,138,0,103,0,5,0,86,0,71,0,0,0,25,0,0,0,228,0,110,0,17,0,14,0,252,0,0,0,211,0,28,0,0,0,61,0,130,0,31,0,9,0,0,0,171,0,52,0,0,0,132,0,199,0,60,0,0,0,116,0,129,0,22,0,204,0,248,0,61,0,226,0,252,0,53,0,0,0,0,0,129,0,252,0,188,0,0,0,138,0,159,0,188,0,0,0,21,0,143,0,239,0,205,0,30,0,251,0,0,0,85,0,176,0,8,0,0,0,109,0,217,0,110,0,130,0,47,0,38,0,6,0,0,0,52,0,35,0,74,0,0,0,0,0,220,0,148,0,76,0,0,0,0,0,35,0,0,0,103,0,57,0,197,0,0,0,238,0,171,0,0,0,58,0,105,0,223,0,9,0,0,0,0,0,82,0,90,0,189,0,0,0,206,0,57,0,0,0,39,0,68,0,237,0,0,0,221,0,250,0,102,0,38,0,43,0,164,0,179,0,0,0,140,0,254,0,153,0,190,0,137,0,71,0,16,0,152,0,105,0,181,0,136,0,174,0,0,0,130,0,93,0,0,0,195,0,210,0,0,0,35,0,86,0,74,0,64,0,0,0,0,0,164,0,223,0,96,0,0,0,87,0,14,0,40,0,138,0,234,0,55,0,139,0,243,0,105,0,131,0,78,0,206,0,120,0,0,0,190,0,183,0,0,0,238,0,186,0,0,0,95,0,246,0,84,0,113,0,0,0,80,0,69,0,0,0,133,0,0,0,118,0,167,0,129,0,253,0,168,0,0,0,63,0,143,0,72,0,186,0,162,0,67,0,231,0,253,0,176,0,0,0,0,0,174,0,36,0,187,0,78,0,200,0,55,0,165,0,110,0,0,0,0,0,164,0,53,0,14,0,254,0,176,0,230,0,31,0,0,0,0,0,193,0,0,0,30,0,83,0,235,0,0,0,248,0,41,0,253,0,253,0,251,0,173,0,0,0,138,0,0,0,151,0,220,0,59,0,76,0,7,0,107,0,92,0,29,0,232,0,88,0,181,0,41,0,177,0,0,0,169,0,222,0,45,0,136,0,44,0);
signal scenario_full  : scenario_type := (0,0,197,31,232,31,232,30,36,31,36,30,36,29,158,31,27,31,242,31,242,30,188,31,185,31,52,31,144,31,192,31,9,31,170,31,96,31,173,31,194,31,11,31,119,31,119,30,119,29,119,28,20,31,49,31,67,31,71,31,73,31,91,31,123,31,189,31,77,31,77,30,159,31,51,31,51,30,60,31,44,31,142,31,230,31,123,31,125,31,195,31,71,31,253,31,253,30,253,29,145,31,243,31,150,31,30,31,30,30,13,31,38,31,38,30,38,29,135,31,228,31,117,31,43,31,43,30,18,31,18,30,77,31,77,30,201,31,201,30,201,29,87,31,87,30,87,29,154,31,159,31,56,31,56,30,220,31,16,31,116,31,37,31,148,31,88,31,248,31,131,31,131,30,86,31,246,31,38,31,76,31,102,31,43,31,173,31,78,31,141,31,101,31,101,30,101,29,106,31,8,31,16,31,154,31,154,30,1,31,1,30,95,31,95,30,112,31,17,31,41,31,41,30,135,31,56,31,246,31,204,31,237,31,237,30,90,31,245,31,171,31,171,30,134,31,150,31,150,30,118,31,143,31,188,31,217,31,234,31,120,31,46,31,174,31,83,31,83,30,83,29,95,31,95,30,95,29,54,31,54,30,54,29,54,28,222,31,115,31,9,31,239,31,239,30,250,31,19,31,23,31,154,31,87,31,10,31,10,30,225,31,225,30,225,29,79,31,128,31,230,31,135,31,139,31,180,31,146,31,83,31,103,31,151,31,135,31,27,31,212,31,2,31,7,31,242,31,53,31,65,31,76,31,134,31,247,31,138,31,205,31,85,31,144,31,144,30,228,31,51,31,133,31,222,31,126,31,161,31,223,31,223,30,153,31,139,31,139,30,139,29,157,31,38,31,14,31,108,31,255,31,89,31,89,30,234,31,116,31,88,31,174,31,174,30,50,31,20,31,101,31,175,31,196,31,87,31,73,31,186,31,186,30,186,29,197,31,18,31,18,30,18,29,104,31,185,31,85,31,23,31,37,31,31,31,254,31,241,31,114,31,130,31,149,31,208,31,98,31,60,31,60,30,128,31,250,31,82,31,177,31,197,31,197,30,129,31,65,31,65,30,77,31,88,31,88,30,10,31,147,31,147,30,127,31,49,31,49,30,254,31,209,31,8,31,18,31,145,31,208,31,116,31,171,31,171,30,100,31,106,31,119,31,101,31,204,31,170,31,206,31,96,31,178,31,178,30,88,31,88,30,117,31,173,31,217,31,217,30,17,31,162,31,162,30,76,31,76,30,6,31,6,30,6,29,6,28,96,31,95,31,231,31,203,31,18,31,18,30,111,31,221,31,211,31,175,31,175,30,151,31,151,30,62,31,190,31,28,31,123,31,102,31,102,30,186,31,42,31,43,31,55,31,156,31,156,30,62,31,218,31,102,31,102,31,102,30,102,29,150,31,222,31,49,31,74,31,218,31,152,31,184,31,237,31,237,30,109,31,253,31,197,31,235,31,225,31,225,30,5,31,162,31,162,30,181,31,85,31,14,31,14,30,14,29,14,28,59,31,201,31,62,31,165,31,8,31,160,31,37,31,37,30,54,31,165,31,53,31,149,31,87,31,91,31,162,31,192,31,173,31,35,31,128,31,124,31,124,30,138,31,215,31,215,30,171,31,199,31,63,31,30,31,72,31,4,31,191,31,191,30,210,31,190,31,208,31,208,30,227,31,111,31,179,31,113,31,235,31,37,31,164,31,212,31,169,31,180,31,180,30,44,31,23,31,98,31,36,31,79,31,205,31,144,31,170,31,243,31,147,31,141,31,96,31,17,31,155,31,7,31,117,31,185,31,236,31,145,31,37,31,252,31,252,30,93,31,93,30,93,29,155,31,228,31,174,31,239,31,239,30,89,31,201,31,201,30,201,29,201,28,201,27,44,31,250,31,250,30,134,31,134,30,134,29,134,28,134,27,156,31,44,31,44,30,62,31,156,31,214,31,7,31,140,31,236,31,236,30,236,29,47,31,209,31,181,31,172,31,43,31,101,31,230,31,230,30,15,31,85,31,239,31,219,31,219,30,183,31,93,31,75,31,186,31,250,31,250,30,137,31,109,31,163,31,81,31,141,31,141,30,99,31,99,30,211,31,211,30,194,31,238,31,221,31,68,31,68,30,225,31,182,31,217,31,68,31,68,30,68,29,141,31,119,31,46,31,111,31,10,31,93,31,93,30,186,31,237,31,141,31,204,31,7,31,160,31,151,31,151,30,151,29,151,28,78,31,192,31,154,31,251,31,181,31,66,31,232,31,177,31,177,30,148,31,244,31,73,31,100,31,57,31,143,31,194,31,194,30,68,31,133,31,2,31,2,30,225,31,83,31,102,31,53,31,98,31,99,31,228,31,8,31,8,30,8,29,8,28,128,31,128,30,104,31,104,30,104,29,47,31,47,30,121,31,10,31,208,31,94,31,10,31,210,31,210,30,145,31,140,31,18,31,18,30,18,29,18,28,18,27,187,31,187,30,100,31,229,31,239,31,8,31,116,31,248,31,248,30,69,31,42,31,89,31,186,31,5,31,5,30,77,31,245,31,238,31,238,30,16,31,216,31,216,30,235,31,235,31,235,30,75,31,75,30,151,31,151,30,69,31,167,31,89,31,186,31,186,30,186,31,94,31,208,31,217,31,49,31,180,31,24,31,24,30,24,29,51,31,63,31,194,31,177,31,71,31,25,31,9,31,9,30,9,29,65,31,239,31,239,30,247,31,83,31,44,31,44,30,206,31,206,30,241,31,194,31,248,31,113,31,247,31,247,30,57,31,127,31,119,31,119,30,218,31,154,31,160,31,211,31,60,31,93,31,23,31,23,30,48,31,48,30,48,29,69,31,69,30,116,31,198,31,198,30,220,31,136,31,232,31,232,30,75,31,127,31,91,31,91,30,123,31,253,31,206,31,237,31,50,31,151,31,125,31,125,30,138,31,103,31,5,31,86,31,71,31,71,30,25,31,25,30,228,31,110,31,17,31,14,31,252,31,252,30,211,31,28,31,28,30,61,31,130,31,31,31,9,31,9,30,171,31,52,31,52,30,132,31,199,31,60,31,60,30,116,31,129,31,22,31,204,31,248,31,61,31,226,31,252,31,53,31,53,30,53,29,129,31,252,31,188,31,188,30,138,31,159,31,188,31,188,30,21,31,143,31,239,31,205,31,30,31,251,31,251,30,85,31,176,31,8,31,8,30,109,31,217,31,110,31,130,31,47,31,38,31,6,31,6,30,52,31,35,31,74,31,74,30,74,29,220,31,148,31,76,31,76,30,76,29,35,31,35,30,103,31,57,31,197,31,197,30,238,31,171,31,171,30,58,31,105,31,223,31,9,31,9,30,9,29,82,31,90,31,189,31,189,30,206,31,57,31,57,30,39,31,68,31,237,31,237,30,221,31,250,31,102,31,38,31,43,31,164,31,179,31,179,30,140,31,254,31,153,31,190,31,137,31,71,31,16,31,152,31,105,31,181,31,136,31,174,31,174,30,130,31,93,31,93,30,195,31,210,31,210,30,35,31,86,31,74,31,64,31,64,30,64,29,164,31,223,31,96,31,96,30,87,31,14,31,40,31,138,31,234,31,55,31,139,31,243,31,105,31,131,31,78,31,206,31,120,31,120,30,190,31,183,31,183,30,238,31,186,31,186,30,95,31,246,31,84,31,113,31,113,30,80,31,69,31,69,30,133,31,133,30,118,31,167,31,129,31,253,31,168,31,168,30,63,31,143,31,72,31,186,31,162,31,67,31,231,31,253,31,176,31,176,30,176,29,174,31,36,31,187,31,78,31,200,31,55,31,165,31,110,31,110,30,110,29,164,31,53,31,14,31,254,31,176,31,230,31,31,31,31,30,31,29,193,31,193,30,30,31,83,31,235,31,235,30,248,31,41,31,253,31,253,31,251,31,173,31,173,30,138,31,138,30,151,31,220,31,59,31,76,31,7,31,107,31,92,31,29,31,232,31,88,31,181,31,41,31,177,31,177,30,169,31,222,31,45,31,136,31,44,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
