-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_581 is
end project_tb_581;

architecture project_tb_arch_581 of project_tb_581 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 717;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,7,0,128,0,102,0,83,0,0,0,230,0,4,0,69,0,88,0,95,0,138,0,161,0,111,0,0,0,0,0,45,0,148,0,230,0,8,0,159,0,214,0,163,0,75,0,62,0,0,0,25,0,168,0,0,0,28,0,139,0,0,0,37,0,183,0,77,0,78,0,0,0,0,0,173,0,71,0,0,0,20,0,0,0,27,0,130,0,18,0,36,0,0,0,227,0,93,0,147,0,0,0,33,0,39,0,184,0,0,0,0,0,85,0,85,0,0,0,0,0,185,0,255,0,0,0,119,0,0,0,41,0,182,0,231,0,120,0,242,0,0,0,242,0,41,0,111,0,0,0,91,0,0,0,233,0,0,0,0,0,209,0,0,0,33,0,158,0,51,0,182,0,171,0,119,0,90,0,203,0,55,0,194,0,122,0,207,0,170,0,206,0,186,0,207,0,8,0,43,0,70,0,0,0,79,0,31,0,144,0,4,0,51,0,138,0,107,0,21,0,15,0,72,0,149,0,130,0,151,0,232,0,76,0,195,0,194,0,158,0,109,0,238,0,0,0,0,0,0,0,183,0,205,0,58,0,131,0,141,0,4,0,0,0,198,0,126,0,26,0,175,0,149,0,243,0,205,0,202,0,220,0,228,0,118,0,102,0,0,0,228,0,200,0,116,0,241,0,118,0,174,0,0,0,0,0,49,0,238,0,249,0,19,0,176,0,0,0,21,0,246,0,59,0,0,0,175,0,87,0,215,0,4,0,0,0,124,0,0,0,166,0,233,0,12,0,87,0,245,0,88,0,56,0,124,0,85,0,76,0,170,0,76,0,157,0,0,0,120,0,11,0,0,0,0,0,14,0,130,0,0,0,0,0,202,0,0,0,194,0,206,0,0,0,126,0,186,0,203,0,150,0,124,0,167,0,89,0,163,0,0,0,0,0,0,0,88,0,52,0,139,0,186,0,252,0,37,0,27,0,0,0,68,0,0,0,0,0,0,0,100,0,82,0,103,0,0,0,118,0,159,0,223,0,196,0,168,0,48,0,48,0,4,0,144,0,139,0,143,0,0,0,22,0,147,0,221,0,150,0,10,0,103,0,61,0,92,0,236,0,44,0,110,0,3,0,0,0,120,0,20,0,199,0,0,0,0,0,0,0,181,0,61,0,254,0,85,0,37,0,180,0,185,0,0,0,0,0,114,0,124,0,0,0,49,0,212,0,0,0,248,0,0,0,149,0,235,0,0,0,38,0,222,0,227,0,214,0,4,0,64,0,87,0,6,0,85,0,59,0,138,0,230,0,241,0,144,0,20,0,197,0,206,0,0,0,128,0,195,0,7,0,73,0,0,0,50,0,0,0,227,0,163,0,33,0,161,0,0,0,156,0,74,0,74,0,160,0,98,0,202,0,214,0,222,0,209,0,193,0,71,0,40,0,94,0,38,0,221,0,97,0,201,0,44,0,222,0,36,0,167,0,0,0,157,0,82,0,231,0,198,0,0,0,172,0,0,0,149,0,235,0,99,0,16,0,60,0,184,0,139,0,99,0,230,0,135,0,146,0,212,0,93,0,0,0,232,0,211,0,14,0,0,0,158,0,230,0,221,0,40,0,0,0,158,0,33,0,0,0,66,0,214,0,6,0,110,0,63,0,15,0,232,0,78,0,133,0,65,0,0,0,223,0,62,0,114,0,23,0,0,0,93,0,74,0,173,0,0,0,81,0,223,0,207,0,191,0,154,0,131,0,148,0,156,0,0,0,251,0,254,0,158,0,243,0,137,0,112,0,54,0,7,0,191,0,0,0,15,0,63,0,100,0,208,0,67,0,233,0,0,0,242,0,141,0,0,0,166,0,106,0,0,0,41,0,98,0,26,0,142,0,0,0,216,0,239,0,118,0,11,0,38,0,46,0,0,0,201,0,0,0,61,0,202,0,41,0,0,0,0,0,221,0,95,0,0,0,229,0,222,0,0,0,48,0,44,0,178,0,107,0,98,0,0,0,0,0,4,0,25,0,0,0,84,0,46,0,233,0,76,0,231,0,150,0,65,0,253,0,213,0,186,0,177,0,106,0,160,0,0,0,247,0,0,0,86,0,248,0,111,0,178,0,51,0,152,0,122,0,0,0,112,0,152,0,22,0,227,0,131,0,192,0,0,0,220,0,0,0,168,0,114,0,232,0,124,0,172,0,55,0,122,0,0,0,0,0,153,0,148,0,101,0,0,0,69,0,132,0,0,0,0,0,140,0,1,0,0,0,67,0,195,0,200,0,169,0,58,0,52,0,64,0,162,0,0,0,15,0,100,0,69,0,76,0,95,0,176,0,185,0,132,0,251,0,75,0,57,0,78,0,237,0,35,0,120,0,189,0,244,0,18,0,72,0,201,0,154,0,76,0,255,0,2,0,56,0,0,0,0,0,191,0,150,0,1,0,0,0,196,0,244,0,128,0,115,0,9,0,0,0,242,0,99,0,245,0,49,0,187,0,165,0,123,0,182,0,126,0,75,0,173,0,0,0,250,0,155,0,57,0,63,0,76,0,217,0,244,0,2,0,0,0,0,0,77,0,0,0,163,0,27,0,0,0,0,0,195,0,225,0,0,0,129,0,92,0,0,0,142,0,220,0,205,0,118,0,73,0,95,0,103,0,154,0,142,0,64,0,168,0,0,0,71,0,74,0,6,0,94,0,76,0,124,0,43,0,33,0,192,0,98,0,156,0,0,0,180,0,100,0,81,0,206,0,124,0,0,0,0,0,0,0,7,0,14,0,0,0,0,0,1,0,56,0,40,0,212,0,58,0,74,0,152,0,176,0,24,0,206,0,248,0,33,0,165,0,178,0,13,0,255,0,192,0,180,0,160,0,0,0,2,0,98,0,225,0,0,0,79,0,49,0,117,0,148,0,0,0,68,0,42,0,254,0,122,0,0,0,120,0,254,0,99,0,173,0,54,0,0,0,83,0,199,0,220,0,133,0,225,0,255,0,0,0,110,0,244,0,239,0,182,0,137,0,106,0,0,0,179,0,213,0,61,0,78,0,194,0,164,0,4,0,87,0,0,0,161,0,107,0,49,0,0,0,144,0,120,0,162,0,125,0,0,0,75,0,252,0,0,0,85,0,216,0,163,0,205,0,0,0,225,0,218,0,0,0,82,0,235,0,77,0,0,0,175,0,82,0,0,0,27,0,0,0,85,0,161,0,124,0,90,0,178,0,3,0,197,0,247,0);
signal scenario_full  : scenario_type := (0,0,7,31,128,31,102,31,83,31,83,30,230,31,4,31,69,31,88,31,95,31,138,31,161,31,111,31,111,30,111,29,45,31,148,31,230,31,8,31,159,31,214,31,163,31,75,31,62,31,62,30,25,31,168,31,168,30,28,31,139,31,139,30,37,31,183,31,77,31,78,31,78,30,78,29,173,31,71,31,71,30,20,31,20,30,27,31,130,31,18,31,36,31,36,30,227,31,93,31,147,31,147,30,33,31,39,31,184,31,184,30,184,29,85,31,85,31,85,30,85,29,185,31,255,31,255,30,119,31,119,30,41,31,182,31,231,31,120,31,242,31,242,30,242,31,41,31,111,31,111,30,91,31,91,30,233,31,233,30,233,29,209,31,209,30,33,31,158,31,51,31,182,31,171,31,119,31,90,31,203,31,55,31,194,31,122,31,207,31,170,31,206,31,186,31,207,31,8,31,43,31,70,31,70,30,79,31,31,31,144,31,4,31,51,31,138,31,107,31,21,31,15,31,72,31,149,31,130,31,151,31,232,31,76,31,195,31,194,31,158,31,109,31,238,31,238,30,238,29,238,28,183,31,205,31,58,31,131,31,141,31,4,31,4,30,198,31,126,31,26,31,175,31,149,31,243,31,205,31,202,31,220,31,228,31,118,31,102,31,102,30,228,31,200,31,116,31,241,31,118,31,174,31,174,30,174,29,49,31,238,31,249,31,19,31,176,31,176,30,21,31,246,31,59,31,59,30,175,31,87,31,215,31,4,31,4,30,124,31,124,30,166,31,233,31,12,31,87,31,245,31,88,31,56,31,124,31,85,31,76,31,170,31,76,31,157,31,157,30,120,31,11,31,11,30,11,29,14,31,130,31,130,30,130,29,202,31,202,30,194,31,206,31,206,30,126,31,186,31,203,31,150,31,124,31,167,31,89,31,163,31,163,30,163,29,163,28,88,31,52,31,139,31,186,31,252,31,37,31,27,31,27,30,68,31,68,30,68,29,68,28,100,31,82,31,103,31,103,30,118,31,159,31,223,31,196,31,168,31,48,31,48,31,4,31,144,31,139,31,143,31,143,30,22,31,147,31,221,31,150,31,10,31,103,31,61,31,92,31,236,31,44,31,110,31,3,31,3,30,120,31,20,31,199,31,199,30,199,29,199,28,181,31,61,31,254,31,85,31,37,31,180,31,185,31,185,30,185,29,114,31,124,31,124,30,49,31,212,31,212,30,248,31,248,30,149,31,235,31,235,30,38,31,222,31,227,31,214,31,4,31,64,31,87,31,6,31,85,31,59,31,138,31,230,31,241,31,144,31,20,31,197,31,206,31,206,30,128,31,195,31,7,31,73,31,73,30,50,31,50,30,227,31,163,31,33,31,161,31,161,30,156,31,74,31,74,31,160,31,98,31,202,31,214,31,222,31,209,31,193,31,71,31,40,31,94,31,38,31,221,31,97,31,201,31,44,31,222,31,36,31,167,31,167,30,157,31,82,31,231,31,198,31,198,30,172,31,172,30,149,31,235,31,99,31,16,31,60,31,184,31,139,31,99,31,230,31,135,31,146,31,212,31,93,31,93,30,232,31,211,31,14,31,14,30,158,31,230,31,221,31,40,31,40,30,158,31,33,31,33,30,66,31,214,31,6,31,110,31,63,31,15,31,232,31,78,31,133,31,65,31,65,30,223,31,62,31,114,31,23,31,23,30,93,31,74,31,173,31,173,30,81,31,223,31,207,31,191,31,154,31,131,31,148,31,156,31,156,30,251,31,254,31,158,31,243,31,137,31,112,31,54,31,7,31,191,31,191,30,15,31,63,31,100,31,208,31,67,31,233,31,233,30,242,31,141,31,141,30,166,31,106,31,106,30,41,31,98,31,26,31,142,31,142,30,216,31,239,31,118,31,11,31,38,31,46,31,46,30,201,31,201,30,61,31,202,31,41,31,41,30,41,29,221,31,95,31,95,30,229,31,222,31,222,30,48,31,44,31,178,31,107,31,98,31,98,30,98,29,4,31,25,31,25,30,84,31,46,31,233,31,76,31,231,31,150,31,65,31,253,31,213,31,186,31,177,31,106,31,160,31,160,30,247,31,247,30,86,31,248,31,111,31,178,31,51,31,152,31,122,31,122,30,112,31,152,31,22,31,227,31,131,31,192,31,192,30,220,31,220,30,168,31,114,31,232,31,124,31,172,31,55,31,122,31,122,30,122,29,153,31,148,31,101,31,101,30,69,31,132,31,132,30,132,29,140,31,1,31,1,30,67,31,195,31,200,31,169,31,58,31,52,31,64,31,162,31,162,30,15,31,100,31,69,31,76,31,95,31,176,31,185,31,132,31,251,31,75,31,57,31,78,31,237,31,35,31,120,31,189,31,244,31,18,31,72,31,201,31,154,31,76,31,255,31,2,31,56,31,56,30,56,29,191,31,150,31,1,31,1,30,196,31,244,31,128,31,115,31,9,31,9,30,242,31,99,31,245,31,49,31,187,31,165,31,123,31,182,31,126,31,75,31,173,31,173,30,250,31,155,31,57,31,63,31,76,31,217,31,244,31,2,31,2,30,2,29,77,31,77,30,163,31,27,31,27,30,27,29,195,31,225,31,225,30,129,31,92,31,92,30,142,31,220,31,205,31,118,31,73,31,95,31,103,31,154,31,142,31,64,31,168,31,168,30,71,31,74,31,6,31,94,31,76,31,124,31,43,31,33,31,192,31,98,31,156,31,156,30,180,31,100,31,81,31,206,31,124,31,124,30,124,29,124,28,7,31,14,31,14,30,14,29,1,31,56,31,40,31,212,31,58,31,74,31,152,31,176,31,24,31,206,31,248,31,33,31,165,31,178,31,13,31,255,31,192,31,180,31,160,31,160,30,2,31,98,31,225,31,225,30,79,31,49,31,117,31,148,31,148,30,68,31,42,31,254,31,122,31,122,30,120,31,254,31,99,31,173,31,54,31,54,30,83,31,199,31,220,31,133,31,225,31,255,31,255,30,110,31,244,31,239,31,182,31,137,31,106,31,106,30,179,31,213,31,61,31,78,31,194,31,164,31,4,31,87,31,87,30,161,31,107,31,49,31,49,30,144,31,120,31,162,31,125,31,125,30,75,31,252,31,252,30,85,31,216,31,163,31,205,31,205,30,225,31,218,31,218,30,82,31,235,31,77,31,77,30,175,31,82,31,82,30,27,31,27,30,85,31,161,31,124,31,90,31,178,31,3,31,197,31,247,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
