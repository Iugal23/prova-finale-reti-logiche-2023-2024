-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1018;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (78,0,87,0,133,0,0,0,106,0,207,0,101,0,110,0,0,0,51,0,198,0,39,0,168,0,134,0,8,0,104,0,24,0,0,0,228,0,97,0,251,0,170,0,142,0,202,0,217,0,0,0,164,0,236,0,0,0,233,0,185,0,240,0,211,0,23,0,59,0,58,0,52,0,110,0,164,0,200,0,0,0,101,0,212,0,241,0,187,0,195,0,25,0,91,0,0,0,1,0,10,0,144,0,145,0,143,0,3,0,247,0,0,0,0,0,160,0,0,0,114,0,173,0,87,0,0,0,237,0,0,0,161,0,0,0,42,0,68,0,209,0,156,0,242,0,102,0,61,0,239,0,28,0,47,0,200,0,64,0,17,0,210,0,50,0,0,0,117,0,49,0,210,0,13,0,109,0,151,0,226,0,112,0,11,0,118,0,71,0,232,0,84,0,0,0,187,0,95,0,102,0,0,0,67,0,224,0,197,0,130,0,109,0,0,0,0,0,181,0,0,0,152,0,127,0,0,0,144,0,49,0,61,0,109,0,88,0,0,0,192,0,99,0,147,0,111,0,245,0,0,0,82,0,255,0,27,0,197,0,0,0,0,0,115,0,109,0,142,0,7,0,0,0,0,0,0,0,142,0,0,0,191,0,75,0,0,0,27,0,138,0,240,0,48,0,28,0,99,0,0,0,235,0,225,0,208,0,7,0,109,0,48,0,250,0,157,0,0,0,0,0,203,0,53,0,105,0,65,0,73,0,180,0,0,0,71,0,0,0,210,0,0,0,77,0,0,0,21,0,185,0,0,0,196,0,155,0,163,0,193,0,46,0,65,0,176,0,228,0,219,0,37,0,29,0,187,0,52,0,91,0,40,0,133,0,219,0,35,0,0,0,0,0,243,0,0,0,173,0,0,0,134,0,34,0,32,0,74,0,198,0,31,0,0,0,69,0,136,0,23,0,219,0,0,0,228,0,144,0,217,0,0,0,221,0,24,0,17,0,145,0,2,0,0,0,135,0,66,0,84,0,0,0,184,0,234,0,7,0,151,0,39,0,255,0,140,0,0,0,47,0,87,0,40,0,94,0,20,0,132,0,0,0,203,0,45,0,167,0,105,0,36,0,43,0,237,0,147,0,120,0,160,0,28,0,132,0,0,0,187,0,138,0,0,0,232,0,120,0,178,0,124,0,63,0,35,0,132,0,86,0,118,0,9,0,0,0,176,0,246,0,159,0,153,0,152,0,43,0,195,0,159,0,245,0,0,0,61,0,0,0,54,0,127,0,130,0,70,0,101,0,179,0,94,0,155,0,0,0,255,0,203,0,241,0,218,0,229,0,235,0,137,0,162,0,129,0,37,0,0,0,199,0,56,0,10,0,136,0,179,0,231,0,201,0,40,0,0,0,244,0,20,0,254,0,57,0,205,0,126,0,175,0,38,0,64,0,0,0,0,0,7,0,0,0,0,0,205,0,97,0,123,0,64,0,177,0,206,0,37,0,43,0,0,0,111,0,227,0,132,0,198,0,106,0,71,0,51,0,44,0,105,0,76,0,236,0,0,0,189,0,34,0,240,0,42,0,14,0,119,0,81,0,86,0,198,0,227,0,33,0,0,0,117,0,252,0,0,0,90,0,193,0,36,0,209,0,0,0,0,0,93,0,161,0,194,0,8,0,13,0,0,0,170,0,222,0,12,0,147,0,22,0,184,0,115,0,113,0,130,0,177,0,172,0,64,0,0,0,0,0,204,0,234,0,87,0,248,0,61,0,84,0,112,0,242,0,116,0,138,0,158,0,225,0,136,0,164,0,155,0,194,0,0,0,34,0,174,0,90,0,128,0,85,0,0,0,199,0,30,0,68,0,66,0,250,0,40,0,1,0,0,0,62,0,222,0,133,0,148,0,176,0,38,0,72,0,187,0,115,0,163,0,0,0,0,0,64,0,0,0,200,0,234,0,112,0,115,0,37,0,246,0,0,0,0,0,0,0,74,0,171,0,0,0,80,0,106,0,247,0,0,0,0,0,76,0,138,0,148,0,120,0,0,0,34,0,0,0,164,0,238,0,246,0,145,0,177,0,0,0,0,0,98,0,77,0,7,0,164,0,16,0,164,0,72,0,224,0,130,0,64,0,5,0,236,0,0,0,226,0,171,0,81,0,0,0,244,0,93,0,143,0,170,0,0,0,0,0,221,0,0,0,11,0,0,0,248,0,178,0,231,0,181,0,0,0,175,0,66,0,104,0,182,0,0,0,143,0,227,0,82,0,0,0,19,0,248,0,0,0,0,0,0,0,33,0,152,0,0,0,103,0,19,0,86,0,172,0,0,0,218,0,97,0,113,0,0,0,63,0,142,0,0,0,0,0,0,0,103,0,174,0,65,0,0,0,202,0,0,0,0,0,124,0,129,0,236,0,249,0,250,0,0,0,127,0,0,0,135,0,124,0,0,0,59,0,232,0,26,0,105,0,178,0,0,0,56,0,0,0,101,0,0,0,71,0,0,0,197,0,200,0,45,0,72,0,3,0,211,0,232,0,0,0,0,0,30,0,229,0,117,0,154,0,53,0,0,0,55,0,208,0,0,0,152,0,158,0,178,0,146,0,12,0,0,0,94,0,68,0,0,0,155,0,147,0,0,0,0,0,96,0,0,0,87,0,0,0,105,0,64,0,145,0,92,0,0,0,0,0,243,0,41,0,0,0,226,0,96,0,184,0,0,0,45,0,48,0,0,0,75,0,96,0,0,0,195,0,230,0,239,0,0,0,11,0,156,0,27,0,185,0,176,0,242,0,222,0,176,0,224,0,138,0,191,0,57,0,102,0,184,0,234,0,91,0,79,0,0,0,128,0,151,0,105,0,109,0,27,0,33,0,78,0,72,0,35,0,37,0,0,0,5,0,25,0,210,0,103,0,37,0,0,0,242,0,98,0,169,0,29,0,224,0,0,0,27,0,149,0,55,0,0,0,201,0,17,0,42,0,102,0,55,0,227,0,224,0,69,0,104,0,36,0,43,0,139,0,64,0,49,0,183,0,164,0,140,0,128,0,0,0,6,0,243,0,71,0,128,0,71,0,5,0,148,0,0,0,237,0,0,0,220,0,252,0,116,0,0,0,221,0,152,0,0,0,243,0,88,0,239,0,228,0,227,0,209,0,18,0,0,0,84,0,0,0,86,0,0,0,0,0,201,0,84,0,174,0,255,0,159,0,86,0,230,0,239,0,93,0,134,0,245,0,116,0,89,0,226,0,120,0,234,0,117,0,223,0,113,0,93,0,178,0,132,0,102,0,36,0,133,0,34,0,253,0,0,0,88,0,0,0,8,0,107,0,7,0,0,0,184,0,85,0,35,0,255,0,25,0,193,0,0,0,15,0,253,0,0,0,0,0,0,0,221,0,2,0,136,0,186,0,6,0,175,0,19,0,0,0,0,0,107,0,165,0,51,0,0,0,0,0,102,0,47,0,137,0,92,0,0,0,120,0,41,0,177,0,141,0,0,0,16,0,0,0,99,0,49,0,0,0,214,0,160,0,232,0,107,0,215,0,51,0,195,0,194,0,110,0,133,0,106,0,16,0,208,0,249,0,34,0,171,0,24,0,236,0,0,0,28,0,0,0,0,0,0,0,0,0,0,0,0,0,61,0,229,0,76,0,194,0,233,0,8,0,0,0,202,0,0,0,127,0,0,0,159,0,0,0,0,0,48,0,237,0,206,0,141,0,52,0,198,0,0,0,150,0,0,0,221,0,44,0,0,0,141,0,25,0,163,0,40,0,38,0,0,0,0,0,38,0,253,0,150,0,197,0,183,0,10,0,227,0,178,0,56,0,54,0,31,0,19,0,21,0,213,0,26,0,239,0,0,0,190,0,232,0,17,0,45,0,92,0,42,0,152,0,50,0,136,0,163,0,228,0,0,0,167,0,182,0,112,0,219,0,67,0,75,0,180,0,50,0,2,0,166,0,0,0,197,0,60,0,7,0,19,0,247,0,129,0,11,0,48,0,58,0,180,0,160,0,169,0,57,0,0,0,113,0,4,0,218,0,215,0,166,0,148,0,0,0,45,0,0,0,38,0,55,0,153,0,109,0,28,0,0,0,0,0,4,0,237,0,176,0,0,0,0,0,154,0,92,0,240,0,143,0,41,0,187,0,0,0,105,0,254,0,79,0,0,0,0,0,0,0,11,0,77,0,0,0,161,0,128,0,163,0,237,0,218,0,6,0,229,0,119,0,95,0,213,0,130,0,0,0,0,0,179,0,170,0,203,0,0,0,12,0,206,0,202,0,139,0,84,0,152,0,108,0,150,0,129,0,0,0,1,0,0,0,0,0,157,0,0,0,125,0,156,0,255,0,0,0,229,0,0,0,120,0,197,0,150,0,107,0,28,0,13,0,89,0,0,0,67,0,54,0,255,0,0,0,144,0,184,0,73,0,70,0,165,0,249,0,105,0,226,0,159,0,247,0,22,0,14,0,44,0,123,0,143,0,241,0,252,0,159,0,194,0,110,0,79,0,33,0,210,0,66,0,0,0,0,0,0,0,129,0,93,0,168,0,11,0,10,0,179,0,170,0,0,0,112,0);
signal scenario_full  : scenario_type := (78,31,87,31,133,31,133,30,106,31,207,31,101,31,110,31,110,30,51,31,198,31,39,31,168,31,134,31,8,31,104,31,24,31,24,30,228,31,97,31,251,31,170,31,142,31,202,31,217,31,217,30,164,31,236,31,236,30,233,31,185,31,240,31,211,31,23,31,59,31,58,31,52,31,110,31,164,31,200,31,200,30,101,31,212,31,241,31,187,31,195,31,25,31,91,31,91,30,1,31,10,31,144,31,145,31,143,31,3,31,247,31,247,30,247,29,160,31,160,30,114,31,173,31,87,31,87,30,237,31,237,30,161,31,161,30,42,31,68,31,209,31,156,31,242,31,102,31,61,31,239,31,28,31,47,31,200,31,64,31,17,31,210,31,50,31,50,30,117,31,49,31,210,31,13,31,109,31,151,31,226,31,112,31,11,31,118,31,71,31,232,31,84,31,84,30,187,31,95,31,102,31,102,30,67,31,224,31,197,31,130,31,109,31,109,30,109,29,181,31,181,30,152,31,127,31,127,30,144,31,49,31,61,31,109,31,88,31,88,30,192,31,99,31,147,31,111,31,245,31,245,30,82,31,255,31,27,31,197,31,197,30,197,29,115,31,109,31,142,31,7,31,7,30,7,29,7,28,142,31,142,30,191,31,75,31,75,30,27,31,138,31,240,31,48,31,28,31,99,31,99,30,235,31,225,31,208,31,7,31,109,31,48,31,250,31,157,31,157,30,157,29,203,31,53,31,105,31,65,31,73,31,180,31,180,30,71,31,71,30,210,31,210,30,77,31,77,30,21,31,185,31,185,30,196,31,155,31,163,31,193,31,46,31,65,31,176,31,228,31,219,31,37,31,29,31,187,31,52,31,91,31,40,31,133,31,219,31,35,31,35,30,35,29,243,31,243,30,173,31,173,30,134,31,34,31,32,31,74,31,198,31,31,31,31,30,69,31,136,31,23,31,219,31,219,30,228,31,144,31,217,31,217,30,221,31,24,31,17,31,145,31,2,31,2,30,135,31,66,31,84,31,84,30,184,31,234,31,7,31,151,31,39,31,255,31,140,31,140,30,47,31,87,31,40,31,94,31,20,31,132,31,132,30,203,31,45,31,167,31,105,31,36,31,43,31,237,31,147,31,120,31,160,31,28,31,132,31,132,30,187,31,138,31,138,30,232,31,120,31,178,31,124,31,63,31,35,31,132,31,86,31,118,31,9,31,9,30,176,31,246,31,159,31,153,31,152,31,43,31,195,31,159,31,245,31,245,30,61,31,61,30,54,31,127,31,130,31,70,31,101,31,179,31,94,31,155,31,155,30,255,31,203,31,241,31,218,31,229,31,235,31,137,31,162,31,129,31,37,31,37,30,199,31,56,31,10,31,136,31,179,31,231,31,201,31,40,31,40,30,244,31,20,31,254,31,57,31,205,31,126,31,175,31,38,31,64,31,64,30,64,29,7,31,7,30,7,29,205,31,97,31,123,31,64,31,177,31,206,31,37,31,43,31,43,30,111,31,227,31,132,31,198,31,106,31,71,31,51,31,44,31,105,31,76,31,236,31,236,30,189,31,34,31,240,31,42,31,14,31,119,31,81,31,86,31,198,31,227,31,33,31,33,30,117,31,252,31,252,30,90,31,193,31,36,31,209,31,209,30,209,29,93,31,161,31,194,31,8,31,13,31,13,30,170,31,222,31,12,31,147,31,22,31,184,31,115,31,113,31,130,31,177,31,172,31,64,31,64,30,64,29,204,31,234,31,87,31,248,31,61,31,84,31,112,31,242,31,116,31,138,31,158,31,225,31,136,31,164,31,155,31,194,31,194,30,34,31,174,31,90,31,128,31,85,31,85,30,199,31,30,31,68,31,66,31,250,31,40,31,1,31,1,30,62,31,222,31,133,31,148,31,176,31,38,31,72,31,187,31,115,31,163,31,163,30,163,29,64,31,64,30,200,31,234,31,112,31,115,31,37,31,246,31,246,30,246,29,246,28,74,31,171,31,171,30,80,31,106,31,247,31,247,30,247,29,76,31,138,31,148,31,120,31,120,30,34,31,34,30,164,31,238,31,246,31,145,31,177,31,177,30,177,29,98,31,77,31,7,31,164,31,16,31,164,31,72,31,224,31,130,31,64,31,5,31,236,31,236,30,226,31,171,31,81,31,81,30,244,31,93,31,143,31,170,31,170,30,170,29,221,31,221,30,11,31,11,30,248,31,178,31,231,31,181,31,181,30,175,31,66,31,104,31,182,31,182,30,143,31,227,31,82,31,82,30,19,31,248,31,248,30,248,29,248,28,33,31,152,31,152,30,103,31,19,31,86,31,172,31,172,30,218,31,97,31,113,31,113,30,63,31,142,31,142,30,142,29,142,28,103,31,174,31,65,31,65,30,202,31,202,30,202,29,124,31,129,31,236,31,249,31,250,31,250,30,127,31,127,30,135,31,124,31,124,30,59,31,232,31,26,31,105,31,178,31,178,30,56,31,56,30,101,31,101,30,71,31,71,30,197,31,200,31,45,31,72,31,3,31,211,31,232,31,232,30,232,29,30,31,229,31,117,31,154,31,53,31,53,30,55,31,208,31,208,30,152,31,158,31,178,31,146,31,12,31,12,30,94,31,68,31,68,30,155,31,147,31,147,30,147,29,96,31,96,30,87,31,87,30,105,31,64,31,145,31,92,31,92,30,92,29,243,31,41,31,41,30,226,31,96,31,184,31,184,30,45,31,48,31,48,30,75,31,96,31,96,30,195,31,230,31,239,31,239,30,11,31,156,31,27,31,185,31,176,31,242,31,222,31,176,31,224,31,138,31,191,31,57,31,102,31,184,31,234,31,91,31,79,31,79,30,128,31,151,31,105,31,109,31,27,31,33,31,78,31,72,31,35,31,37,31,37,30,5,31,25,31,210,31,103,31,37,31,37,30,242,31,98,31,169,31,29,31,224,31,224,30,27,31,149,31,55,31,55,30,201,31,17,31,42,31,102,31,55,31,227,31,224,31,69,31,104,31,36,31,43,31,139,31,64,31,49,31,183,31,164,31,140,31,128,31,128,30,6,31,243,31,71,31,128,31,71,31,5,31,148,31,148,30,237,31,237,30,220,31,252,31,116,31,116,30,221,31,152,31,152,30,243,31,88,31,239,31,228,31,227,31,209,31,18,31,18,30,84,31,84,30,86,31,86,30,86,29,201,31,84,31,174,31,255,31,159,31,86,31,230,31,239,31,93,31,134,31,245,31,116,31,89,31,226,31,120,31,234,31,117,31,223,31,113,31,93,31,178,31,132,31,102,31,36,31,133,31,34,31,253,31,253,30,88,31,88,30,8,31,107,31,7,31,7,30,184,31,85,31,35,31,255,31,25,31,193,31,193,30,15,31,253,31,253,30,253,29,253,28,221,31,2,31,136,31,186,31,6,31,175,31,19,31,19,30,19,29,107,31,165,31,51,31,51,30,51,29,102,31,47,31,137,31,92,31,92,30,120,31,41,31,177,31,141,31,141,30,16,31,16,30,99,31,49,31,49,30,214,31,160,31,232,31,107,31,215,31,51,31,195,31,194,31,110,31,133,31,106,31,16,31,208,31,249,31,34,31,171,31,24,31,236,31,236,30,28,31,28,30,28,29,28,28,28,27,28,26,28,25,61,31,229,31,76,31,194,31,233,31,8,31,8,30,202,31,202,30,127,31,127,30,159,31,159,30,159,29,48,31,237,31,206,31,141,31,52,31,198,31,198,30,150,31,150,30,221,31,44,31,44,30,141,31,25,31,163,31,40,31,38,31,38,30,38,29,38,31,253,31,150,31,197,31,183,31,10,31,227,31,178,31,56,31,54,31,31,31,19,31,21,31,213,31,26,31,239,31,239,30,190,31,232,31,17,31,45,31,92,31,42,31,152,31,50,31,136,31,163,31,228,31,228,30,167,31,182,31,112,31,219,31,67,31,75,31,180,31,50,31,2,31,166,31,166,30,197,31,60,31,7,31,19,31,247,31,129,31,11,31,48,31,58,31,180,31,160,31,169,31,57,31,57,30,113,31,4,31,218,31,215,31,166,31,148,31,148,30,45,31,45,30,38,31,55,31,153,31,109,31,28,31,28,30,28,29,4,31,237,31,176,31,176,30,176,29,154,31,92,31,240,31,143,31,41,31,187,31,187,30,105,31,254,31,79,31,79,30,79,29,79,28,11,31,77,31,77,30,161,31,128,31,163,31,237,31,218,31,6,31,229,31,119,31,95,31,213,31,130,31,130,30,130,29,179,31,170,31,203,31,203,30,12,31,206,31,202,31,139,31,84,31,152,31,108,31,150,31,129,31,129,30,1,31,1,30,1,29,157,31,157,30,125,31,156,31,255,31,255,30,229,31,229,30,120,31,197,31,150,31,107,31,28,31,13,31,89,31,89,30,67,31,54,31,255,31,255,30,144,31,184,31,73,31,70,31,165,31,249,31,105,31,226,31,159,31,247,31,22,31,14,31,44,31,123,31,143,31,241,31,252,31,159,31,194,31,110,31,79,31,33,31,210,31,66,31,66,30,66,29,66,28,129,31,93,31,168,31,11,31,10,31,179,31,170,31,170,30,112,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
