-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_735 is
end project_tb_735;

architecture project_tb_arch_735 of project_tb_735 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 621;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (71,0,215,0,254,0,181,0,66,0,172,0,204,0,0,0,53,0,46,0,238,0,77,0,162,0,9,0,0,0,128,0,173,0,132,0,80,0,201,0,4,0,0,0,0,0,140,0,136,0,0,0,247,0,51,0,163,0,218,0,0,0,214,0,188,0,30,0,0,0,47,0,169,0,13,0,190,0,23,0,29,0,196,0,120,0,114,0,138,0,131,0,170,0,0,0,150,0,239,0,77,0,254,0,218,0,0,0,126,0,20,0,0,0,155,0,40,0,154,0,0,0,0,0,0,0,111,0,63,0,185,0,0,0,0,0,3,0,217,0,0,0,0,0,0,0,245,0,185,0,165,0,0,0,223,0,0,0,203,0,199,0,248,0,118,0,251,0,112,0,115,0,199,0,251,0,173,0,0,0,160,0,0,0,163,0,63,0,76,0,38,0,154,0,103,0,107,0,239,0,164,0,0,0,0,0,29,0,0,0,24,0,142,0,222,0,105,0,246,0,250,0,241,0,231,0,0,0,231,0,91,0,110,0,0,0,0,0,46,0,248,0,165,0,77,0,127,0,253,0,83,0,202,0,237,0,44,0,159,0,132,0,227,0,190,0,203,0,121,0,75,0,6,0,33,0,228,0,44,0,0,0,34,0,189,0,167,0,254,0,238,0,198,0,0,0,174,0,0,0,37,0,52,0,134,0,102,0,0,0,22,0,0,0,6,0,120,0,0,0,28,0,242,0,179,0,76,0,140,0,0,0,91,0,0,0,166,0,138,0,198,0,100,0,230,0,85,0,156,0,3,0,69,0,237,0,28,0,48,0,132,0,93,0,100,0,196,0,5,0,105,0,0,0,180,0,183,0,0,0,219,0,104,0,0,0,78,0,0,0,84,0,138,0,223,0,0,0,0,0,0,0,194,0,190,0,0,0,0,0,177,0,165,0,89,0,137,0,2,0,236,0,159,0,43,0,127,0,159,0,148,0,227,0,124,0,65,0,58,0,132,0,206,0,143,0,0,0,240,0,193,0,33,0,126,0,148,0,127,0,0,0,16,0,21,0,56,0,72,0,210,0,202,0,176,0,97,0,141,0,148,0,184,0,117,0,129,0,221,0,0,0,0,0,216,0,78,0,0,0,0,0,197,0,183,0,0,0,163,0,36,0,207,0,0,0,18,0,0,0,0,0,19,0,107,0,67,0,133,0,228,0,27,0,190,0,197,0,239,0,89,0,202,0,176,0,172,0,19,0,35,0,233,0,186,0,255,0,229,0,39,0,133,0,83,0,0,0,0,0,103,0,0,0,228,0,202,0,0,0,105,0,0,0,122,0,217,0,188,0,171,0,187,0,0,0,134,0,66,0,0,0,0,0,0,0,232,0,150,0,0,0,0,0,14,0,92,0,154,0,183,0,19,0,0,0,6,0,234,0,150,0,0,0,86,0,71,0,89,0,63,0,2,0,121,0,49,0,0,0,201,0,249,0,0,0,21,0,58,0,96,0,92,0,114,0,74,0,210,0,159,0,38,0,118,0,191,0,204,0,57,0,210,0,207,0,0,0,0,0,66,0,143,0,129,0,0,0,206,0,100,0,11,0,136,0,30,0,0,0,65,0,0,0,160,0,0,0,240,0,18,0,255,0,0,0,98,0,34,0,0,0,44,0,7,0,200,0,56,0,247,0,183,0,166,0,84,0,106,0,74,0,166,0,137,0,57,0,191,0,157,0,0,0,48,0,0,0,114,0,0,0,54,0,119,0,232,0,196,0,254,0,29,0,171,0,120,0,105,0,146,0,169,0,116,0,110,0,206,0,143,0,177,0,191,0,77,0,0,0,66,0,150,0,0,0,36,0,142,0,178,0,204,0,234,0,95,0,99,0,104,0,0,0,131,0,62,0,0,0,0,0,135,0,0,0,184,0,252,0,16,0,0,0,142,0,208,0,0,0,94,0,0,0,38,0,80,0,15,0,107,0,66,0,236,0,136,0,0,0,51,0,154,0,99,0,85,0,124,0,244,0,225,0,0,0,0,0,86,0,91,0,164,0,206,0,0,0,234,0,217,0,57,0,198,0,194,0,0,0,61,0,72,0,246,0,89,0,0,0,131,0,62,0,41,0,240,0,94,0,221,0,0,0,79,0,0,0,154,0,117,0,41,0,73,0,0,0,203,0,96,0,255,0,140,0,163,0,69,0,35,0,233,0,211,0,219,0,126,0,102,0,109,0,27,0,0,0,116,0,65,0,12,0,0,0,0,0,205,0,0,0,167,0,93,0,137,0,0,0,245,0,0,0,0,0,249,0,159,0,30,0,69,0,0,0,0,0,0,0,232,0,230,0,238,0,247,0,1,0,207,0,89,0,91,0,212,0,31,0,50,0,213,0,157,0,17,0,94,0,0,0,20,0,140,0,211,0,226,0,166,0,0,0,203,0,251,0,134,0,0,0,0,0,177,0,239,0,137,0,215,0,98,0,79,0,33,0,186,0,21,0,127,0,0,0,0,0,193,0,0,0,185,0,181,0,188,0,33,0,49,0,233,0,0,0,224,0,232,0,163,0,194,0,242,0,130,0,0,0,45,0,0,0,1,0,68,0,110,0,194,0,171,0,94,0,157,0,137,0,122,0,114,0,0,0,7,0,0,0,93,0,155,0,0,0,128,0,48,0,14,0,0,0,107,0,21,0,59,0,0,0,55,0,193,0,136,0,248,0,82,0,0,0,244,0,158,0,84,0,122,0,49,0,177,0,42,0,0,0,118,0,0,0,220,0,48,0,226,0,0,0,242,0,216,0,211,0,0,0,0,0);
signal scenario_full  : scenario_type := (71,31,215,31,254,31,181,31,66,31,172,31,204,31,204,30,53,31,46,31,238,31,77,31,162,31,9,31,9,30,128,31,173,31,132,31,80,31,201,31,4,31,4,30,4,29,140,31,136,31,136,30,247,31,51,31,163,31,218,31,218,30,214,31,188,31,30,31,30,30,47,31,169,31,13,31,190,31,23,31,29,31,196,31,120,31,114,31,138,31,131,31,170,31,170,30,150,31,239,31,77,31,254,31,218,31,218,30,126,31,20,31,20,30,155,31,40,31,154,31,154,30,154,29,154,28,111,31,63,31,185,31,185,30,185,29,3,31,217,31,217,30,217,29,217,28,245,31,185,31,165,31,165,30,223,31,223,30,203,31,199,31,248,31,118,31,251,31,112,31,115,31,199,31,251,31,173,31,173,30,160,31,160,30,163,31,63,31,76,31,38,31,154,31,103,31,107,31,239,31,164,31,164,30,164,29,29,31,29,30,24,31,142,31,222,31,105,31,246,31,250,31,241,31,231,31,231,30,231,31,91,31,110,31,110,30,110,29,46,31,248,31,165,31,77,31,127,31,253,31,83,31,202,31,237,31,44,31,159,31,132,31,227,31,190,31,203,31,121,31,75,31,6,31,33,31,228,31,44,31,44,30,34,31,189,31,167,31,254,31,238,31,198,31,198,30,174,31,174,30,37,31,52,31,134,31,102,31,102,30,22,31,22,30,6,31,120,31,120,30,28,31,242,31,179,31,76,31,140,31,140,30,91,31,91,30,166,31,138,31,198,31,100,31,230,31,85,31,156,31,3,31,69,31,237,31,28,31,48,31,132,31,93,31,100,31,196,31,5,31,105,31,105,30,180,31,183,31,183,30,219,31,104,31,104,30,78,31,78,30,84,31,138,31,223,31,223,30,223,29,223,28,194,31,190,31,190,30,190,29,177,31,165,31,89,31,137,31,2,31,236,31,159,31,43,31,127,31,159,31,148,31,227,31,124,31,65,31,58,31,132,31,206,31,143,31,143,30,240,31,193,31,33,31,126,31,148,31,127,31,127,30,16,31,21,31,56,31,72,31,210,31,202,31,176,31,97,31,141,31,148,31,184,31,117,31,129,31,221,31,221,30,221,29,216,31,78,31,78,30,78,29,197,31,183,31,183,30,163,31,36,31,207,31,207,30,18,31,18,30,18,29,19,31,107,31,67,31,133,31,228,31,27,31,190,31,197,31,239,31,89,31,202,31,176,31,172,31,19,31,35,31,233,31,186,31,255,31,229,31,39,31,133,31,83,31,83,30,83,29,103,31,103,30,228,31,202,31,202,30,105,31,105,30,122,31,217,31,188,31,171,31,187,31,187,30,134,31,66,31,66,30,66,29,66,28,232,31,150,31,150,30,150,29,14,31,92,31,154,31,183,31,19,31,19,30,6,31,234,31,150,31,150,30,86,31,71,31,89,31,63,31,2,31,121,31,49,31,49,30,201,31,249,31,249,30,21,31,58,31,96,31,92,31,114,31,74,31,210,31,159,31,38,31,118,31,191,31,204,31,57,31,210,31,207,31,207,30,207,29,66,31,143,31,129,31,129,30,206,31,100,31,11,31,136,31,30,31,30,30,65,31,65,30,160,31,160,30,240,31,18,31,255,31,255,30,98,31,34,31,34,30,44,31,7,31,200,31,56,31,247,31,183,31,166,31,84,31,106,31,74,31,166,31,137,31,57,31,191,31,157,31,157,30,48,31,48,30,114,31,114,30,54,31,119,31,232,31,196,31,254,31,29,31,171,31,120,31,105,31,146,31,169,31,116,31,110,31,206,31,143,31,177,31,191,31,77,31,77,30,66,31,150,31,150,30,36,31,142,31,178,31,204,31,234,31,95,31,99,31,104,31,104,30,131,31,62,31,62,30,62,29,135,31,135,30,184,31,252,31,16,31,16,30,142,31,208,31,208,30,94,31,94,30,38,31,80,31,15,31,107,31,66,31,236,31,136,31,136,30,51,31,154,31,99,31,85,31,124,31,244,31,225,31,225,30,225,29,86,31,91,31,164,31,206,31,206,30,234,31,217,31,57,31,198,31,194,31,194,30,61,31,72,31,246,31,89,31,89,30,131,31,62,31,41,31,240,31,94,31,221,31,221,30,79,31,79,30,154,31,117,31,41,31,73,31,73,30,203,31,96,31,255,31,140,31,163,31,69,31,35,31,233,31,211,31,219,31,126,31,102,31,109,31,27,31,27,30,116,31,65,31,12,31,12,30,12,29,205,31,205,30,167,31,93,31,137,31,137,30,245,31,245,30,245,29,249,31,159,31,30,31,69,31,69,30,69,29,69,28,232,31,230,31,238,31,247,31,1,31,207,31,89,31,91,31,212,31,31,31,50,31,213,31,157,31,17,31,94,31,94,30,20,31,140,31,211,31,226,31,166,31,166,30,203,31,251,31,134,31,134,30,134,29,177,31,239,31,137,31,215,31,98,31,79,31,33,31,186,31,21,31,127,31,127,30,127,29,193,31,193,30,185,31,181,31,188,31,33,31,49,31,233,31,233,30,224,31,232,31,163,31,194,31,242,31,130,31,130,30,45,31,45,30,1,31,68,31,110,31,194,31,171,31,94,31,157,31,137,31,122,31,114,31,114,30,7,31,7,30,93,31,155,31,155,30,128,31,48,31,14,31,14,30,107,31,21,31,59,31,59,30,55,31,193,31,136,31,248,31,82,31,82,30,244,31,158,31,84,31,122,31,49,31,177,31,42,31,42,30,118,31,118,30,220,31,48,31,226,31,226,30,242,31,216,31,211,31,211,30,211,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
