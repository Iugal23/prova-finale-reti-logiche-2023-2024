-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_486 is
end project_tb_486;

architecture project_tb_arch_486 of project_tb_486 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 783;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (93,0,202,0,183,0,0,0,252,0,0,0,144,0,146,0,155,0,224,0,211,0,59,0,0,0,238,0,138,0,97,0,143,0,116,0,72,0,0,0,38,0,0,0,0,0,203,0,191,0,62,0,202,0,58,0,0,0,0,0,244,0,49,0,16,0,253,0,230,0,54,0,88,0,108,0,55,0,149,0,62,0,164,0,58,0,0,0,106,0,61,0,172,0,6,0,0,0,66,0,153,0,182,0,242,0,137,0,77,0,0,0,59,0,156,0,101,0,0,0,0,0,161,0,116,0,179,0,89,0,109,0,56,0,207,0,140,0,90,0,84,0,0,0,65,0,30,0,98,0,200,0,179,0,94,0,145,0,85,0,0,0,253,0,0,0,102,0,0,0,220,0,249,0,154,0,213,0,141,0,146,0,104,0,0,0,208,0,142,0,208,0,147,0,202,0,209,0,0,0,81,0,208,0,96,0,0,0,125,0,79,0,0,0,82,0,0,0,234,0,128,0,0,0,219,0,221,0,211,0,0,0,0,0,160,0,57,0,200,0,145,0,142,0,6,0,47,0,55,0,49,0,230,0,52,0,0,0,0,0,20,0,120,0,226,0,223,0,0,0,27,0,142,0,98,0,75,0,110,0,90,0,233,0,16,0,199,0,154,0,255,0,123,0,240,0,12,0,0,0,156,0,108,0,17,0,28,0,164,0,182,0,40,0,7,0,0,0,0,0,243,0,0,0,31,0,132,0,87,0,0,0,123,0,76,0,90,0,100,0,146,0,105,0,209,0,70,0,0,0,203,0,190,0,71,0,183,0,186,0,137,0,0,0,148,0,55,0,241,0,168,0,188,0,56,0,0,0,194,0,169,0,0,0,31,0,0,0,42,0,220,0,90,0,21,0,0,0,154,0,60,0,0,0,0,0,123,0,136,0,147,0,131,0,117,0,74,0,171,0,0,0,108,0,192,0,249,0,124,0,145,0,97,0,145,0,0,0,14,0,25,0,154,0,239,0,183,0,249,0,0,0,107,0,63,0,78,0,112,0,178,0,222,0,5,0,62,0,134,0,219,0,251,0,78,0,158,0,28,0,95,0,0,0,54,0,187,0,158,0,33,0,52,0,0,0,155,0,0,0,236,0,233,0,237,0,116,0,195,0,65,0,215,0,116,0,17,0,82,0,207,0,101,0,89,0,0,0,0,0,135,0,0,0,0,0,0,0,90,0,73,0,120,0,193,0,78,0,249,0,0,0,214,0,246,0,0,0,249,0,145,0,0,0,95,0,101,0,173,0,102,0,106,0,236,0,0,0,18,0,20,0,0,0,0,0,0,0,0,0,24,0,94,0,0,0,27,0,16,0,143,0,65,0,187,0,0,0,109,0,218,0,125,0,16,0,23,0,6,0,218,0,2,0,53,0,236,0,108,0,0,0,52,0,255,0,3,0,82,0,126,0,0,0,144,0,62,0,239,0,197,0,84,0,0,0,242,0,100,0,208,0,99,0,211,0,180,0,225,0,0,0,113,0,60,0,129,0,0,0,2,0,126,0,13,0,152,0,0,0,92,0,0,0,102,0,197,0,134,0,157,0,0,0,128,0,0,0,0,0,9,0,66,0,43,0,249,0,0,0,63,0,36,0,0,0,38,0,0,0,121,0,37,0,205,0,26,0,0,0,4,0,130,0,63,0,13,0,28,0,190,0,208,0,0,0,30,0,12,0,208,0,24,0,53,0,54,0,0,0,149,0,0,0,0,0,213,0,102,0,17,0,0,0,72,0,121,0,77,0,119,0,227,0,114,0,70,0,241,0,0,0,143,0,238,0,0,0,15,0,0,0,182,0,55,0,250,0,168,0,113,0,0,0,245,0,8,0,236,0,100,0,255,0,204,0,183,0,139,0,0,0,0,0,32,0,147,0,1,0,18,0,117,0,203,0,174,0,21,0,0,0,207,0,195,0,112,0,6,0,213,0,56,0,182,0,0,0,3,0,178,0,173,0,86,0,172,0,0,0,151,0,198,0,172,0,125,0,79,0,0,0,114,0,77,0,93,0,180,0,50,0,0,0,0,0,0,0,114,0,87,0,0,0,134,0,0,0,119,0,30,0,178,0,14,0,112,0,246,0,0,0,124,0,213,0,212,0,0,0,0,0,0,0,57,0,198,0,58,0,0,0,74,0,0,0,26,0,33,0,59,0,196,0,0,0,216,0,138,0,33,0,29,0,131,0,240,0,0,0,0,0,241,0,189,0,13,0,130,0,0,0,180,0,0,0,0,0,16,0,0,0,16,0,185,0,83,0,97,0,235,0,67,0,86,0,0,0,232,0,0,0,0,0,251,0,151,0,240,0,0,0,148,0,0,0,62,0,0,0,51,0,144,0,181,0,47,0,0,0,254,0,203,0,0,0,51,0,129,0,0,0,8,0,166,0,222,0,183,0,128,0,152,0,176,0,178,0,234,0,80,0,9,0,0,0,97,0,140,0,14,0,0,0,41,0,0,0,236,0,250,0,37,0,18,0,174,0,236,0,137,0,205,0,233,0,22,0,227,0,2,0,136,0,58,0,89,0,170,0,9,0,71,0,242,0,5,0,225,0,118,0,247,0,61,0,10,0,165,0,143,0,19,0,226,0,76,0,232,0,247,0,74,0,238,0,0,0,48,0,43,0,0,0,32,0,53,0,4,0,205,0,79,0,43,0,4,0,0,0,56,0,0,0,92,0,133,0,74,0,72,0,253,0,176,0,51,0,0,0,2,0,177,0,176,0,156,0,250,0,0,0,0,0,165,0,193,0,0,0,160,0,73,0,0,0,186,0,173,0,229,0,0,0,0,0,0,0,150,0,161,0,219,0,21,0,253,0,46,0,236,0,30,0,0,0,65,0,213,0,22,0,135,0,35,0,113,0,67,0,163,0,22,0,4,0,11,0,135,0,40,0,215,0,0,0,42,0,0,0,46,0,201,0,0,0,223,0,131,0,165,0,130,0,0,0,0,0,7,0,251,0,64,0,39,0,70,0,87,0,122,0,246,0,174,0,227,0,0,0,163,0,185,0,23,0,113,0,0,0,97,0,0,0,202,0,182,0,165,0,41,0,64,0,173,0,0,0,240,0,41,0,177,0,0,0,0,0,42,0,0,0,62,0,0,0,0,0,3,0,0,0,0,0,233,0,23,0,171,0,42,0,231,0,144,0,0,0,45,0,2,0,173,0,206,0,128,0,42,0,206,0,190,0,0,0,15,0,134,0,19,0,234,0,58,0,176,0,169,0,234,0,26,0,49,0,246,0,0,0,209,0,132,0,84,0,200,0,93,0,0,0,96,0,208,0,100,0,0,0,203,0,242,0,1,0,0,0,207,0,123,0,0,0,199,0,42,0,29,0,179,0,140,0,201,0,222,0,0,0,0,0,146,0,210,0,176,0,253,0,96,0,114,0,218,0,247,0,173,0,69,0,156,0,2,0,185,0,134,0,230,0,229,0,209,0,129,0,0,0,3,0,70,0,211,0,202,0,0,0,40,0,225,0,58,0);
signal scenario_full  : scenario_type := (93,31,202,31,183,31,183,30,252,31,252,30,144,31,146,31,155,31,224,31,211,31,59,31,59,30,238,31,138,31,97,31,143,31,116,31,72,31,72,30,38,31,38,30,38,29,203,31,191,31,62,31,202,31,58,31,58,30,58,29,244,31,49,31,16,31,253,31,230,31,54,31,88,31,108,31,55,31,149,31,62,31,164,31,58,31,58,30,106,31,61,31,172,31,6,31,6,30,66,31,153,31,182,31,242,31,137,31,77,31,77,30,59,31,156,31,101,31,101,30,101,29,161,31,116,31,179,31,89,31,109,31,56,31,207,31,140,31,90,31,84,31,84,30,65,31,30,31,98,31,200,31,179,31,94,31,145,31,85,31,85,30,253,31,253,30,102,31,102,30,220,31,249,31,154,31,213,31,141,31,146,31,104,31,104,30,208,31,142,31,208,31,147,31,202,31,209,31,209,30,81,31,208,31,96,31,96,30,125,31,79,31,79,30,82,31,82,30,234,31,128,31,128,30,219,31,221,31,211,31,211,30,211,29,160,31,57,31,200,31,145,31,142,31,6,31,47,31,55,31,49,31,230,31,52,31,52,30,52,29,20,31,120,31,226,31,223,31,223,30,27,31,142,31,98,31,75,31,110,31,90,31,233,31,16,31,199,31,154,31,255,31,123,31,240,31,12,31,12,30,156,31,108,31,17,31,28,31,164,31,182,31,40,31,7,31,7,30,7,29,243,31,243,30,31,31,132,31,87,31,87,30,123,31,76,31,90,31,100,31,146,31,105,31,209,31,70,31,70,30,203,31,190,31,71,31,183,31,186,31,137,31,137,30,148,31,55,31,241,31,168,31,188,31,56,31,56,30,194,31,169,31,169,30,31,31,31,30,42,31,220,31,90,31,21,31,21,30,154,31,60,31,60,30,60,29,123,31,136,31,147,31,131,31,117,31,74,31,171,31,171,30,108,31,192,31,249,31,124,31,145,31,97,31,145,31,145,30,14,31,25,31,154,31,239,31,183,31,249,31,249,30,107,31,63,31,78,31,112,31,178,31,222,31,5,31,62,31,134,31,219,31,251,31,78,31,158,31,28,31,95,31,95,30,54,31,187,31,158,31,33,31,52,31,52,30,155,31,155,30,236,31,233,31,237,31,116,31,195,31,65,31,215,31,116,31,17,31,82,31,207,31,101,31,89,31,89,30,89,29,135,31,135,30,135,29,135,28,90,31,73,31,120,31,193,31,78,31,249,31,249,30,214,31,246,31,246,30,249,31,145,31,145,30,95,31,101,31,173,31,102,31,106,31,236,31,236,30,18,31,20,31,20,30,20,29,20,28,20,27,24,31,94,31,94,30,27,31,16,31,143,31,65,31,187,31,187,30,109,31,218,31,125,31,16,31,23,31,6,31,218,31,2,31,53,31,236,31,108,31,108,30,52,31,255,31,3,31,82,31,126,31,126,30,144,31,62,31,239,31,197,31,84,31,84,30,242,31,100,31,208,31,99,31,211,31,180,31,225,31,225,30,113,31,60,31,129,31,129,30,2,31,126,31,13,31,152,31,152,30,92,31,92,30,102,31,197,31,134,31,157,31,157,30,128,31,128,30,128,29,9,31,66,31,43,31,249,31,249,30,63,31,36,31,36,30,38,31,38,30,121,31,37,31,205,31,26,31,26,30,4,31,130,31,63,31,13,31,28,31,190,31,208,31,208,30,30,31,12,31,208,31,24,31,53,31,54,31,54,30,149,31,149,30,149,29,213,31,102,31,17,31,17,30,72,31,121,31,77,31,119,31,227,31,114,31,70,31,241,31,241,30,143,31,238,31,238,30,15,31,15,30,182,31,55,31,250,31,168,31,113,31,113,30,245,31,8,31,236,31,100,31,255,31,204,31,183,31,139,31,139,30,139,29,32,31,147,31,1,31,18,31,117,31,203,31,174,31,21,31,21,30,207,31,195,31,112,31,6,31,213,31,56,31,182,31,182,30,3,31,178,31,173,31,86,31,172,31,172,30,151,31,198,31,172,31,125,31,79,31,79,30,114,31,77,31,93,31,180,31,50,31,50,30,50,29,50,28,114,31,87,31,87,30,134,31,134,30,119,31,30,31,178,31,14,31,112,31,246,31,246,30,124,31,213,31,212,31,212,30,212,29,212,28,57,31,198,31,58,31,58,30,74,31,74,30,26,31,33,31,59,31,196,31,196,30,216,31,138,31,33,31,29,31,131,31,240,31,240,30,240,29,241,31,189,31,13,31,130,31,130,30,180,31,180,30,180,29,16,31,16,30,16,31,185,31,83,31,97,31,235,31,67,31,86,31,86,30,232,31,232,30,232,29,251,31,151,31,240,31,240,30,148,31,148,30,62,31,62,30,51,31,144,31,181,31,47,31,47,30,254,31,203,31,203,30,51,31,129,31,129,30,8,31,166,31,222,31,183,31,128,31,152,31,176,31,178,31,234,31,80,31,9,31,9,30,97,31,140,31,14,31,14,30,41,31,41,30,236,31,250,31,37,31,18,31,174,31,236,31,137,31,205,31,233,31,22,31,227,31,2,31,136,31,58,31,89,31,170,31,9,31,71,31,242,31,5,31,225,31,118,31,247,31,61,31,10,31,165,31,143,31,19,31,226,31,76,31,232,31,247,31,74,31,238,31,238,30,48,31,43,31,43,30,32,31,53,31,4,31,205,31,79,31,43,31,4,31,4,30,56,31,56,30,92,31,133,31,74,31,72,31,253,31,176,31,51,31,51,30,2,31,177,31,176,31,156,31,250,31,250,30,250,29,165,31,193,31,193,30,160,31,73,31,73,30,186,31,173,31,229,31,229,30,229,29,229,28,150,31,161,31,219,31,21,31,253,31,46,31,236,31,30,31,30,30,65,31,213,31,22,31,135,31,35,31,113,31,67,31,163,31,22,31,4,31,11,31,135,31,40,31,215,31,215,30,42,31,42,30,46,31,201,31,201,30,223,31,131,31,165,31,130,31,130,30,130,29,7,31,251,31,64,31,39,31,70,31,87,31,122,31,246,31,174,31,227,31,227,30,163,31,185,31,23,31,113,31,113,30,97,31,97,30,202,31,182,31,165,31,41,31,64,31,173,31,173,30,240,31,41,31,177,31,177,30,177,29,42,31,42,30,62,31,62,30,62,29,3,31,3,30,3,29,233,31,23,31,171,31,42,31,231,31,144,31,144,30,45,31,2,31,173,31,206,31,128,31,42,31,206,31,190,31,190,30,15,31,134,31,19,31,234,31,58,31,176,31,169,31,234,31,26,31,49,31,246,31,246,30,209,31,132,31,84,31,200,31,93,31,93,30,96,31,208,31,100,31,100,30,203,31,242,31,1,31,1,30,207,31,123,31,123,30,199,31,42,31,29,31,179,31,140,31,201,31,222,31,222,30,222,29,146,31,210,31,176,31,253,31,96,31,114,31,218,31,247,31,173,31,69,31,156,31,2,31,185,31,134,31,230,31,229,31,209,31,129,31,129,30,3,31,70,31,211,31,202,31,202,30,40,31,225,31,58,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
