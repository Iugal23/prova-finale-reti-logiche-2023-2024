-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_346 is
end project_tb_346;

architecture project_tb_arch_346 of project_tb_346 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 471;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (122,0,0,0,175,0,25,0,67,0,222,0,0,0,0,0,0,0,0,0,0,0,19,0,84,0,71,0,170,0,32,0,0,0,141,0,0,0,95,0,64,0,206,0,117,0,0,0,181,0,221,0,82,0,36,0,119,0,234,0,0,0,0,0,21,0,133,0,36,0,149,0,56,0,198,0,63,0,101,0,98,0,71,0,164,0,129,0,223,0,69,0,80,0,23,0,0,0,0,0,102,0,231,0,0,0,40,0,183,0,0,0,0,0,157,0,7,0,174,0,245,0,107,0,191,0,208,0,73,0,32,0,74,0,0,0,184,0,86,0,233,0,227,0,88,0,248,0,153,0,0,0,52,0,106,0,146,0,58,0,9,0,92,0,16,0,19,0,109,0,166,0,200,0,136,0,0,0,215,0,145,0,12,0,140,0,238,0,55,0,80,0,142,0,188,0,147,0,0,0,27,0,109,0,28,0,0,0,0,0,198,0,3,0,253,0,0,0,206,0,255,0,25,0,55,0,77,0,0,0,12,0,191,0,89,0,119,0,11,0,244,0,137,0,129,0,179,0,146,0,152,0,75,0,147,0,34,0,76,0,160,0,1,0,159,0,11,0,222,0,0,0,216,0,79,0,114,0,96,0,101,0,0,0,253,0,209,0,0,0,146,0,114,0,129,0,53,0,14,0,98,0,5,0,156,0,97,0,0,0,158,0,133,0,171,0,0,0,107,0,171,0,0,0,0,0,237,0,106,0,188,0,73,0,225,0,0,0,73,0,42,0,236,0,0,0,0,0,121,0,21,0,248,0,0,0,203,0,5,0,0,0,214,0,23,0,149,0,0,0,77,0,87,0,76,0,0,0,186,0,197,0,204,0,0,0,79,0,97,0,41,0,189,0,238,0,45,0,186,0,224,0,46,0,138,0,53,0,214,0,101,0,172,0,78,0,179,0,12,0,45,0,145,0,0,0,242,0,126,0,205,0,17,0,149,0,163,0,49,0,173,0,36,0,75,0,227,0,168,0,0,0,230,0,22,0,90,0,0,0,176,0,197,0,94,0,250,0,131,0,149,0,75,0,0,0,0,0,0,0,185,0,0,0,0,0,0,0,209,0,189,0,34,0,16,0,61,0,231,0,15,0,58,0,112,0,0,0,224,0,251,0,242,0,211,0,38,0,1,0,10,0,0,0,190,0,240,0,79,0,182,0,0,0,113,0,129,0,60,0,158,0,251,0,0,0,188,0,99,0,161,0,64,0,204,0,123,0,249,0,151,0,197,0,222,0,171,0,171,0,216,0,4,0,193,0,48,0,252,0,63,0,162,0,156,0,40,0,222,0,165,0,26,0,90,0,104,0,88,0,91,0,182,0,83,0,33,0,135,0,250,0,231,0,13,0,0,0,37,0,31,0,0,0,25,0,254,0,0,0,212,0,181,0,0,0,0,0,186,0,147,0,94,0,122,0,121,0,27,0,119,0,107,0,77,0,49,0,138,0,15,0,52,0,87,0,132,0,134,0,85,0,174,0,81,0,75,0,206,0,68,0,0,0,95,0,163,0,134,0,0,0,206,0,191,0,0,0,24,0,203,0,0,0,224,0,121,0,0,0,0,0,47,0,67,0,173,0,251,0,186,0,239,0,159,0,202,0,69,0,222,0,70,0,149,0,162,0,245,0,0,0,175,0,30,0,217,0,14,0,220,0,68,0,0,0,118,0,0,0,0,0,0,0,0,0,186,0,55,0,0,0,91,0,86,0,237,0,42,0,163,0,90,0,225,0,0,0,216,0,218,0,0,0,111,0,163,0,13,0,0,0,200,0,94,0,200,0,0,0,107,0,0,0,154,0,0,0,111,0,208,0,60,0,0,0,6,0,0,0,119,0,110,0,191,0,178,0,254,0,225,0,81,0,129,0,206,0,51,0,119,0,155,0,121,0,97,0,127,0,40,0,218,0,0,0,41,0,243,0,134,0,164,0,99,0,0,0,0,0,30,0,0,0,0,0,0,0,224,0,246,0,107,0,164,0,27,0,17,0,228,0,246,0,54,0,0,0,194,0,236,0,0,0,226,0,130,0,175,0,0,0,39,0,206,0,30,0,121,0,0,0,60,0,202,0,166,0,3,0,105,0);
signal scenario_full  : scenario_type := (122,31,122,30,175,31,25,31,67,31,222,31,222,30,222,29,222,28,222,27,222,26,19,31,84,31,71,31,170,31,32,31,32,30,141,31,141,30,95,31,64,31,206,31,117,31,117,30,181,31,221,31,82,31,36,31,119,31,234,31,234,30,234,29,21,31,133,31,36,31,149,31,56,31,198,31,63,31,101,31,98,31,71,31,164,31,129,31,223,31,69,31,80,31,23,31,23,30,23,29,102,31,231,31,231,30,40,31,183,31,183,30,183,29,157,31,7,31,174,31,245,31,107,31,191,31,208,31,73,31,32,31,74,31,74,30,184,31,86,31,233,31,227,31,88,31,248,31,153,31,153,30,52,31,106,31,146,31,58,31,9,31,92,31,16,31,19,31,109,31,166,31,200,31,136,31,136,30,215,31,145,31,12,31,140,31,238,31,55,31,80,31,142,31,188,31,147,31,147,30,27,31,109,31,28,31,28,30,28,29,198,31,3,31,253,31,253,30,206,31,255,31,25,31,55,31,77,31,77,30,12,31,191,31,89,31,119,31,11,31,244,31,137,31,129,31,179,31,146,31,152,31,75,31,147,31,34,31,76,31,160,31,1,31,159,31,11,31,222,31,222,30,216,31,79,31,114,31,96,31,101,31,101,30,253,31,209,31,209,30,146,31,114,31,129,31,53,31,14,31,98,31,5,31,156,31,97,31,97,30,158,31,133,31,171,31,171,30,107,31,171,31,171,30,171,29,237,31,106,31,188,31,73,31,225,31,225,30,73,31,42,31,236,31,236,30,236,29,121,31,21,31,248,31,248,30,203,31,5,31,5,30,214,31,23,31,149,31,149,30,77,31,87,31,76,31,76,30,186,31,197,31,204,31,204,30,79,31,97,31,41,31,189,31,238,31,45,31,186,31,224,31,46,31,138,31,53,31,214,31,101,31,172,31,78,31,179,31,12,31,45,31,145,31,145,30,242,31,126,31,205,31,17,31,149,31,163,31,49,31,173,31,36,31,75,31,227,31,168,31,168,30,230,31,22,31,90,31,90,30,176,31,197,31,94,31,250,31,131,31,149,31,75,31,75,30,75,29,75,28,185,31,185,30,185,29,185,28,209,31,189,31,34,31,16,31,61,31,231,31,15,31,58,31,112,31,112,30,224,31,251,31,242,31,211,31,38,31,1,31,10,31,10,30,190,31,240,31,79,31,182,31,182,30,113,31,129,31,60,31,158,31,251,31,251,30,188,31,99,31,161,31,64,31,204,31,123,31,249,31,151,31,197,31,222,31,171,31,171,31,216,31,4,31,193,31,48,31,252,31,63,31,162,31,156,31,40,31,222,31,165,31,26,31,90,31,104,31,88,31,91,31,182,31,83,31,33,31,135,31,250,31,231,31,13,31,13,30,37,31,31,31,31,30,25,31,254,31,254,30,212,31,181,31,181,30,181,29,186,31,147,31,94,31,122,31,121,31,27,31,119,31,107,31,77,31,49,31,138,31,15,31,52,31,87,31,132,31,134,31,85,31,174,31,81,31,75,31,206,31,68,31,68,30,95,31,163,31,134,31,134,30,206,31,191,31,191,30,24,31,203,31,203,30,224,31,121,31,121,30,121,29,47,31,67,31,173,31,251,31,186,31,239,31,159,31,202,31,69,31,222,31,70,31,149,31,162,31,245,31,245,30,175,31,30,31,217,31,14,31,220,31,68,31,68,30,118,31,118,30,118,29,118,28,118,27,186,31,55,31,55,30,91,31,86,31,237,31,42,31,163,31,90,31,225,31,225,30,216,31,218,31,218,30,111,31,163,31,13,31,13,30,200,31,94,31,200,31,200,30,107,31,107,30,154,31,154,30,111,31,208,31,60,31,60,30,6,31,6,30,119,31,110,31,191,31,178,31,254,31,225,31,81,31,129,31,206,31,51,31,119,31,155,31,121,31,97,31,127,31,40,31,218,31,218,30,41,31,243,31,134,31,164,31,99,31,99,30,99,29,30,31,30,30,30,29,30,28,224,31,246,31,107,31,164,31,27,31,17,31,228,31,246,31,54,31,54,30,194,31,236,31,236,30,226,31,130,31,175,31,175,30,39,31,206,31,30,31,121,31,121,30,60,31,202,31,166,31,3,31,105,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
