-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 933;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (245,0,79,0,0,0,119,0,46,0,69,0,251,0,0,0,196,0,0,0,91,0,96,0,0,0,164,0,4,0,173,0,244,0,114,0,112,0,0,0,0,0,0,0,38,0,186,0,247,0,0,0,162,0,160,0,92,0,0,0,228,0,0,0,143,0,91,0,232,0,123,0,140,0,0,0,240,0,144,0,0,0,232,0,171,0,92,0,2,0,234,0,219,0,188,0,143,0,157,0,191,0,0,0,250,0,0,0,204,0,95,0,0,0,0,0,59,0,12,0,179,0,249,0,0,0,63,0,38,0,92,0,194,0,127,0,139,0,225,0,0,0,247,0,171,0,145,0,147,0,159,0,144,0,122,0,32,0,41,0,47,0,41,0,232,0,121,0,169,0,56,0,226,0,123,0,207,0,99,0,228,0,0,0,156,0,0,0,164,0,198,0,244,0,233,0,178,0,0,0,0,0,116,0,77,0,38,0,203,0,0,0,195,0,6,0,73,0,0,0,222,0,196,0,0,0,216,0,86,0,18,0,116,0,134,0,161,0,228,0,0,0,29,0,23,0,223,0,12,0,83,0,0,0,241,0,0,0,75,0,25,0,124,0,28,0,232,0,52,0,34,0,0,0,0,0,56,0,209,0,0,0,244,0,213,0,121,0,255,0,129,0,3,0,0,0,237,0,120,0,47,0,141,0,181,0,251,0,126,0,0,0,103,0,0,0,127,0,159,0,158,0,94,0,130,0,45,0,62,0,0,0,0,0,24,0,151,0,249,0,182,0,142,0,63,0,98,0,27,0,20,0,104,0,155,0,65,0,154,0,197,0,251,0,185,0,196,0,163,0,0,0,0,0,178,0,0,0,235,0,0,0,34,0,58,0,255,0,100,0,0,0,6,0,193,0,0,0,19,0,125,0,55,0,105,0,240,0,119,0,76,0,0,0,129,0,21,0,0,0,184,0,171,0,181,0,0,0,115,0,64,0,117,0,212,0,159,0,248,0,197,0,208,0,158,0,192,0,161,0,106,0,222,0,249,0,198,0,135,0,163,0,140,0,57,0,150,0,239,0,172,0,159,0,247,0,0,0,235,0,148,0,234,0,236,0,42,0,212,0,220,0,19,0,0,0,156,0,177,0,90,0,212,0,0,0,41,0,171,0,85,0,205,0,233,0,149,0,0,0,58,0,117,0,52,0,108,0,49,0,65,0,0,0,133,0,147,0,143,0,202,0,0,0,0,0,59,0,27,0,0,0,27,0,117,0,192,0,230,0,45,0,36,0,0,0,0,0,119,0,0,0,9,0,101,0,35,0,0,0,203,0,200,0,0,0,159,0,98,0,233,0,0,0,51,0,34,0,213,0,141,0,0,0,200,0,85,0,64,0,0,0,88,0,98,0,7,0,37,0,15,0,150,0,205,0,110,0,0,0,250,0,0,0,11,0,2,0,0,0,190,0,97,0,245,0,245,0,136,0,246,0,150,0,73,0,0,0,155,0,254,0,221,0,71,0,60,0,47,0,0,0,173,0,115,0,28,0,52,0,252,0,184,0,176,0,105,0,2,0,104,0,242,0,74,0,81,0,190,0,0,0,112,0,17,0,228,0,18,0,11,0,52,0,222,0,172,0,0,0,69,0,36,0,163,0,8,0,64,0,0,0,242,0,14,0,30,0,168,0,26,0,252,0,0,0,34,0,144,0,31,0,114,0,226,0,44,0,41,0,249,0,215,0,111,0,101,0,192,0,7,0,0,0,155,0,255,0,229,0,0,0,0,0,0,0,55,0,183,0,45,0,0,0,231,0,203,0,244,0,206,0,0,0,233,0,124,0,84,0,214,0,32,0,60,0,174,0,139,0,139,0,8,0,9,0,77,0,143,0,132,0,172,0,130,0,196,0,130,0,68,0,148,0,97,0,214,0,55,0,152,0,0,0,93,0,243,0,172,0,165,0,0,0,0,0,192,0,177,0,0,0,0,0,222,0,96,0,126,0,8,0,115,0,166,0,0,0,219,0,28,0,41,0,38,0,59,0,202,0,42,0,134,0,199,0,0,0,230,0,17,0,0,0,149,0,56,0,174,0,0,0,204,0,151,0,62,0,195,0,201,0,48,0,124,0,52,0,110,0,144,0,52,0,24,0,0,0,75,0,230,0,0,0,95,0,143,0,243,0,0,0,0,0,90,0,176,0,93,0,223,0,217,0,11,0,31,0,56,0,164,0,13,0,50,0,104,0,0,0,194,0,83,0,37,0,233,0,115,0,138,0,196,0,99,0,195,0,113,0,89,0,124,0,0,0,103,0,0,0,224,0,13,0,235,0,103,0,0,0,235,0,151,0,200,0,198,0,143,0,0,0,0,0,82,0,0,0,140,0,242,0,88,0,66,0,224,0,0,0,140,0,134,0,228,0,48,0,171,0,100,0,232,0,0,0,43,0,5,0,0,0,0,0,0,0,0,0,140,0,82,0,40,0,197,0,131,0,67,0,41,0,132,0,192,0,233,0,217,0,0,0,0,0,180,0,58,0,0,0,133,0,46,0,166,0,253,0,66,0,27,0,58,0,68,0,230,0,0,0,140,0,227,0,22,0,108,0,193,0,0,0,55,0,47,0,162,0,52,0,127,0,0,0,0,0,84,0,0,0,120,0,4,0,21,0,243,0,17,0,151,0,97,0,24,0,244,0,46,0,23,0,68,0,112,0,192,0,76,0,161,0,178,0,25,0,204,0,125,0,55,0,153,0,0,0,0,0,88,0,137,0,187,0,76,0,16,0,58,0,139,0,0,0,154,0,138,0,0,0,0,0,0,0,0,0,120,0,149,0,0,0,152,0,230,0,149,0,69,0,54,0,187,0,72,0,0,0,0,0,153,0,124,0,0,0,0,0,24,0,0,0,238,0,0,0,0,0,147,0,116,0,247,0,170,0,54,0,0,0,154,0,24,0,0,0,250,0,144,0,0,0,0,0,58,0,58,0,10,0,157,0,0,0,225,0,223,0,138,0,0,0,0,0,16,0,97,0,95,0,213,0,0,0,153,0,18,0,145,0,0,0,82,0,2,0,161,0,108,0,51,0,144,0,182,0,201,0,0,0,205,0,73,0,44,0,184,0,142,0,0,0,107,0,119,0,234,0,100,0,89,0,199,0,19,0,225,0,87,0,145,0,3,0,0,0,170,0,44,0,88,0,2,0,160,0,197,0,208,0,7,0,0,0,0,0,161,0,26,0,56,0,240,0,235,0,0,0,47,0,175,0,235,0,142,0,150,0,0,0,208,0,88,0,0,0,141,0,249,0,247,0,162,0,11,0,0,0,167,0,179,0,0,0,196,0,107,0,0,0,76,0,19,0,230,0,176,0,47,0,218,0,0,0,0,0,0,0,154,0,0,0,93,0,0,0,119,0,219,0,0,0,12,0,184,0,228,0,88,0,47,0,0,0,165,0,0,0,243,0,42,0,238,0,95,0,0,0,110,0,69,0,185,0,0,0,217,0,71,0,177,0,12,0,97,0,0,0,124,0,11,0,199,0,121,0,112,0,76,0,0,0,101,0,189,0,0,0,242,0,139,0,202,0,155,0,170,0,0,0,38,0,0,0,0,0,45,0,20,0,56,0,20,0,217,0,0,0,156,0,41,0,228,0,155,0,36,0,77,0,209,0,76,0,0,0,0,0,186,0,107,0,73,0,237,0,233,0,10,0,0,0,26,0,235,0,183,0,95,0,176,0,108,0,133,0,12,0,75,0,38,0,0,0,15,0,0,0,0,0,217,0,112,0,45,0,0,0,63,0,0,0,227,0,152,0,233,0,81,0,149,0,74,0,0,0,99,0,96,0,181,0,118,0,37,0,26,0,209,0,0,0,77,0,65,0,0,0,207,0,25,0,244,0,156,0,54,0,186,0,170,0,0,0,0,0,52,0,138,0,2,0,0,0,233,0,244,0,0,0,176,0,122,0,0,0,224,0,102,0,0,0,93,0,95,0,52,0,109,0,5,0,0,0,38,0,119,0,199,0,248,0,45,0,169,0,254,0,116,0,250,0,0,0,41,0,181,0,241,0,0,0,103,0,162,0,254,0,122,0,169,0,59,0,4,0,121,0,43,0,32,0,62,0,0,0,247,0,223,0,98,0,88,0,0,0,81,0,116,0,193,0,217,0,0,0,115,0,35,0,0,0,142,0,233,0,232,0,89,0,52,0,68,0,252,0);
signal scenario_full  : scenario_type := (245,31,79,31,79,30,119,31,46,31,69,31,251,31,251,30,196,31,196,30,91,31,96,31,96,30,164,31,4,31,173,31,244,31,114,31,112,31,112,30,112,29,112,28,38,31,186,31,247,31,247,30,162,31,160,31,92,31,92,30,228,31,228,30,143,31,91,31,232,31,123,31,140,31,140,30,240,31,144,31,144,30,232,31,171,31,92,31,2,31,234,31,219,31,188,31,143,31,157,31,191,31,191,30,250,31,250,30,204,31,95,31,95,30,95,29,59,31,12,31,179,31,249,31,249,30,63,31,38,31,92,31,194,31,127,31,139,31,225,31,225,30,247,31,171,31,145,31,147,31,159,31,144,31,122,31,32,31,41,31,47,31,41,31,232,31,121,31,169,31,56,31,226,31,123,31,207,31,99,31,228,31,228,30,156,31,156,30,164,31,198,31,244,31,233,31,178,31,178,30,178,29,116,31,77,31,38,31,203,31,203,30,195,31,6,31,73,31,73,30,222,31,196,31,196,30,216,31,86,31,18,31,116,31,134,31,161,31,228,31,228,30,29,31,23,31,223,31,12,31,83,31,83,30,241,31,241,30,75,31,25,31,124,31,28,31,232,31,52,31,34,31,34,30,34,29,56,31,209,31,209,30,244,31,213,31,121,31,255,31,129,31,3,31,3,30,237,31,120,31,47,31,141,31,181,31,251,31,126,31,126,30,103,31,103,30,127,31,159,31,158,31,94,31,130,31,45,31,62,31,62,30,62,29,24,31,151,31,249,31,182,31,142,31,63,31,98,31,27,31,20,31,104,31,155,31,65,31,154,31,197,31,251,31,185,31,196,31,163,31,163,30,163,29,178,31,178,30,235,31,235,30,34,31,58,31,255,31,100,31,100,30,6,31,193,31,193,30,19,31,125,31,55,31,105,31,240,31,119,31,76,31,76,30,129,31,21,31,21,30,184,31,171,31,181,31,181,30,115,31,64,31,117,31,212,31,159,31,248,31,197,31,208,31,158,31,192,31,161,31,106,31,222,31,249,31,198,31,135,31,163,31,140,31,57,31,150,31,239,31,172,31,159,31,247,31,247,30,235,31,148,31,234,31,236,31,42,31,212,31,220,31,19,31,19,30,156,31,177,31,90,31,212,31,212,30,41,31,171,31,85,31,205,31,233,31,149,31,149,30,58,31,117,31,52,31,108,31,49,31,65,31,65,30,133,31,147,31,143,31,202,31,202,30,202,29,59,31,27,31,27,30,27,31,117,31,192,31,230,31,45,31,36,31,36,30,36,29,119,31,119,30,9,31,101,31,35,31,35,30,203,31,200,31,200,30,159,31,98,31,233,31,233,30,51,31,34,31,213,31,141,31,141,30,200,31,85,31,64,31,64,30,88,31,98,31,7,31,37,31,15,31,150,31,205,31,110,31,110,30,250,31,250,30,11,31,2,31,2,30,190,31,97,31,245,31,245,31,136,31,246,31,150,31,73,31,73,30,155,31,254,31,221,31,71,31,60,31,47,31,47,30,173,31,115,31,28,31,52,31,252,31,184,31,176,31,105,31,2,31,104,31,242,31,74,31,81,31,190,31,190,30,112,31,17,31,228,31,18,31,11,31,52,31,222,31,172,31,172,30,69,31,36,31,163,31,8,31,64,31,64,30,242,31,14,31,30,31,168,31,26,31,252,31,252,30,34,31,144,31,31,31,114,31,226,31,44,31,41,31,249,31,215,31,111,31,101,31,192,31,7,31,7,30,155,31,255,31,229,31,229,30,229,29,229,28,55,31,183,31,45,31,45,30,231,31,203,31,244,31,206,31,206,30,233,31,124,31,84,31,214,31,32,31,60,31,174,31,139,31,139,31,8,31,9,31,77,31,143,31,132,31,172,31,130,31,196,31,130,31,68,31,148,31,97,31,214,31,55,31,152,31,152,30,93,31,243,31,172,31,165,31,165,30,165,29,192,31,177,31,177,30,177,29,222,31,96,31,126,31,8,31,115,31,166,31,166,30,219,31,28,31,41,31,38,31,59,31,202,31,42,31,134,31,199,31,199,30,230,31,17,31,17,30,149,31,56,31,174,31,174,30,204,31,151,31,62,31,195,31,201,31,48,31,124,31,52,31,110,31,144,31,52,31,24,31,24,30,75,31,230,31,230,30,95,31,143,31,243,31,243,30,243,29,90,31,176,31,93,31,223,31,217,31,11,31,31,31,56,31,164,31,13,31,50,31,104,31,104,30,194,31,83,31,37,31,233,31,115,31,138,31,196,31,99,31,195,31,113,31,89,31,124,31,124,30,103,31,103,30,224,31,13,31,235,31,103,31,103,30,235,31,151,31,200,31,198,31,143,31,143,30,143,29,82,31,82,30,140,31,242,31,88,31,66,31,224,31,224,30,140,31,134,31,228,31,48,31,171,31,100,31,232,31,232,30,43,31,5,31,5,30,5,29,5,28,5,27,140,31,82,31,40,31,197,31,131,31,67,31,41,31,132,31,192,31,233,31,217,31,217,30,217,29,180,31,58,31,58,30,133,31,46,31,166,31,253,31,66,31,27,31,58,31,68,31,230,31,230,30,140,31,227,31,22,31,108,31,193,31,193,30,55,31,47,31,162,31,52,31,127,31,127,30,127,29,84,31,84,30,120,31,4,31,21,31,243,31,17,31,151,31,97,31,24,31,244,31,46,31,23,31,68,31,112,31,192,31,76,31,161,31,178,31,25,31,204,31,125,31,55,31,153,31,153,30,153,29,88,31,137,31,187,31,76,31,16,31,58,31,139,31,139,30,154,31,138,31,138,30,138,29,138,28,138,27,120,31,149,31,149,30,152,31,230,31,149,31,69,31,54,31,187,31,72,31,72,30,72,29,153,31,124,31,124,30,124,29,24,31,24,30,238,31,238,30,238,29,147,31,116,31,247,31,170,31,54,31,54,30,154,31,24,31,24,30,250,31,144,31,144,30,144,29,58,31,58,31,10,31,157,31,157,30,225,31,223,31,138,31,138,30,138,29,16,31,97,31,95,31,213,31,213,30,153,31,18,31,145,31,145,30,82,31,2,31,161,31,108,31,51,31,144,31,182,31,201,31,201,30,205,31,73,31,44,31,184,31,142,31,142,30,107,31,119,31,234,31,100,31,89,31,199,31,19,31,225,31,87,31,145,31,3,31,3,30,170,31,44,31,88,31,2,31,160,31,197,31,208,31,7,31,7,30,7,29,161,31,26,31,56,31,240,31,235,31,235,30,47,31,175,31,235,31,142,31,150,31,150,30,208,31,88,31,88,30,141,31,249,31,247,31,162,31,11,31,11,30,167,31,179,31,179,30,196,31,107,31,107,30,76,31,19,31,230,31,176,31,47,31,218,31,218,30,218,29,218,28,154,31,154,30,93,31,93,30,119,31,219,31,219,30,12,31,184,31,228,31,88,31,47,31,47,30,165,31,165,30,243,31,42,31,238,31,95,31,95,30,110,31,69,31,185,31,185,30,217,31,71,31,177,31,12,31,97,31,97,30,124,31,11,31,199,31,121,31,112,31,76,31,76,30,101,31,189,31,189,30,242,31,139,31,202,31,155,31,170,31,170,30,38,31,38,30,38,29,45,31,20,31,56,31,20,31,217,31,217,30,156,31,41,31,228,31,155,31,36,31,77,31,209,31,76,31,76,30,76,29,186,31,107,31,73,31,237,31,233,31,10,31,10,30,26,31,235,31,183,31,95,31,176,31,108,31,133,31,12,31,75,31,38,31,38,30,15,31,15,30,15,29,217,31,112,31,45,31,45,30,63,31,63,30,227,31,152,31,233,31,81,31,149,31,74,31,74,30,99,31,96,31,181,31,118,31,37,31,26,31,209,31,209,30,77,31,65,31,65,30,207,31,25,31,244,31,156,31,54,31,186,31,170,31,170,30,170,29,52,31,138,31,2,31,2,30,233,31,244,31,244,30,176,31,122,31,122,30,224,31,102,31,102,30,93,31,95,31,52,31,109,31,5,31,5,30,38,31,119,31,199,31,248,31,45,31,169,31,254,31,116,31,250,31,250,30,41,31,181,31,241,31,241,30,103,31,162,31,254,31,122,31,169,31,59,31,4,31,121,31,43,31,32,31,62,31,62,30,247,31,223,31,98,31,88,31,88,30,81,31,116,31,193,31,217,31,217,30,115,31,35,31,35,30,142,31,233,31,232,31,89,31,52,31,68,31,252,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
