-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 725;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (223,0,57,0,108,0,170,0,114,0,52,0,75,0,187,0,1,0,19,0,12,0,210,0,0,0,0,0,125,0,13,0,104,0,12,0,30,0,7,0,253,0,102,0,24,0,168,0,122,0,129,0,38,0,0,0,0,0,0,0,153,0,140,0,238,0,0,0,0,0,184,0,205,0,164,0,183,0,21,0,5,0,223,0,235,0,0,0,215,0,72,0,69,0,135,0,197,0,176,0,245,0,0,0,156,0,108,0,0,0,0,0,177,0,202,0,145,0,0,0,0,0,207,0,213,0,113,0,12,0,204,0,184,0,0,0,0,0,55,0,144,0,215,0,36,0,211,0,136,0,98,0,34,0,123,0,141,0,19,0,104,0,0,0,78,0,43,0,103,0,253,0,23,0,156,0,75,0,189,0,36,0,62,0,100,0,102,0,170,0,169,0,51,0,59,0,46,0,0,0,185,0,246,0,118,0,0,0,0,0,228,0,135,0,36,0,99,0,182,0,159,0,60,0,244,0,0,0,194,0,37,0,221,0,152,0,0,0,0,0,187,0,0,0,27,0,183,0,117,0,71,0,0,0,0,0,0,0,0,0,161,0,63,0,146,0,128,0,139,0,87,0,183,0,247,0,0,0,58,0,64,0,91,0,53,0,104,0,85,0,182,0,246,0,0,0,147,0,144,0,85,0,40,0,211,0,141,0,106,0,0,0,122,0,187,0,0,0,0,0,0,0,0,0,27,0,87,0,0,0,0,0,207,0,75,0,234,0,4,0,104,0,187,0,240,0,0,0,31,0,0,0,199,0,215,0,131,0,0,0,83,0,0,0,0,0,77,0,41,0,150,0,213,0,34,0,38,0,127,0,0,0,45,0,0,0,166,0,38,0,0,0,40,0,36,0,11,0,94,0,77,0,90,0,195,0,64,0,87,0,178,0,230,0,13,0,113,0,200,0,52,0,165,0,84,0,238,0,14,0,149,0,53,0,95,0,120,0,103,0,0,0,51,0,69,0,87,0,0,0,0,0,219,0,46,0,16,0,4,0,0,0,0,0,0,0,28,0,48,0,209,0,0,0,168,0,78,0,61,0,0,0,89,0,172,0,55,0,44,0,253,0,117,0,88,0,180,0,236,0,0,0,232,0,141,0,31,0,206,0,149,0,233,0,21,0,0,0,225,0,0,0,30,0,0,0,3,0,64,0,183,0,200,0,102,0,51,0,32,0,186,0,63,0,149,0,139,0,225,0,187,0,247,0,174,0,95,0,192,0,20,0,74,0,160,0,145,0,217,0,237,0,114,0,144,0,181,0,188,0,64,0,216,0,155,0,0,0,0,0,0,0,207,0,114,0,0,0,83,0,27,0,142,0,85,0,82,0,104,0,46,0,67,0,101,0,183,0,77,0,185,0,220,0,14,0,246,0,76,0,0,0,119,0,215,0,74,0,83,0,0,0,54,0,36,0,182,0,225,0,0,0,251,0,0,0,159,0,120,0,37,0,82,0,219,0,235,0,84,0,142,0,165,0,98,0,0,0,207,0,0,0,0,0,65,0,173,0,0,0,0,0,105,0,150,0,83,0,0,0,225,0,236,0,126,0,122,0,241,0,20,0,123,0,39,0,253,0,0,0,89,0,0,0,253,0,255,0,0,0,234,0,252,0,186,0,52,0,111,0,224,0,245,0,0,0,173,0,73,0,236,0,245,0,189,0,178,0,0,0,0,0,248,0,191,0,77,0,100,0,19,0,55,0,167,0,238,0,65,0,34,0,0,0,236,0,0,0,0,0,0,0,30,0,73,0,144,0,100,0,8,0,0,0,0,0,137,0,0,0,19,0,58,0,0,0,165,0,115,0,199,0,119,0,239,0,169,0,17,0,77,0,53,0,160,0,0,0,0,0,65,0,99,0,219,0,3,0,206,0,20,0,0,0,95,0,66,0,162,0,0,0,0,0,199,0,92,0,52,0,8,0,179,0,13,0,171,0,67,0,222,0,185,0,246,0,72,0,115,0,121,0,96,0,0,0,61,0,167,0,152,0,0,0,91,0,120,0,43,0,176,0,8,0,0,0,111,0,227,0,0,0,36,0,12,0,11,0,134,0,91,0,225,0,0,0,82,0,239,0,227,0,133,0,222,0,0,0,84,0,0,0,158,0,197,0,156,0,82,0,0,0,177,0,0,0,0,0,0,0,0,0,246,0,100,0,52,0,198,0,241,0,74,0,55,0,146,0,55,0,135,0,0,0,0,0,0,0,46,0,210,0,0,0,157,0,90,0,0,0,85,0,126,0,56,0,0,0,245,0,250,0,198,0,183,0,0,0,154,0,34,0,208,0,0,0,131,0,70,0,123,0,209,0,223,0,20,0,0,0,141,0,164,0,0,0,157,0,200,0,208,0,83,0,71,0,234,0,176,0,0,0,0,0,112,0,59,0,48,0,113,0,39,0,103,0,141,0,0,0,0,0,94,0,43,0,79,0,112,0,0,0,201,0,132,0,111,0,0,0,208,0,78,0,10,0,0,0,169,0,0,0,46,0,102,0,252,0,219,0,41,0,88,0,230,0,54,0,121,0,164,0,87,0,71,0,0,0,190,0,161,0,0,0,214,0,162,0,0,0,0,0,0,0,86,0,224,0,114,0,0,0,199,0,0,0,189,0,0,0,116,0,79,0,0,0,93,0,0,0,224,0,6,0,105,0,0,0,249,0,116,0,0,0,177,0,0,0,11,0,0,0,154,0,49,0,136,0,88,0,7,0,60,0,246,0,70,0,212,0,3,0,89,0,19,0,113,0,0,0,0,0,122,0,183,0,174,0,87,0,11,0,168,0,102,0,193,0,0,0,0,0,93,0,70,0,0,0,152,0,28,0,3,0,200,0,0,0,0,0,123,0,0,0,197,0,234,0,87,0,236,0,116,0,122,0,74,0,23,0,113,0,134,0,198,0,190,0,139,0,21,0,214,0,181,0,0,0,92,0,255,0,16,0,110,0,63,0,2,0,247,0,0,0,0,0,136,0,146,0,25,0,163,0,227,0,219,0,70,0,37,0,58,0,180,0,158,0,152,0,0,0,80,0,134,0,169,0,85,0,117,0,0,0,69,0,198,0,0,0,0,0,152,0,103,0,193,0,183,0,154,0,24,0,118,0,36,0,182,0,0,0,20,0,192,0,86,0,189,0,0,0,89,0,84,0,0,0,223,0,0,0,178,0,172,0,74,0,81,0,0,0,150,0,9,0,83,0,196,0,179,0,18,0,0,0,134,0,5,0);
signal scenario_full  : scenario_type := (223,31,57,31,108,31,170,31,114,31,52,31,75,31,187,31,1,31,19,31,12,31,210,31,210,30,210,29,125,31,13,31,104,31,12,31,30,31,7,31,253,31,102,31,24,31,168,31,122,31,129,31,38,31,38,30,38,29,38,28,153,31,140,31,238,31,238,30,238,29,184,31,205,31,164,31,183,31,21,31,5,31,223,31,235,31,235,30,215,31,72,31,69,31,135,31,197,31,176,31,245,31,245,30,156,31,108,31,108,30,108,29,177,31,202,31,145,31,145,30,145,29,207,31,213,31,113,31,12,31,204,31,184,31,184,30,184,29,55,31,144,31,215,31,36,31,211,31,136,31,98,31,34,31,123,31,141,31,19,31,104,31,104,30,78,31,43,31,103,31,253,31,23,31,156,31,75,31,189,31,36,31,62,31,100,31,102,31,170,31,169,31,51,31,59,31,46,31,46,30,185,31,246,31,118,31,118,30,118,29,228,31,135,31,36,31,99,31,182,31,159,31,60,31,244,31,244,30,194,31,37,31,221,31,152,31,152,30,152,29,187,31,187,30,27,31,183,31,117,31,71,31,71,30,71,29,71,28,71,27,161,31,63,31,146,31,128,31,139,31,87,31,183,31,247,31,247,30,58,31,64,31,91,31,53,31,104,31,85,31,182,31,246,31,246,30,147,31,144,31,85,31,40,31,211,31,141,31,106,31,106,30,122,31,187,31,187,30,187,29,187,28,187,27,27,31,87,31,87,30,87,29,207,31,75,31,234,31,4,31,104,31,187,31,240,31,240,30,31,31,31,30,199,31,215,31,131,31,131,30,83,31,83,30,83,29,77,31,41,31,150,31,213,31,34,31,38,31,127,31,127,30,45,31,45,30,166,31,38,31,38,30,40,31,36,31,11,31,94,31,77,31,90,31,195,31,64,31,87,31,178,31,230,31,13,31,113,31,200,31,52,31,165,31,84,31,238,31,14,31,149,31,53,31,95,31,120,31,103,31,103,30,51,31,69,31,87,31,87,30,87,29,219,31,46,31,16,31,4,31,4,30,4,29,4,28,28,31,48,31,209,31,209,30,168,31,78,31,61,31,61,30,89,31,172,31,55,31,44,31,253,31,117,31,88,31,180,31,236,31,236,30,232,31,141,31,31,31,206,31,149,31,233,31,21,31,21,30,225,31,225,30,30,31,30,30,3,31,64,31,183,31,200,31,102,31,51,31,32,31,186,31,63,31,149,31,139,31,225,31,187,31,247,31,174,31,95,31,192,31,20,31,74,31,160,31,145,31,217,31,237,31,114,31,144,31,181,31,188,31,64,31,216,31,155,31,155,30,155,29,155,28,207,31,114,31,114,30,83,31,27,31,142,31,85,31,82,31,104,31,46,31,67,31,101,31,183,31,77,31,185,31,220,31,14,31,246,31,76,31,76,30,119,31,215,31,74,31,83,31,83,30,54,31,36,31,182,31,225,31,225,30,251,31,251,30,159,31,120,31,37,31,82,31,219,31,235,31,84,31,142,31,165,31,98,31,98,30,207,31,207,30,207,29,65,31,173,31,173,30,173,29,105,31,150,31,83,31,83,30,225,31,236,31,126,31,122,31,241,31,20,31,123,31,39,31,253,31,253,30,89,31,89,30,253,31,255,31,255,30,234,31,252,31,186,31,52,31,111,31,224,31,245,31,245,30,173,31,73,31,236,31,245,31,189,31,178,31,178,30,178,29,248,31,191,31,77,31,100,31,19,31,55,31,167,31,238,31,65,31,34,31,34,30,236,31,236,30,236,29,236,28,30,31,73,31,144,31,100,31,8,31,8,30,8,29,137,31,137,30,19,31,58,31,58,30,165,31,115,31,199,31,119,31,239,31,169,31,17,31,77,31,53,31,160,31,160,30,160,29,65,31,99,31,219,31,3,31,206,31,20,31,20,30,95,31,66,31,162,31,162,30,162,29,199,31,92,31,52,31,8,31,179,31,13,31,171,31,67,31,222,31,185,31,246,31,72,31,115,31,121,31,96,31,96,30,61,31,167,31,152,31,152,30,91,31,120,31,43,31,176,31,8,31,8,30,111,31,227,31,227,30,36,31,12,31,11,31,134,31,91,31,225,31,225,30,82,31,239,31,227,31,133,31,222,31,222,30,84,31,84,30,158,31,197,31,156,31,82,31,82,30,177,31,177,30,177,29,177,28,177,27,246,31,100,31,52,31,198,31,241,31,74,31,55,31,146,31,55,31,135,31,135,30,135,29,135,28,46,31,210,31,210,30,157,31,90,31,90,30,85,31,126,31,56,31,56,30,245,31,250,31,198,31,183,31,183,30,154,31,34,31,208,31,208,30,131,31,70,31,123,31,209,31,223,31,20,31,20,30,141,31,164,31,164,30,157,31,200,31,208,31,83,31,71,31,234,31,176,31,176,30,176,29,112,31,59,31,48,31,113,31,39,31,103,31,141,31,141,30,141,29,94,31,43,31,79,31,112,31,112,30,201,31,132,31,111,31,111,30,208,31,78,31,10,31,10,30,169,31,169,30,46,31,102,31,252,31,219,31,41,31,88,31,230,31,54,31,121,31,164,31,87,31,71,31,71,30,190,31,161,31,161,30,214,31,162,31,162,30,162,29,162,28,86,31,224,31,114,31,114,30,199,31,199,30,189,31,189,30,116,31,79,31,79,30,93,31,93,30,224,31,6,31,105,31,105,30,249,31,116,31,116,30,177,31,177,30,11,31,11,30,154,31,49,31,136,31,88,31,7,31,60,31,246,31,70,31,212,31,3,31,89,31,19,31,113,31,113,30,113,29,122,31,183,31,174,31,87,31,11,31,168,31,102,31,193,31,193,30,193,29,93,31,70,31,70,30,152,31,28,31,3,31,200,31,200,30,200,29,123,31,123,30,197,31,234,31,87,31,236,31,116,31,122,31,74,31,23,31,113,31,134,31,198,31,190,31,139,31,21,31,214,31,181,31,181,30,92,31,255,31,16,31,110,31,63,31,2,31,247,31,247,30,247,29,136,31,146,31,25,31,163,31,227,31,219,31,70,31,37,31,58,31,180,31,158,31,152,31,152,30,80,31,134,31,169,31,85,31,117,31,117,30,69,31,198,31,198,30,198,29,152,31,103,31,193,31,183,31,154,31,24,31,118,31,36,31,182,31,182,30,20,31,192,31,86,31,189,31,189,30,89,31,84,31,84,30,223,31,223,30,178,31,172,31,74,31,81,31,81,30,150,31,9,31,83,31,196,31,179,31,18,31,18,30,134,31,5,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
