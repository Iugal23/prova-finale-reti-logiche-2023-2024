-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_270 is
end project_tb_270;

architecture project_tb_arch_270 of project_tb_270 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 276;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (122,0,107,0,17,0,212,0,6,0,80,0,27,0,133,0,241,0,0,0,112,0,171,0,157,0,224,0,33,0,241,0,0,0,0,0,92,0,108,0,145,0,251,0,204,0,56,0,30,0,0,0,0,0,104,0,47,0,9,0,0,0,252,0,135,0,17,0,0,0,22,0,0,0,148,0,206,0,73,0,207,0,0,0,94,0,0,0,121,0,122,0,137,0,177,0,157,0,0,0,167,0,182,0,159,0,5,0,193,0,0,0,113,0,108,0,155,0,0,0,29,0,215,0,0,0,208,0,218,0,0,0,233,0,250,0,74,0,178,0,0,0,0,0,0,0,145,0,0,0,0,0,239,0,240,0,254,0,84,0,0,0,217,0,130,0,255,0,37,0,160,0,86,0,173,0,109,0,91,0,0,0,130,0,174,0,125,0,251,0,255,0,28,0,39,0,101,0,125,0,0,0,110,0,146,0,237,0,53,0,0,0,46,0,213,0,50,0,46,0,185,0,0,0,76,0,48,0,114,0,107,0,136,0,226,0,15,0,0,0,154,0,189,0,246,0,88,0,204,0,250,0,194,0,0,0,237,0,187,0,61,0,212,0,54,0,0,0,104,0,0,0,149,0,76,0,146,0,122,0,151,0,232,0,211,0,67,0,231,0,146,0,0,0,158,0,117,0,0,0,42,0,96,0,162,0,27,0,0,0,224,0,114,0,104,0,174,0,216,0,223,0,0,0,63,0,170,0,236,0,0,0,0,0,183,0,0,0,250,0,196,0,0,0,127,0,210,0,106,0,82,0,162,0,20,0,241,0,0,0,9,0,219,0,93,0,135,0,170,0,45,0,102,0,225,0,8,0,50,0,182,0,65,0,0,0,161,0,233,0,0,0,0,0,129,0,101,0,179,0,0,0,36,0,29,0,0,0,0,0,0,0,140,0,64,0,241,0,207,0,166,0,254,0,134,0,119,0,103,0,242,0,0,0,0,0,98,0,4,0,239,0,147,0,160,0,45,0,90,0,243,0,55,0,0,0,42,0,182,0,84,0,0,0,230,0,80,0,226,0,51,0,101,0,129,0,116,0,131,0,95,0,73,0,248,0,60,0,159,0,0,0,0,0,0,0,246,0,0,0,26,0,125,0,0,0,110,0,243,0,128,0,227,0,76,0,238,0,132,0,128,0,243,0,83,0,0,0,15,0,34,0,0,0,17,0,81,0,218,0,50,0,25,0,22,0,130,0,19,0,23,0);
signal scenario_full  : scenario_type := (122,31,107,31,17,31,212,31,6,31,80,31,27,31,133,31,241,31,241,30,112,31,171,31,157,31,224,31,33,31,241,31,241,30,241,29,92,31,108,31,145,31,251,31,204,31,56,31,30,31,30,30,30,29,104,31,47,31,9,31,9,30,252,31,135,31,17,31,17,30,22,31,22,30,148,31,206,31,73,31,207,31,207,30,94,31,94,30,121,31,122,31,137,31,177,31,157,31,157,30,167,31,182,31,159,31,5,31,193,31,193,30,113,31,108,31,155,31,155,30,29,31,215,31,215,30,208,31,218,31,218,30,233,31,250,31,74,31,178,31,178,30,178,29,178,28,145,31,145,30,145,29,239,31,240,31,254,31,84,31,84,30,217,31,130,31,255,31,37,31,160,31,86,31,173,31,109,31,91,31,91,30,130,31,174,31,125,31,251,31,255,31,28,31,39,31,101,31,125,31,125,30,110,31,146,31,237,31,53,31,53,30,46,31,213,31,50,31,46,31,185,31,185,30,76,31,48,31,114,31,107,31,136,31,226,31,15,31,15,30,154,31,189,31,246,31,88,31,204,31,250,31,194,31,194,30,237,31,187,31,61,31,212,31,54,31,54,30,104,31,104,30,149,31,76,31,146,31,122,31,151,31,232,31,211,31,67,31,231,31,146,31,146,30,158,31,117,31,117,30,42,31,96,31,162,31,27,31,27,30,224,31,114,31,104,31,174,31,216,31,223,31,223,30,63,31,170,31,236,31,236,30,236,29,183,31,183,30,250,31,196,31,196,30,127,31,210,31,106,31,82,31,162,31,20,31,241,31,241,30,9,31,219,31,93,31,135,31,170,31,45,31,102,31,225,31,8,31,50,31,182,31,65,31,65,30,161,31,233,31,233,30,233,29,129,31,101,31,179,31,179,30,36,31,29,31,29,30,29,29,29,28,140,31,64,31,241,31,207,31,166,31,254,31,134,31,119,31,103,31,242,31,242,30,242,29,98,31,4,31,239,31,147,31,160,31,45,31,90,31,243,31,55,31,55,30,42,31,182,31,84,31,84,30,230,31,80,31,226,31,51,31,101,31,129,31,116,31,131,31,95,31,73,31,248,31,60,31,159,31,159,30,159,29,159,28,246,31,246,30,26,31,125,31,125,30,110,31,243,31,128,31,227,31,76,31,238,31,132,31,128,31,243,31,83,31,83,30,15,31,34,31,34,30,17,31,81,31,218,31,50,31,25,31,22,31,130,31,19,31,23,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
