-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 617;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (146,0,202,0,179,0,95,0,91,0,215,0,0,0,227,0,69,0,231,0,5,0,209,0,36,0,0,0,193,0,0,0,155,0,96,0,169,0,225,0,127,0,196,0,239,0,156,0,18,0,0,0,70,0,56,0,131,0,165,0,187,0,0,0,222,0,216,0,115,0,169,0,71,0,46,0,0,0,0,0,95,0,210,0,12,0,0,0,6,0,168,0,19,0,63,0,71,0,0,0,116,0,236,0,229,0,13,0,162,0,36,0,244,0,0,0,250,0,106,0,0,0,107,0,61,0,104,0,11,0,112,0,86,0,79,0,221,0,232,0,174,0,0,0,195,0,145,0,65,0,72,0,90,0,240,0,104,0,77,0,134,0,0,0,196,0,174,0,66,0,186,0,45,0,77,0,0,0,162,0,0,0,56,0,137,0,184,0,99,0,0,0,0,0,239,0,179,0,0,0,36,0,201,0,128,0,104,0,109,0,148,0,103,0,100,0,188,0,130,0,72,0,0,0,98,0,5,0,176,0,0,0,160,0,117,0,100,0,38,0,0,0,76,0,154,0,0,0,137,0,176,0,0,0,24,0,75,0,185,0,189,0,158,0,65,0,83,0,1,0,104,0,0,0,227,0,208,0,150,0,88,0,143,0,0,0,75,0,5,0,89,0,235,0,252,0,61,0,106,0,38,0,33,0,90,0,104,0,2,0,48,0,29,0,94,0,72,0,171,0,0,0,93,0,165,0,220,0,134,0,191,0,146,0,0,0,98,0,85,0,227,0,153,0,191,0,74,0,213,0,245,0,50,0,113,0,62,0,0,0,0,0,137,0,205,0,174,0,26,0,30,0,244,0,49,0,250,0,82,0,144,0,85,0,154,0,36,0,0,0,9,0,0,0,0,0,0,0,234,0,0,0,88,0,24,0,163,0,232,0,87,0,219,0,96,0,104,0,23,0,8,0,70,0,0,0,0,0,127,0,0,0,83,0,221,0,57,0,175,0,152,0,233,0,0,0,170,0,186,0,50,0,176,0,42,0,192,0,182,0,1,0,83,0,0,0,174,0,250,0,24,0,17,0,182,0,211,0,211,0,2,0,0,0,181,0,126,0,41,0,92,0,250,0,98,0,152,0,4,0,165,0,0,0,91,0,241,0,223,0,0,0,205,0,0,0,203,0,86,0,217,0,139,0,128,0,28,0,40,0,13,0,207,0,46,0,83,0,71,0,159,0,239,0,38,0,139,0,112,0,183,0,0,0,0,0,205,0,102,0,22,0,0,0,54,0,197,0,0,0,0,0,0,0,8,0,97,0,81,0,132,0,0,0,168,0,86,0,1,0,48,0,223,0,0,0,183,0,88,0,122,0,159,0,42,0,226,0,25,0,62,0,119,0,130,0,70,0,0,0,101,0,216,0,141,0,94,0,232,0,192,0,0,0,188,0,0,0,78,0,158,0,0,0,119,0,0,0,35,0,0,0,0,0,219,0,74,0,76,0,97,0,0,0,102,0,28,0,102,0,91,0,0,0,0,0,139,0,0,0,20,0,99,0,46,0,211,0,3,0,105,0,144,0,87,0,236,0,5,0,192,0,0,0,0,0,0,0,24,0,233,0,203,0,166,0,2,0,203,0,0,0,114,0,100,0,53,0,232,0,38,0,0,0,204,0,0,0,245,0,92,0,242,0,0,0,3,0,0,0,243,0,252,0,176,0,223,0,210,0,195,0,0,0,0,0,105,0,176,0,89,0,89,0,212,0,11,0,0,0,0,0,226,0,28,0,192,0,0,0,205,0,121,0,117,0,87,0,116,0,45,0,0,0,28,0,148,0,0,0,55,0,244,0,24,0,118,0,142,0,17,0,0,0,71,0,171,0,0,0,221,0,19,0,202,0,183,0,153,0,71,0,115,0,73,0,0,0,246,0,194,0,44,0,0,0,0,0,103,0,71,0,210,0,40,0,96,0,14,0,0,0,158,0,70,0,146,0,0,0,0,0,113,0,13,0,232,0,0,0,19,0,29,0,30,0,249,0,251,0,150,0,79,0,202,0,0,0,42,0,126,0,0,0,0,0,155,0,0,0,38,0,252,0,102,0,11,0,69,0,141,0,66,0,162,0,0,0,105,0,204,0,88,0,46,0,6,0,75,0,59,0,81,0,208,0,220,0,129,0,0,0,0,0,187,0,123,0,0,0,213,0,101,0,221,0,0,0,215,0,233,0,0,0,0,0,0,0,0,0,234,0,227,0,18,0,0,0,219,0,41,0,0,0,88,0,129,0,249,0,97,0,122,0,0,0,126,0,0,0,0,0,132,0,83,0,133,0,182,0,90,0,3,0,146,0,206,0,240,0,122,0,177,0,79,0,228,0,239,0,190,0,100,0,179,0,140,0,0,0,0,0,0,0,106,0,58,0,195,0,75,0,0,0,236,0,0,0,120,0,89,0,188,0,197,0,0,0,130,0,43,0,167,0,219,0,233,0,0,0,162,0,161,0,217,0,125,0,176,0,142,0,60,0,20,0,157,0,150,0,50,0,15,0,169,0,178,0,39,0,56,0,143,0,86,0,0,0,82,0,177,0,88,0,49,0,0,0,254,0,165,0,0,0,7,0,43,0,27,0,226,0,62,0,61,0,193,0,0,0,60,0,30,0,53,0,51,0,0,0,4,0,14,0,189,0,209,0,96,0,195,0,61,0,0,0,0,0,0,0,195,0,101,0,0,0,54,0,0,0,163,0,4,0,159,0,14,0,154,0,127,0,226,0,199,0,211,0,58,0,0,0,230,0);
signal scenario_full  : scenario_type := (146,31,202,31,179,31,95,31,91,31,215,31,215,30,227,31,69,31,231,31,5,31,209,31,36,31,36,30,193,31,193,30,155,31,96,31,169,31,225,31,127,31,196,31,239,31,156,31,18,31,18,30,70,31,56,31,131,31,165,31,187,31,187,30,222,31,216,31,115,31,169,31,71,31,46,31,46,30,46,29,95,31,210,31,12,31,12,30,6,31,168,31,19,31,63,31,71,31,71,30,116,31,236,31,229,31,13,31,162,31,36,31,244,31,244,30,250,31,106,31,106,30,107,31,61,31,104,31,11,31,112,31,86,31,79,31,221,31,232,31,174,31,174,30,195,31,145,31,65,31,72,31,90,31,240,31,104,31,77,31,134,31,134,30,196,31,174,31,66,31,186,31,45,31,77,31,77,30,162,31,162,30,56,31,137,31,184,31,99,31,99,30,99,29,239,31,179,31,179,30,36,31,201,31,128,31,104,31,109,31,148,31,103,31,100,31,188,31,130,31,72,31,72,30,98,31,5,31,176,31,176,30,160,31,117,31,100,31,38,31,38,30,76,31,154,31,154,30,137,31,176,31,176,30,24,31,75,31,185,31,189,31,158,31,65,31,83,31,1,31,104,31,104,30,227,31,208,31,150,31,88,31,143,31,143,30,75,31,5,31,89,31,235,31,252,31,61,31,106,31,38,31,33,31,90,31,104,31,2,31,48,31,29,31,94,31,72,31,171,31,171,30,93,31,165,31,220,31,134,31,191,31,146,31,146,30,98,31,85,31,227,31,153,31,191,31,74,31,213,31,245,31,50,31,113,31,62,31,62,30,62,29,137,31,205,31,174,31,26,31,30,31,244,31,49,31,250,31,82,31,144,31,85,31,154,31,36,31,36,30,9,31,9,30,9,29,9,28,234,31,234,30,88,31,24,31,163,31,232,31,87,31,219,31,96,31,104,31,23,31,8,31,70,31,70,30,70,29,127,31,127,30,83,31,221,31,57,31,175,31,152,31,233,31,233,30,170,31,186,31,50,31,176,31,42,31,192,31,182,31,1,31,83,31,83,30,174,31,250,31,24,31,17,31,182,31,211,31,211,31,2,31,2,30,181,31,126,31,41,31,92,31,250,31,98,31,152,31,4,31,165,31,165,30,91,31,241,31,223,31,223,30,205,31,205,30,203,31,86,31,217,31,139,31,128,31,28,31,40,31,13,31,207,31,46,31,83,31,71,31,159,31,239,31,38,31,139,31,112,31,183,31,183,30,183,29,205,31,102,31,22,31,22,30,54,31,197,31,197,30,197,29,197,28,8,31,97,31,81,31,132,31,132,30,168,31,86,31,1,31,48,31,223,31,223,30,183,31,88,31,122,31,159,31,42,31,226,31,25,31,62,31,119,31,130,31,70,31,70,30,101,31,216,31,141,31,94,31,232,31,192,31,192,30,188,31,188,30,78,31,158,31,158,30,119,31,119,30,35,31,35,30,35,29,219,31,74,31,76,31,97,31,97,30,102,31,28,31,102,31,91,31,91,30,91,29,139,31,139,30,20,31,99,31,46,31,211,31,3,31,105,31,144,31,87,31,236,31,5,31,192,31,192,30,192,29,192,28,24,31,233,31,203,31,166,31,2,31,203,31,203,30,114,31,100,31,53,31,232,31,38,31,38,30,204,31,204,30,245,31,92,31,242,31,242,30,3,31,3,30,243,31,252,31,176,31,223,31,210,31,195,31,195,30,195,29,105,31,176,31,89,31,89,31,212,31,11,31,11,30,11,29,226,31,28,31,192,31,192,30,205,31,121,31,117,31,87,31,116,31,45,31,45,30,28,31,148,31,148,30,55,31,244,31,24,31,118,31,142,31,17,31,17,30,71,31,171,31,171,30,221,31,19,31,202,31,183,31,153,31,71,31,115,31,73,31,73,30,246,31,194,31,44,31,44,30,44,29,103,31,71,31,210,31,40,31,96,31,14,31,14,30,158,31,70,31,146,31,146,30,146,29,113,31,13,31,232,31,232,30,19,31,29,31,30,31,249,31,251,31,150,31,79,31,202,31,202,30,42,31,126,31,126,30,126,29,155,31,155,30,38,31,252,31,102,31,11,31,69,31,141,31,66,31,162,31,162,30,105,31,204,31,88,31,46,31,6,31,75,31,59,31,81,31,208,31,220,31,129,31,129,30,129,29,187,31,123,31,123,30,213,31,101,31,221,31,221,30,215,31,233,31,233,30,233,29,233,28,233,27,234,31,227,31,18,31,18,30,219,31,41,31,41,30,88,31,129,31,249,31,97,31,122,31,122,30,126,31,126,30,126,29,132,31,83,31,133,31,182,31,90,31,3,31,146,31,206,31,240,31,122,31,177,31,79,31,228,31,239,31,190,31,100,31,179,31,140,31,140,30,140,29,140,28,106,31,58,31,195,31,75,31,75,30,236,31,236,30,120,31,89,31,188,31,197,31,197,30,130,31,43,31,167,31,219,31,233,31,233,30,162,31,161,31,217,31,125,31,176,31,142,31,60,31,20,31,157,31,150,31,50,31,15,31,169,31,178,31,39,31,56,31,143,31,86,31,86,30,82,31,177,31,88,31,49,31,49,30,254,31,165,31,165,30,7,31,43,31,27,31,226,31,62,31,61,31,193,31,193,30,60,31,30,31,53,31,51,31,51,30,4,31,14,31,189,31,209,31,96,31,195,31,61,31,61,30,61,29,61,28,195,31,101,31,101,30,54,31,54,30,163,31,4,31,159,31,14,31,154,31,127,31,226,31,199,31,211,31,58,31,58,30,230,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
