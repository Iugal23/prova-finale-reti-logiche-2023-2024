-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 696;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,54,0,0,0,125,0,0,0,0,0,0,0,0,0,0,0,216,0,0,0,132,0,199,0,0,0,221,0,50,0,250,0,1,0,0,0,98,0,166,0,34,0,100,0,37,0,203,0,220,0,9,0,54,0,135,0,217,0,242,0,0,0,108,0,178,0,0,0,227,0,77,0,238,0,0,0,251,0,0,0,102,0,230,0,54,0,184,0,34,0,137,0,102,0,124,0,232,0,75,0,0,0,190,0,232,0,34,0,204,0,129,0,0,0,247,0,228,0,61,0,45,0,86,0,253,0,208,0,97,0,114,0,0,0,0,0,70,0,0,0,165,0,176,0,227,0,68,0,69,0,248,0,0,0,228,0,0,0,183,0,0,0,120,0,0,0,216,0,137,0,213,0,70,0,231,0,132,0,0,0,0,0,98,0,196,0,0,0,59,0,173,0,238,0,0,0,210,0,201,0,92,0,0,0,175,0,0,0,0,0,209,0,238,0,102,0,146,0,70,0,100,0,0,0,235,0,0,0,0,0,23,0,221,0,164,0,79,0,134,0,140,0,252,0,119,0,169,0,233,0,4,0,0,0,118,0,132,0,121,0,230,0,0,0,18,0,16,0,0,0,16,0,225,0,97,0,142,0,244,0,0,0,218,0,0,0,218,0,85,0,209,0,254,0,0,0,92,0,207,0,0,0,221,0,7,0,0,0,35,0,241,0,0,0,96,0,83,0,3,0,0,0,184,0,195,0,24,0,123,0,33,0,146,0,0,0,191,0,0,0,0,0,3,0,203,0,145,0,211,0,39,0,1,0,104,0,101,0,0,0,0,0,0,0,177,0,0,0,42,0,22,0,234,0,132,0,21,0,49,0,201,0,227,0,153,0,25,0,0,0,170,0,0,0,0,0,196,0,96,0,70,0,195,0,99,0,0,0,61,0,4,0,48,0,78,0,60,0,217,0,0,0,24,0,0,0,212,0,238,0,0,0,126,0,218,0,143,0,217,0,56,0,0,0,120,0,0,0,139,0,103,0,0,0,162,0,50,0,55,0,219,0,254,0,119,0,44,0,0,0,107,0,0,0,0,0,117,0,212,0,0,0,221,0,240,0,249,0,229,0,238,0,217,0,48,0,0,0,155,0,245,0,122,0,219,0,25,0,52,0,245,0,82,0,83,0,0,0,0,0,241,0,245,0,79,0,65,0,20,0,54,0,201,0,207,0,26,0,0,0,0,0,32,0,88,0,158,0,13,0,2,0,35,0,174,0,0,0,246,0,0,0,66,0,109,0,0,0,0,0,143,0,147,0,95,0,3,0,183,0,146,0,110,0,137,0,170,0,156,0,212,0,114,0,153,0,187,0,136,0,163,0,152,0,18,0,24,0,63,0,246,0,211,0,45,0,194,0,94,0,221,0,89,0,29,0,45,0,125,0,173,0,0,0,218,0,156,0,55,0,117,0,180,0,63,0,47,0,255,0,0,0,234,0,119,0,251,0,64,0,161,0,241,0,7,0,0,0,41,0,148,0,255,0,161,0,0,0,0,0,70,0,120,0,244,0,0,0,218,0,191,0,246,0,63,0,186,0,0,0,121,0,140,0,0,0,158,0,130,0,109,0,118,0,213,0,129,0,0,0,127,0,45,0,206,0,38,0,212,0,236,0,192,0,0,0,71,0,0,0,52,0,128,0,176,0,224,0,230,0,76,0,242,0,203,0,9,0,242,0,132,0,245,0,222,0,196,0,16,0,40,0,111,0,242,0,164,0,134,0,0,0,48,0,25,0,0,0,184,0,31,0,215,0,199,0,46,0,87,0,7,0,0,0,40,0,187,0,23,0,173,0,13,0,216,0,44,0,161,0,161,0,51,0,15,0,28,0,0,0,204,0,0,0,171,0,0,0,131,0,23,0,237,0,207,0,11,0,197,0,0,0,79,0,22,0,130,0,84,0,195,0,238,0,123,0,56,0,221,0,10,0,127,0,154,0,173,0,236,0,128,0,0,0,182,0,47,0,242,0,0,0,167,0,178,0,41,0,217,0,121,0,68,0,176,0,211,0,25,0,159,0,76,0,0,0,68,0,0,0,178,0,17,0,18,0,71,0,159,0,1,0,0,0,0,0,0,0,184,0,0,0,224,0,186,0,0,0,186,0,0,0,0,0,154,0,229,0,222,0,159,0,223,0,253,0,59,0,32,0,159,0,152,0,77,0,0,0,242,0,0,0,98,0,20,0,59,0,0,0,88,0,50,0,29,0,206,0,112,0,245,0,209,0,48,0,237,0,176,0,155,0,95,0,1,0,159,0,70,0,222,0,147,0,74,0,104,0,169,0,181,0,126,0,144,0,159,0,29,0,41,0,0,0,214,0,116,0,0,0,0,0,160,0,10,0,46,0,13,0,147,0,74,0,241,0,173,0,79,0,147,0,61,0,77,0,0,0,235,0,118,0,36,0,0,0,0,0,0,0,109,0,135,0,0,0,30,0,31,0,117,0,230,0,0,0,172,0,0,0,245,0,42,0,61,0,239,0,0,0,0,0,76,0,28,0,233,0,105,0,117,0,0,0,0,0,184,0,0,0,41,0,177,0,106,0,136,0,127,0,0,0,126,0,103,0,74,0,42,0,201,0,0,0,0,0,178,0,0,0,16,0,0,0,0,0,0,0,66,0,237,0,39,0,21,0,23,0,34,0,0,0,188,0,51,0,0,0,188,0,170,0,168,0,71,0,0,0,107,0,90,0,0,0,30,0,141,0,115,0,29,0,111,0,93,0,201,0,0,0,0,0,25,0,0,0,53,0,175,0,34,0,84,0,223,0,85,0,22,0,0,0,75,0,0,0,91,0,78,0,253,0,71,0,137,0,100,0,251,0,72,0,154,0,230,0,214,0,206,0,0,0,238,0,210,0,0,0,168,0,58,0,162,0,10,0,0,0,111,0,237,0,232,0,156,0,150,0,34,0,61,0,114,0,108,0,0,0,140,0,37,0,78,0,146,0,36,0,148,0,63,0,195,0,23,0,27,0,185,0,0,0,152,0,0,0,143,0,0,0,230,0,26,0,162,0,129,0,231,0,165,0,0,0,0,0,114,0,206,0,167,0,95,0,86,0,0,0,142,0,0,0,0,0,199,0,72,0,246,0);
signal scenario_full  : scenario_type := (0,0,54,31,54,30,125,31,125,30,125,29,125,28,125,27,125,26,216,31,216,30,132,31,199,31,199,30,221,31,50,31,250,31,1,31,1,30,98,31,166,31,34,31,100,31,37,31,203,31,220,31,9,31,54,31,135,31,217,31,242,31,242,30,108,31,178,31,178,30,227,31,77,31,238,31,238,30,251,31,251,30,102,31,230,31,54,31,184,31,34,31,137,31,102,31,124,31,232,31,75,31,75,30,190,31,232,31,34,31,204,31,129,31,129,30,247,31,228,31,61,31,45,31,86,31,253,31,208,31,97,31,114,31,114,30,114,29,70,31,70,30,165,31,176,31,227,31,68,31,69,31,248,31,248,30,228,31,228,30,183,31,183,30,120,31,120,30,216,31,137,31,213,31,70,31,231,31,132,31,132,30,132,29,98,31,196,31,196,30,59,31,173,31,238,31,238,30,210,31,201,31,92,31,92,30,175,31,175,30,175,29,209,31,238,31,102,31,146,31,70,31,100,31,100,30,235,31,235,30,235,29,23,31,221,31,164,31,79,31,134,31,140,31,252,31,119,31,169,31,233,31,4,31,4,30,118,31,132,31,121,31,230,31,230,30,18,31,16,31,16,30,16,31,225,31,97,31,142,31,244,31,244,30,218,31,218,30,218,31,85,31,209,31,254,31,254,30,92,31,207,31,207,30,221,31,7,31,7,30,35,31,241,31,241,30,96,31,83,31,3,31,3,30,184,31,195,31,24,31,123,31,33,31,146,31,146,30,191,31,191,30,191,29,3,31,203,31,145,31,211,31,39,31,1,31,104,31,101,31,101,30,101,29,101,28,177,31,177,30,42,31,22,31,234,31,132,31,21,31,49,31,201,31,227,31,153,31,25,31,25,30,170,31,170,30,170,29,196,31,96,31,70,31,195,31,99,31,99,30,61,31,4,31,48,31,78,31,60,31,217,31,217,30,24,31,24,30,212,31,238,31,238,30,126,31,218,31,143,31,217,31,56,31,56,30,120,31,120,30,139,31,103,31,103,30,162,31,50,31,55,31,219,31,254,31,119,31,44,31,44,30,107,31,107,30,107,29,117,31,212,31,212,30,221,31,240,31,249,31,229,31,238,31,217,31,48,31,48,30,155,31,245,31,122,31,219,31,25,31,52,31,245,31,82,31,83,31,83,30,83,29,241,31,245,31,79,31,65,31,20,31,54,31,201,31,207,31,26,31,26,30,26,29,32,31,88,31,158,31,13,31,2,31,35,31,174,31,174,30,246,31,246,30,66,31,109,31,109,30,109,29,143,31,147,31,95,31,3,31,183,31,146,31,110,31,137,31,170,31,156,31,212,31,114,31,153,31,187,31,136,31,163,31,152,31,18,31,24,31,63,31,246,31,211,31,45,31,194,31,94,31,221,31,89,31,29,31,45,31,125,31,173,31,173,30,218,31,156,31,55,31,117,31,180,31,63,31,47,31,255,31,255,30,234,31,119,31,251,31,64,31,161,31,241,31,7,31,7,30,41,31,148,31,255,31,161,31,161,30,161,29,70,31,120,31,244,31,244,30,218,31,191,31,246,31,63,31,186,31,186,30,121,31,140,31,140,30,158,31,130,31,109,31,118,31,213,31,129,31,129,30,127,31,45,31,206,31,38,31,212,31,236,31,192,31,192,30,71,31,71,30,52,31,128,31,176,31,224,31,230,31,76,31,242,31,203,31,9,31,242,31,132,31,245,31,222,31,196,31,16,31,40,31,111,31,242,31,164,31,134,31,134,30,48,31,25,31,25,30,184,31,31,31,215,31,199,31,46,31,87,31,7,31,7,30,40,31,187,31,23,31,173,31,13,31,216,31,44,31,161,31,161,31,51,31,15,31,28,31,28,30,204,31,204,30,171,31,171,30,131,31,23,31,237,31,207,31,11,31,197,31,197,30,79,31,22,31,130,31,84,31,195,31,238,31,123,31,56,31,221,31,10,31,127,31,154,31,173,31,236,31,128,31,128,30,182,31,47,31,242,31,242,30,167,31,178,31,41,31,217,31,121,31,68,31,176,31,211,31,25,31,159,31,76,31,76,30,68,31,68,30,178,31,17,31,18,31,71,31,159,31,1,31,1,30,1,29,1,28,184,31,184,30,224,31,186,31,186,30,186,31,186,30,186,29,154,31,229,31,222,31,159,31,223,31,253,31,59,31,32,31,159,31,152,31,77,31,77,30,242,31,242,30,98,31,20,31,59,31,59,30,88,31,50,31,29,31,206,31,112,31,245,31,209,31,48,31,237,31,176,31,155,31,95,31,1,31,159,31,70,31,222,31,147,31,74,31,104,31,169,31,181,31,126,31,144,31,159,31,29,31,41,31,41,30,214,31,116,31,116,30,116,29,160,31,10,31,46,31,13,31,147,31,74,31,241,31,173,31,79,31,147,31,61,31,77,31,77,30,235,31,118,31,36,31,36,30,36,29,36,28,109,31,135,31,135,30,30,31,31,31,117,31,230,31,230,30,172,31,172,30,245,31,42,31,61,31,239,31,239,30,239,29,76,31,28,31,233,31,105,31,117,31,117,30,117,29,184,31,184,30,41,31,177,31,106,31,136,31,127,31,127,30,126,31,103,31,74,31,42,31,201,31,201,30,201,29,178,31,178,30,16,31,16,30,16,29,16,28,66,31,237,31,39,31,21,31,23,31,34,31,34,30,188,31,51,31,51,30,188,31,170,31,168,31,71,31,71,30,107,31,90,31,90,30,30,31,141,31,115,31,29,31,111,31,93,31,201,31,201,30,201,29,25,31,25,30,53,31,175,31,34,31,84,31,223,31,85,31,22,31,22,30,75,31,75,30,91,31,78,31,253,31,71,31,137,31,100,31,251,31,72,31,154,31,230,31,214,31,206,31,206,30,238,31,210,31,210,30,168,31,58,31,162,31,10,31,10,30,111,31,237,31,232,31,156,31,150,31,34,31,61,31,114,31,108,31,108,30,140,31,37,31,78,31,146,31,36,31,148,31,63,31,195,31,23,31,27,31,185,31,185,30,152,31,152,30,143,31,143,30,230,31,26,31,162,31,129,31,231,31,165,31,165,30,165,29,114,31,206,31,167,31,95,31,86,31,86,30,142,31,142,30,142,29,199,31,72,31,246,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
