-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_90 is
end project_tb_90;

architecture project_tb_arch_90 of project_tb_90 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 999;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (182,0,6,0,106,0,224,0,0,0,24,0,46,0,0,0,21,0,0,0,8,0,149,0,104,0,0,0,0,0,0,0,37,0,0,0,0,0,83,0,140,0,199,0,0,0,106,0,60,0,0,0,5,0,178,0,0,0,157,0,68,0,240,0,100,0,134,0,147,0,0,0,0,0,90,0,103,0,250,0,244,0,0,0,0,0,95,0,90,0,39,0,117,0,126,0,169,0,0,0,175,0,1,0,107,0,198,0,47,0,147,0,24,0,141,0,245,0,126,0,198,0,114,0,16,0,54,0,234,0,131,0,48,0,242,0,0,0,175,0,0,0,191,0,129,0,98,0,115,0,137,0,0,0,204,0,147,0,0,0,250,0,0,0,245,0,0,0,32,0,0,0,0,0,0,0,95,0,0,0,112,0,122,0,88,0,109,0,138,0,0,0,222,0,204,0,161,0,0,0,0,0,24,0,120,0,174,0,246,0,0,0,29,0,0,0,44,0,25,0,0,0,184,0,213,0,0,0,165,0,174,0,64,0,0,0,88,0,107,0,229,0,217,0,206,0,240,0,97,0,230,0,240,0,101,0,0,0,92,0,112,0,180,0,207,0,233,0,0,0,0,0,38,0,0,0,52,0,193,0,52,0,170,0,34,0,4,0,215,0,90,0,0,0,66,0,181,0,29,0,81,0,243,0,242,0,0,0,14,0,122,0,118,0,61,0,184,0,0,0,128,0,8,0,86,0,74,0,44,0,0,0,64,0,0,0,0,0,12,0,0,0,108,0,0,0,0,0,184,0,34,0,151,0,113,0,242,0,222,0,202,0,240,0,69,0,0,0,0,0,0,0,197,0,41,0,108,0,148,0,247,0,0,0,0,0,188,0,99,0,0,0,145,0,252,0,206,0,155,0,79,0,152,0,0,0,216,0,0,0,217,0,248,0,40,0,0,0,240,0,57,0,91,0,225,0,77,0,245,0,158,0,94,0,0,0,174,0,39,0,203,0,237,0,78,0,0,0,144,0,168,0,0,0,62,0,151,0,139,0,225,0,68,0,219,0,58,0,118,0,246,0,221,0,5,0,22,0,67,0,192,0,236,0,111,0,0,0,146,0,100,0,212,0,96,0,77,0,62,0,102,0,53,0,45,0,143,0,222,0,237,0,181,0,0,0,22,0,19,0,0,0,76,0,38,0,44,0,0,0,226,0,60,0,92,0,46,0,106,0,51,0,234,0,228,0,153,0,0,0,141,0,212,0,0,0,106,0,124,0,81,0,6,0,0,0,109,0,0,0,42,0,228,0,146,0,0,0,90,0,74,0,161,0,95,0,164,0,0,0,192,0,5,0,25,0,0,0,101,0,179,0,251,0,24,0,154,0,127,0,0,0,197,0,67,0,67,0,136,0,72,0,173,0,0,0,0,0,0,0,47,0,14,0,125,0,216,0,0,0,12,0,0,0,17,0,0,0,211,0,0,0,0,0,115,0,29,0,38,0,0,0,0,0,253,0,166,0,73,0,147,0,171,0,141,0,0,0,0,0,224,0,203,0,0,0,153,0,0,0,212,0,180,0,85,0,239,0,255,0,216,0,25,0,142,0,246,0,0,0,59,0,21,0,60,0,70,0,0,0,4,0,21,0,242,0,195,0,200,0,0,0,37,0,0,0,139,0,55,0,198,0,173,0,0,0,66,0,43,0,41,0,12,0,78,0,191,0,95,0,117,0,0,0,10,0,224,0,251,0,53,0,218,0,0,0,16,0,84,0,72,0,210,0,182,0,248,0,95,0,26,0,0,0,99,0,115,0,247,0,220,0,9,0,9,0,255,0,104,0,0,0,0,0,224,0,244,0,184,0,39,0,43,0,170,0,0,0,0,0,127,0,238,0,0,0,28,0,183,0,179,0,124,0,103,0,160,0,36,0,100,0,72,0,97,0,223,0,52,0,0,0,233,0,190,0,178,0,251,0,134,0,0,0,110,0,7,0,189,0,163,0,130,0,49,0,76,0,232,0,184,0,225,0,154,0,194,0,170,0,0,0,241,0,0,0,237,0,0,0,0,0,53,0,29,0,110,0,248,0,114,0,206,0,29,0,160,0,200,0,61,0,10,0,236,0,199,0,100,0,0,0,52,0,233,0,168,0,0,0,44,0,86,0,48,0,8,0,24,0,253,0,16,0,0,0,0,0,122,0,3,0,184,0,14,0,249,0,114,0,0,0,239,0,239,0,53,0,0,0,77,0,18,0,198,0,36,0,15,0,6,0,82,0,141,0,33,0,10,0,132,0,35,0,11,0,166,0,206,0,117,0,140,0,139,0,165,0,141,0,0,0,0,0,187,0,204,0,179,0,0,0,248,0,0,0,26,0,0,0,0,0,239,0,189,0,57,0,221,0,0,0,139,0,89,0,0,0,52,0,62,0,67,0,189,0,176,0,124,0,82,0,189,0,245,0,19,0,110,0,119,0,169,0,164,0,176,0,0,0,12,0,157,0,210,0,88,0,97,0,0,0,14,0,59,0,204,0,146,0,89,0,0,0,0,0,123,0,205,0,40,0,74,0,39,0,189,0,159,0,162,0,205,0,28,0,0,0,108,0,0,0,250,0,189,0,218,0,0,0,78,0,226,0,210,0,44,0,16,0,39,0,96,0,195,0,145,0,0,0,92,0,12,0,185,0,150,0,0,0,27,0,0,0,46,0,39,0,0,0,88,0,254,0,0,0,0,0,36,0,93,0,170,0,217,0,117,0,191,0,246,0,84,0,0,0,177,0,0,0,0,0,0,0,71,0,63,0,0,0,0,0,195,0,0,0,234,0,90,0,75,0,205,0,30,0,195,0,42,0,232,0,0,0,157,0,0,0,137,0,192,0,206,0,100,0,143,0,107,0,169,0,168,0,224,0,78,0,0,0,1,0,168,0,64,0,175,0,5,0,54,0,177,0,104,0,0,0,16,0,0,0,131,0,240,0,21,0,20,0,23,0,66,0,0,0,163,0,0,0,62,0,90,0,6,0,65,0,60,0,0,0,85,0,94,0,147,0,150,0,0,0,0,0,39,0,0,0,236,0,185,0,58,0,145,0,94,0,32,0,38,0,0,0,0,0,57,0,0,0,84,0,120,0,171,0,124,0,61,0,0,0,218,0,53,0,146,0,100,0,155,0,253,0,234,0,230,0,197,0,7,0,8,0,0,0,0,0,0,0,24,0,247,0,133,0,207,0,213,0,91,0,127,0,0,0,139,0,0,0,249,0,187,0,254,0,0,0,14,0,210,0,0,0,184,0,179,0,42,0,235,0,220,0,205,0,188,0,73,0,146,0,152,0,92,0,2,0,255,0,0,0,90,0,69,0,61,0,159,0,0,0,127,0,0,0,37,0,122,0,99,0,29,0,0,0,213,0,247,0,0,0,96,0,5,0,46,0,0,0,91,0,202,0,55,0,0,0,150,0,219,0,190,0,31,0,89,0,91,0,51,0,232,0,137,0,31,0,102,0,18,0,14,0,213,0,231,0,84,0,232,0,83,0,132,0,110,0,0,0,4,0,86,0,0,0,0,0,45,0,0,0,170,0,103,0,206,0,252,0,199,0,0,0,0,0,0,0,189,0,43,0,240,0,143,0,3,0,20,0,98,0,18,0,0,0,178,0,59,0,62,0,129,0,38,0,0,0,69,0,77,0,205,0,216,0,127,0,89,0,174,0,13,0,61,0,16,0,226,0,236,0,89,0,253,0,0,0,119,0,235,0,104,0,231,0,120,0,85,0,218,0,0,0,188,0,79,0,23,0,104,0,24,0,24,0,132,0,0,0,218,0,236,0,106,0,0,0,169,0,135,0,0,0,175,0,10,0,214,0,194,0,0,0,58,0,226,0,14,0,75,0,141,0,58,0,63,0,0,0,211,0,0,0,0,0,40,0,11,0,0,0,167,0,66,0,0,0,110,0,37,0,137,0,123,0,69,0,0,0,64,0,133,0,204,0,0,0,224,0,71,0,83,0,66,0,174,0,0,0,207,0,73,0,0,0,120,0,82,0,220,0,93,0,131,0,0,0,106,0,24,0,43,0,0,0,15,0,79,0,68,0,108,0,168,0,0,0,128,0,90,0,45,0,88,0,181,0,70,0,109,0,0,0,115,0,88,0,126,0,129,0,84,0,121,0,0,0,84,0,104,0,165,0,0,0,172,0,42,0,214,0,61,0,102,0,35,0,227,0,137,0,71,0,156,0,18,0,29,0,54,0,228,0,0,0,111,0,146,0,0,0,43,0,94,0,0,0,0,0,173,0,57,0,87,0,233,0,0,0,35,0,43,0,203,0,114,0,190,0,245,0,111,0,126,0,177,0,37,0,191,0,75,0,0,0,67,0,139,0,169,0,140,0,0,0,192,0,87,0,22,0,121,0,209,0,160,0,239,0,218,0,0,0,204,0,157,0,74,0,202,0,4,0,3,0,0,0,90,0,249,0,0,0,109,0,54,0,247,0,254,0,172,0,219,0,237,0);
signal scenario_full  : scenario_type := (182,31,6,31,106,31,224,31,224,30,24,31,46,31,46,30,21,31,21,30,8,31,149,31,104,31,104,30,104,29,104,28,37,31,37,30,37,29,83,31,140,31,199,31,199,30,106,31,60,31,60,30,5,31,178,31,178,30,157,31,68,31,240,31,100,31,134,31,147,31,147,30,147,29,90,31,103,31,250,31,244,31,244,30,244,29,95,31,90,31,39,31,117,31,126,31,169,31,169,30,175,31,1,31,107,31,198,31,47,31,147,31,24,31,141,31,245,31,126,31,198,31,114,31,16,31,54,31,234,31,131,31,48,31,242,31,242,30,175,31,175,30,191,31,129,31,98,31,115,31,137,31,137,30,204,31,147,31,147,30,250,31,250,30,245,31,245,30,32,31,32,30,32,29,32,28,95,31,95,30,112,31,122,31,88,31,109,31,138,31,138,30,222,31,204,31,161,31,161,30,161,29,24,31,120,31,174,31,246,31,246,30,29,31,29,30,44,31,25,31,25,30,184,31,213,31,213,30,165,31,174,31,64,31,64,30,88,31,107,31,229,31,217,31,206,31,240,31,97,31,230,31,240,31,101,31,101,30,92,31,112,31,180,31,207,31,233,31,233,30,233,29,38,31,38,30,52,31,193,31,52,31,170,31,34,31,4,31,215,31,90,31,90,30,66,31,181,31,29,31,81,31,243,31,242,31,242,30,14,31,122,31,118,31,61,31,184,31,184,30,128,31,8,31,86,31,74,31,44,31,44,30,64,31,64,30,64,29,12,31,12,30,108,31,108,30,108,29,184,31,34,31,151,31,113,31,242,31,222,31,202,31,240,31,69,31,69,30,69,29,69,28,197,31,41,31,108,31,148,31,247,31,247,30,247,29,188,31,99,31,99,30,145,31,252,31,206,31,155,31,79,31,152,31,152,30,216,31,216,30,217,31,248,31,40,31,40,30,240,31,57,31,91,31,225,31,77,31,245,31,158,31,94,31,94,30,174,31,39,31,203,31,237,31,78,31,78,30,144,31,168,31,168,30,62,31,151,31,139,31,225,31,68,31,219,31,58,31,118,31,246,31,221,31,5,31,22,31,67,31,192,31,236,31,111,31,111,30,146,31,100,31,212,31,96,31,77,31,62,31,102,31,53,31,45,31,143,31,222,31,237,31,181,31,181,30,22,31,19,31,19,30,76,31,38,31,44,31,44,30,226,31,60,31,92,31,46,31,106,31,51,31,234,31,228,31,153,31,153,30,141,31,212,31,212,30,106,31,124,31,81,31,6,31,6,30,109,31,109,30,42,31,228,31,146,31,146,30,90,31,74,31,161,31,95,31,164,31,164,30,192,31,5,31,25,31,25,30,101,31,179,31,251,31,24,31,154,31,127,31,127,30,197,31,67,31,67,31,136,31,72,31,173,31,173,30,173,29,173,28,47,31,14,31,125,31,216,31,216,30,12,31,12,30,17,31,17,30,211,31,211,30,211,29,115,31,29,31,38,31,38,30,38,29,253,31,166,31,73,31,147,31,171,31,141,31,141,30,141,29,224,31,203,31,203,30,153,31,153,30,212,31,180,31,85,31,239,31,255,31,216,31,25,31,142,31,246,31,246,30,59,31,21,31,60,31,70,31,70,30,4,31,21,31,242,31,195,31,200,31,200,30,37,31,37,30,139,31,55,31,198,31,173,31,173,30,66,31,43,31,41,31,12,31,78,31,191,31,95,31,117,31,117,30,10,31,224,31,251,31,53,31,218,31,218,30,16,31,84,31,72,31,210,31,182,31,248,31,95,31,26,31,26,30,99,31,115,31,247,31,220,31,9,31,9,31,255,31,104,31,104,30,104,29,224,31,244,31,184,31,39,31,43,31,170,31,170,30,170,29,127,31,238,31,238,30,28,31,183,31,179,31,124,31,103,31,160,31,36,31,100,31,72,31,97,31,223,31,52,31,52,30,233,31,190,31,178,31,251,31,134,31,134,30,110,31,7,31,189,31,163,31,130,31,49,31,76,31,232,31,184,31,225,31,154,31,194,31,170,31,170,30,241,31,241,30,237,31,237,30,237,29,53,31,29,31,110,31,248,31,114,31,206,31,29,31,160,31,200,31,61,31,10,31,236,31,199,31,100,31,100,30,52,31,233,31,168,31,168,30,44,31,86,31,48,31,8,31,24,31,253,31,16,31,16,30,16,29,122,31,3,31,184,31,14,31,249,31,114,31,114,30,239,31,239,31,53,31,53,30,77,31,18,31,198,31,36,31,15,31,6,31,82,31,141,31,33,31,10,31,132,31,35,31,11,31,166,31,206,31,117,31,140,31,139,31,165,31,141,31,141,30,141,29,187,31,204,31,179,31,179,30,248,31,248,30,26,31,26,30,26,29,239,31,189,31,57,31,221,31,221,30,139,31,89,31,89,30,52,31,62,31,67,31,189,31,176,31,124,31,82,31,189,31,245,31,19,31,110,31,119,31,169,31,164,31,176,31,176,30,12,31,157,31,210,31,88,31,97,31,97,30,14,31,59,31,204,31,146,31,89,31,89,30,89,29,123,31,205,31,40,31,74,31,39,31,189,31,159,31,162,31,205,31,28,31,28,30,108,31,108,30,250,31,189,31,218,31,218,30,78,31,226,31,210,31,44,31,16,31,39,31,96,31,195,31,145,31,145,30,92,31,12,31,185,31,150,31,150,30,27,31,27,30,46,31,39,31,39,30,88,31,254,31,254,30,254,29,36,31,93,31,170,31,217,31,117,31,191,31,246,31,84,31,84,30,177,31,177,30,177,29,177,28,71,31,63,31,63,30,63,29,195,31,195,30,234,31,90,31,75,31,205,31,30,31,195,31,42,31,232,31,232,30,157,31,157,30,137,31,192,31,206,31,100,31,143,31,107,31,169,31,168,31,224,31,78,31,78,30,1,31,168,31,64,31,175,31,5,31,54,31,177,31,104,31,104,30,16,31,16,30,131,31,240,31,21,31,20,31,23,31,66,31,66,30,163,31,163,30,62,31,90,31,6,31,65,31,60,31,60,30,85,31,94,31,147,31,150,31,150,30,150,29,39,31,39,30,236,31,185,31,58,31,145,31,94,31,32,31,38,31,38,30,38,29,57,31,57,30,84,31,120,31,171,31,124,31,61,31,61,30,218,31,53,31,146,31,100,31,155,31,253,31,234,31,230,31,197,31,7,31,8,31,8,30,8,29,8,28,24,31,247,31,133,31,207,31,213,31,91,31,127,31,127,30,139,31,139,30,249,31,187,31,254,31,254,30,14,31,210,31,210,30,184,31,179,31,42,31,235,31,220,31,205,31,188,31,73,31,146,31,152,31,92,31,2,31,255,31,255,30,90,31,69,31,61,31,159,31,159,30,127,31,127,30,37,31,122,31,99,31,29,31,29,30,213,31,247,31,247,30,96,31,5,31,46,31,46,30,91,31,202,31,55,31,55,30,150,31,219,31,190,31,31,31,89,31,91,31,51,31,232,31,137,31,31,31,102,31,18,31,14,31,213,31,231,31,84,31,232,31,83,31,132,31,110,31,110,30,4,31,86,31,86,30,86,29,45,31,45,30,170,31,103,31,206,31,252,31,199,31,199,30,199,29,199,28,189,31,43,31,240,31,143,31,3,31,20,31,98,31,18,31,18,30,178,31,59,31,62,31,129,31,38,31,38,30,69,31,77,31,205,31,216,31,127,31,89,31,174,31,13,31,61,31,16,31,226,31,236,31,89,31,253,31,253,30,119,31,235,31,104,31,231,31,120,31,85,31,218,31,218,30,188,31,79,31,23,31,104,31,24,31,24,31,132,31,132,30,218,31,236,31,106,31,106,30,169,31,135,31,135,30,175,31,10,31,214,31,194,31,194,30,58,31,226,31,14,31,75,31,141,31,58,31,63,31,63,30,211,31,211,30,211,29,40,31,11,31,11,30,167,31,66,31,66,30,110,31,37,31,137,31,123,31,69,31,69,30,64,31,133,31,204,31,204,30,224,31,71,31,83,31,66,31,174,31,174,30,207,31,73,31,73,30,120,31,82,31,220,31,93,31,131,31,131,30,106,31,24,31,43,31,43,30,15,31,79,31,68,31,108,31,168,31,168,30,128,31,90,31,45,31,88,31,181,31,70,31,109,31,109,30,115,31,88,31,126,31,129,31,84,31,121,31,121,30,84,31,104,31,165,31,165,30,172,31,42,31,214,31,61,31,102,31,35,31,227,31,137,31,71,31,156,31,18,31,29,31,54,31,228,31,228,30,111,31,146,31,146,30,43,31,94,31,94,30,94,29,173,31,57,31,87,31,233,31,233,30,35,31,43,31,203,31,114,31,190,31,245,31,111,31,126,31,177,31,37,31,191,31,75,31,75,30,67,31,139,31,169,31,140,31,140,30,192,31,87,31,22,31,121,31,209,31,160,31,239,31,218,31,218,30,204,31,157,31,74,31,202,31,4,31,3,31,3,30,90,31,249,31,249,30,109,31,54,31,247,31,254,31,172,31,219,31,237,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
