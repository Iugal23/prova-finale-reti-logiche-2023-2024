-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 891;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,2,0,0,0,119,0,83,0,0,0,188,0,96,0,0,0,140,0,226,0,54,0,0,0,184,0,0,0,110,0,38,0,31,0,255,0,0,0,163,0,0,0,0,0,133,0,198,0,102,0,0,0,0,0,83,0,0,0,142,0,0,0,0,0,137,0,105,0,77,0,221,0,18,0,182,0,0,0,62,0,2,0,0,0,219,0,255,0,44,0,0,0,245,0,73,0,175,0,151,0,2,0,0,0,0,0,6,0,57,0,67,0,214,0,0,0,20,0,216,0,187,0,212,0,91,0,204,0,126,0,177,0,0,0,159,0,93,0,0,0,194,0,185,0,0,0,143,0,68,0,0,0,226,0,72,0,11,0,0,0,77,0,74,0,229,0,132,0,161,0,136,0,0,0,37,0,80,0,0,0,42,0,248,0,22,0,0,0,206,0,240,0,175,0,106,0,140,0,0,0,93,0,55,0,16,0,54,0,23,0,213,0,46,0,193,0,182,0,7,0,46,0,72,0,83,0,179,0,254,0,230,0,31,0,166,0,0,0,70,0,0,0,80,0,203,0,111,0,110,0,206,0,124,0,86,0,0,0,187,0,238,0,108,0,0,0,49,0,25,0,0,0,97,0,25,0,148,0,121,0,0,0,64,0,0,0,168,0,83,0,0,0,164,0,73,0,127,0,0,0,0,0,166,0,0,0,205,0,0,0,38,0,0,0,143,0,157,0,105,0,0,0,141,0,0,0,192,0,5,0,77,0,17,0,0,0,165,0,182,0,0,0,0,0,9,0,118,0,143,0,0,0,0,0,233,0,154,0,222,0,194,0,22,0,185,0,0,0,86,0,3,0,14,0,179,0,117,0,37,0,0,0,0,0,0,0,79,0,160,0,0,0,253,0,26,0,106,0,132,0,81,0,78,0,0,0,167,0,255,0,65,0,240,0,23,0,57,0,0,0,92,0,214,0,143,0,0,0,68,0,3,0,166,0,140,0,148,0,94,0,226,0,57,0,143,0,70,0,0,0,122,0,149,0,182,0,196,0,96,0,161,0,0,0,213,0,236,0,250,0,63,0,185,0,198,0,0,0,102,0,114,0,96,0,114,0,65,0,184,0,95,0,0,0,70,0,24,0,22,0,50,0,113,0,0,0,37,0,171,0,191,0,161,0,3,0,199,0,248,0,186,0,0,0,146,0,234,0,38,0,118,0,135,0,233,0,226,0,244,0,180,0,190,0,132,0,88,0,140,0,40,0,154,0,0,0,222,0,20,0,118,0,0,0,150,0,0,0,200,0,150,0,130,0,88,0,199,0,226,0,9,0,237,0,184,0,142,0,0,0,96,0,171,0,229,0,217,0,0,0,154,0,69,0,180,0,79,0,222,0,0,0,75,0,90,0,13,0,10,0,0,0,190,0,0,0,218,0,206,0,204,0,221,0,237,0,0,0,32,0,103,0,0,0,85,0,197,0,170,0,75,0,124,0,97,0,167,0,202,0,167,0,103,0,172,0,205,0,72,0,148,0,229,0,96,0,202,0,240,0,91,0,141,0,77,0,87,0,252,0,172,0,80,0,0,0,179,0,169,0,73,0,139,0,0,0,39,0,99,0,11,0,216,0,139,0,129,0,162,0,9,0,60,0,42,0,227,0,0,0,97,0,133,0,111,0,0,0,174,0,115,0,0,0,15,0,204,0,227,0,66,0,0,0,164,0,112,0,53,0,147,0,122,0,17,0,51,0,0,0,186,0,55,0,107,0,3,0,26,0,62,0,0,0,0,0,237,0,114,0,137,0,251,0,165,0,176,0,237,0,47,0,118,0,0,0,69,0,222,0,235,0,13,0,142,0,55,0,124,0,150,0,49,0,58,0,177,0,190,0,55,0,0,0,35,0,47,0,0,0,194,0,84,0,216,0,233,0,49,0,219,0,55,0,0,0,31,0,191,0,107,0,176,0,0,0,66,0,205,0,0,0,247,0,119,0,101,0,185,0,97,0,0,0,101,0,12,0,49,0,180,0,150,0,45,0,246,0,13,0,215,0,124,0,199,0,0,0,66,0,104,0,171,0,0,0,0,0,193,0,0,0,163,0,44,0,119,0,224,0,239,0,238,0,114,0,130,0,0,0,0,0,0,0,0,0,125,0,134,0,85,0,70,0,29,0,174,0,31,0,6,0,164,0,201,0,87,0,0,0,0,0,214,0,211,0,175,0,46,0,0,0,32,0,235,0,80,0,0,0,217,0,0,0,0,0,153,0,58,0,18,0,114,0,225,0,140,0,31,0,143,0,102,0,58,0,186,0,201,0,132,0,234,0,44,0,0,0,97,0,0,0,234,0,0,0,229,0,0,0,32,0,184,0,59,0,48,0,145,0,26,0,0,0,244,0,148,0,141,0,0,0,70,0,243,0,5,0,183,0,0,0,249,0,95,0,231,0,230,0,46,0,63,0,104,0,203,0,80,0,0,0,0,0,0,0,114,0,171,0,48,0,15,0,55,0,12,0,35,0,5,0,55,0,211,0,231,0,183,0,0,0,105,0,85,0,231,0,190,0,65,0,175,0,125,0,150,0,90,0,0,0,33,0,0,0,0,0,216,0,122,0,196,0,54,0,0,0,232,0,242,0,72,0,151,0,36,0,44,0,0,0,49,0,201,0,67,0,219,0,234,0,0,0,110,0,147,0,0,0,213,0,245,0,22,0,69,0,5,0,44,0,80,0,47,0,0,0,213,0,194,0,0,0,176,0,0,0,0,0,67,0,172,0,89,0,113,0,0,0,0,0,209,0,29,0,40,0,28,0,15,0,74,0,148,0,10,0,0,0,129,0,125,0,0,0,196,0,210,0,208,0,0,0,36,0,201,0,179,0,196,0,0,0,55,0,99,0,144,0,97,0,40,0,48,0,126,0,112,0,41,0,132,0,121,0,217,0,48,0,94,0,0,0,111,0,0,0,29,0,181,0,0,0,188,0,0,0,208,0,194,0,178,0,80,0,29,0,0,0,188,0,153,0,255,0,96,0,167,0,0,0,219,0,70,0,220,0,148,0,0,0,87,0,121,0,0,0,59,0,0,0,74,0,0,0,0,0,6,0,0,0,240,0,53,0,0,0,197,0,172,0,16,0,99,0,104,0,45,0,8,0,212,0,27,0,232,0,126,0,15,0,16,0,81,0,0,0,0,0,73,0,0,0,241,0,46,0,0,0,147,0,15,0,0,0,154,0,213,0,0,0,0,0,138,0,76,0,12,0,1,0,45,0,48,0,141,0,182,0,0,0,46,0,0,0,0,0,152,0,237,0,0,0,0,0,27,0,139,0,245,0,48,0,254,0,199,0,0,0,0,0,143,0,86,0,192,0,102,0,84,0,81,0,159,0,31,0,110,0,25,0,169,0,0,0,49,0,240,0,211,0,56,0,237,0,121,0,35,0,192,0,165,0,40,0,50,0,208,0,250,0,104,0,171,0,69,0,0,0,211,0,13,0,206,0,157,0,250,0,14,0,159,0,0,0,176,0,0,0,0,0,91,0,209,0,164,0,0,0,72,0,195,0,145,0,0,0,147,0,158,0,181,0,210,0,78,0,78,0,208,0,68,0,0,0,196,0,161,0,19,0,209,0,5,0,224,0,172,0,224,0,45,0,185,0,0,0,30,0,224,0,0,0,217,0,175,0,23,0,0,0,0,0,0,0,115,0,5,0,41,0,200,0,211,0,206,0,204,0,33,0,0,0,26,0,55,0,225,0,19,0,185,0,132,0,0,0,74,0,44,0,236,0,57,0,84,0,0,0,0,0,163,0,68,0,66,0,0,0,230,0,235,0,23,0,95,0,0,0,223,0,17,0,40,0,101,0,238,0,255,0,210,0,136,0,194,0,209,0,23,0,118,0,0,0,108,0,0,0,191,0,167,0,248,0,17,0,37,0,182,0,165,0,136,0,233,0,220,0,0,0,232,0,161,0,0,0,120,0,35,0,7,0,49,0,71,0,141,0,235,0,200,0,191,0,183,0,203,0);
signal scenario_full  : scenario_type := (0,0,2,31,2,30,119,31,83,31,83,30,188,31,96,31,96,30,140,31,226,31,54,31,54,30,184,31,184,30,110,31,38,31,31,31,255,31,255,30,163,31,163,30,163,29,133,31,198,31,102,31,102,30,102,29,83,31,83,30,142,31,142,30,142,29,137,31,105,31,77,31,221,31,18,31,182,31,182,30,62,31,2,31,2,30,219,31,255,31,44,31,44,30,245,31,73,31,175,31,151,31,2,31,2,30,2,29,6,31,57,31,67,31,214,31,214,30,20,31,216,31,187,31,212,31,91,31,204,31,126,31,177,31,177,30,159,31,93,31,93,30,194,31,185,31,185,30,143,31,68,31,68,30,226,31,72,31,11,31,11,30,77,31,74,31,229,31,132,31,161,31,136,31,136,30,37,31,80,31,80,30,42,31,248,31,22,31,22,30,206,31,240,31,175,31,106,31,140,31,140,30,93,31,55,31,16,31,54,31,23,31,213,31,46,31,193,31,182,31,7,31,46,31,72,31,83,31,179,31,254,31,230,31,31,31,166,31,166,30,70,31,70,30,80,31,203,31,111,31,110,31,206,31,124,31,86,31,86,30,187,31,238,31,108,31,108,30,49,31,25,31,25,30,97,31,25,31,148,31,121,31,121,30,64,31,64,30,168,31,83,31,83,30,164,31,73,31,127,31,127,30,127,29,166,31,166,30,205,31,205,30,38,31,38,30,143,31,157,31,105,31,105,30,141,31,141,30,192,31,5,31,77,31,17,31,17,30,165,31,182,31,182,30,182,29,9,31,118,31,143,31,143,30,143,29,233,31,154,31,222,31,194,31,22,31,185,31,185,30,86,31,3,31,14,31,179,31,117,31,37,31,37,30,37,29,37,28,79,31,160,31,160,30,253,31,26,31,106,31,132,31,81,31,78,31,78,30,167,31,255,31,65,31,240,31,23,31,57,31,57,30,92,31,214,31,143,31,143,30,68,31,3,31,166,31,140,31,148,31,94,31,226,31,57,31,143,31,70,31,70,30,122,31,149,31,182,31,196,31,96,31,161,31,161,30,213,31,236,31,250,31,63,31,185,31,198,31,198,30,102,31,114,31,96,31,114,31,65,31,184,31,95,31,95,30,70,31,24,31,22,31,50,31,113,31,113,30,37,31,171,31,191,31,161,31,3,31,199,31,248,31,186,31,186,30,146,31,234,31,38,31,118,31,135,31,233,31,226,31,244,31,180,31,190,31,132,31,88,31,140,31,40,31,154,31,154,30,222,31,20,31,118,31,118,30,150,31,150,30,200,31,150,31,130,31,88,31,199,31,226,31,9,31,237,31,184,31,142,31,142,30,96,31,171,31,229,31,217,31,217,30,154,31,69,31,180,31,79,31,222,31,222,30,75,31,90,31,13,31,10,31,10,30,190,31,190,30,218,31,206,31,204,31,221,31,237,31,237,30,32,31,103,31,103,30,85,31,197,31,170,31,75,31,124,31,97,31,167,31,202,31,167,31,103,31,172,31,205,31,72,31,148,31,229,31,96,31,202,31,240,31,91,31,141,31,77,31,87,31,252,31,172,31,80,31,80,30,179,31,169,31,73,31,139,31,139,30,39,31,99,31,11,31,216,31,139,31,129,31,162,31,9,31,60,31,42,31,227,31,227,30,97,31,133,31,111,31,111,30,174,31,115,31,115,30,15,31,204,31,227,31,66,31,66,30,164,31,112,31,53,31,147,31,122,31,17,31,51,31,51,30,186,31,55,31,107,31,3,31,26,31,62,31,62,30,62,29,237,31,114,31,137,31,251,31,165,31,176,31,237,31,47,31,118,31,118,30,69,31,222,31,235,31,13,31,142,31,55,31,124,31,150,31,49,31,58,31,177,31,190,31,55,31,55,30,35,31,47,31,47,30,194,31,84,31,216,31,233,31,49,31,219,31,55,31,55,30,31,31,191,31,107,31,176,31,176,30,66,31,205,31,205,30,247,31,119,31,101,31,185,31,97,31,97,30,101,31,12,31,49,31,180,31,150,31,45,31,246,31,13,31,215,31,124,31,199,31,199,30,66,31,104,31,171,31,171,30,171,29,193,31,193,30,163,31,44,31,119,31,224,31,239,31,238,31,114,31,130,31,130,30,130,29,130,28,130,27,125,31,134,31,85,31,70,31,29,31,174,31,31,31,6,31,164,31,201,31,87,31,87,30,87,29,214,31,211,31,175,31,46,31,46,30,32,31,235,31,80,31,80,30,217,31,217,30,217,29,153,31,58,31,18,31,114,31,225,31,140,31,31,31,143,31,102,31,58,31,186,31,201,31,132,31,234,31,44,31,44,30,97,31,97,30,234,31,234,30,229,31,229,30,32,31,184,31,59,31,48,31,145,31,26,31,26,30,244,31,148,31,141,31,141,30,70,31,243,31,5,31,183,31,183,30,249,31,95,31,231,31,230,31,46,31,63,31,104,31,203,31,80,31,80,30,80,29,80,28,114,31,171,31,48,31,15,31,55,31,12,31,35,31,5,31,55,31,211,31,231,31,183,31,183,30,105,31,85,31,231,31,190,31,65,31,175,31,125,31,150,31,90,31,90,30,33,31,33,30,33,29,216,31,122,31,196,31,54,31,54,30,232,31,242,31,72,31,151,31,36,31,44,31,44,30,49,31,201,31,67,31,219,31,234,31,234,30,110,31,147,31,147,30,213,31,245,31,22,31,69,31,5,31,44,31,80,31,47,31,47,30,213,31,194,31,194,30,176,31,176,30,176,29,67,31,172,31,89,31,113,31,113,30,113,29,209,31,29,31,40,31,28,31,15,31,74,31,148,31,10,31,10,30,129,31,125,31,125,30,196,31,210,31,208,31,208,30,36,31,201,31,179,31,196,31,196,30,55,31,99,31,144,31,97,31,40,31,48,31,126,31,112,31,41,31,132,31,121,31,217,31,48,31,94,31,94,30,111,31,111,30,29,31,181,31,181,30,188,31,188,30,208,31,194,31,178,31,80,31,29,31,29,30,188,31,153,31,255,31,96,31,167,31,167,30,219,31,70,31,220,31,148,31,148,30,87,31,121,31,121,30,59,31,59,30,74,31,74,30,74,29,6,31,6,30,240,31,53,31,53,30,197,31,172,31,16,31,99,31,104,31,45,31,8,31,212,31,27,31,232,31,126,31,15,31,16,31,81,31,81,30,81,29,73,31,73,30,241,31,46,31,46,30,147,31,15,31,15,30,154,31,213,31,213,30,213,29,138,31,76,31,12,31,1,31,45,31,48,31,141,31,182,31,182,30,46,31,46,30,46,29,152,31,237,31,237,30,237,29,27,31,139,31,245,31,48,31,254,31,199,31,199,30,199,29,143,31,86,31,192,31,102,31,84,31,81,31,159,31,31,31,110,31,25,31,169,31,169,30,49,31,240,31,211,31,56,31,237,31,121,31,35,31,192,31,165,31,40,31,50,31,208,31,250,31,104,31,171,31,69,31,69,30,211,31,13,31,206,31,157,31,250,31,14,31,159,31,159,30,176,31,176,30,176,29,91,31,209,31,164,31,164,30,72,31,195,31,145,31,145,30,147,31,158,31,181,31,210,31,78,31,78,31,208,31,68,31,68,30,196,31,161,31,19,31,209,31,5,31,224,31,172,31,224,31,45,31,185,31,185,30,30,31,224,31,224,30,217,31,175,31,23,31,23,30,23,29,23,28,115,31,5,31,41,31,200,31,211,31,206,31,204,31,33,31,33,30,26,31,55,31,225,31,19,31,185,31,132,31,132,30,74,31,44,31,236,31,57,31,84,31,84,30,84,29,163,31,68,31,66,31,66,30,230,31,235,31,23,31,95,31,95,30,223,31,17,31,40,31,101,31,238,31,255,31,210,31,136,31,194,31,209,31,23,31,118,31,118,30,108,31,108,30,191,31,167,31,248,31,17,31,37,31,182,31,165,31,136,31,233,31,220,31,220,30,232,31,161,31,161,30,120,31,35,31,7,31,49,31,71,31,141,31,235,31,200,31,191,31,183,31,203,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
