-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_606 is
end project_tb_606;

architecture project_tb_arch_606 of project_tb_606 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 867;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,59,0,101,0,209,0,1,0,0,0,22,0,22,0,205,0,0,0,60,0,122,0,211,0,198,0,112,0,118,0,109,0,0,0,0,0,251,0,182,0,144,0,119,0,75,0,72,0,23,0,75,0,74,0,203,0,0,0,213,0,235,0,65,0,65,0,0,0,195,0,17,0,205,0,45,0,98,0,146,0,158,0,133,0,0,0,175,0,135,0,241,0,73,0,139,0,0,0,183,0,37,0,76,0,61,0,0,0,249,0,86,0,0,0,233,0,0,0,17,0,127,0,45,0,0,0,62,0,74,0,238,0,0,0,89,0,18,0,0,0,183,0,236,0,143,0,43,0,190,0,125,0,43,0,187,0,23,0,240,0,43,0,206,0,213,0,0,0,47,0,182,0,0,0,216,0,126,0,0,0,5,0,101,0,75,0,151,0,47,0,135,0,96,0,94,0,0,0,172,0,33,0,139,0,96,0,211,0,120,0,177,0,225,0,115,0,0,0,0,0,9,0,203,0,144,0,0,0,0,0,44,0,58,0,0,0,0,0,103,0,102,0,27,0,251,0,134,0,156,0,198,0,81,0,0,0,250,0,47,0,178,0,0,0,201,0,221,0,22,0,19,0,247,0,186,0,219,0,211,0,14,0,210,0,121,0,29,0,0,0,200,0,66,0,58,0,123,0,254,0,85,0,5,0,235,0,25,0,238,0,0,0,96,0,194,0,0,0,246,0,158,0,26,0,158,0,13,0,138,0,169,0,97,0,40,0,108,0,87,0,71,0,0,0,0,0,170,0,226,0,226,0,158,0,0,0,185,0,66,0,153,0,127,0,105,0,80,0,0,0,0,0,49,0,141,0,37,0,54,0,87,0,176,0,58,0,149,0,27,0,97,0,48,0,191,0,210,0,141,0,137,0,93,0,14,0,0,0,227,0,101,0,166,0,49,0,86,0,65,0,0,0,140,0,134,0,202,0,204,0,141,0,251,0,214,0,33,0,175,0,176,0,20,0,95,0,0,0,100,0,186,0,0,0,173,0,175,0,28,0,91,0,17,0,84,0,141,0,54,0,104,0,105,0,60,0,158,0,234,0,42,0,108,0,209,0,148,0,190,0,0,0,0,0,124,0,234,0,221,0,138,0,131,0,222,0,0,0,0,0,48,0,77,0,207,0,0,0,217,0,205,0,146,0,118,0,171,0,0,0,84,0,0,0,0,0,187,0,188,0,84,0,249,0,0,0,97,0,251,0,164,0,96,0,188,0,148,0,67,0,145,0,13,0,133,0,149,0,53,0,0,0,37,0,216,0,70,0,36,0,212,0,192,0,170,0,115,0,31,0,2,0,21,0,0,0,74,0,98,0,92,0,92,0,212,0,0,0,5,0,140,0,221,0,182,0,166,0,117,0,131,0,32,0,108,0,75,0,0,0,60,0,219,0,0,0,0,0,71,0,252,0,28,0,13,0,128,0,249,0,255,0,164,0,111,0,82,0,248,0,26,0,0,0,53,0,134,0,232,0,187,0,101,0,0,0,20,0,54,0,36,0,158,0,204,0,83,0,130,0,0,0,138,0,240,0,242,0,104,0,139,0,137,0,218,0,60,0,0,0,172,0,0,0,0,0,148,0,0,0,0,0,158,0,80,0,0,0,180,0,0,0,99,0,206,0,0,0,37,0,0,0,0,0,20,0,166,0,115,0,211,0,142,0,232,0,152,0,132,0,194,0,223,0,0,0,143,0,0,0,80,0,125,0,58,0,0,0,72,0,159,0,0,0,239,0,172,0,229,0,48,0,0,0,111,0,164,0,0,0,39,0,155,0,210,0,92,0,65,0,200,0,64,0,205,0,77,0,0,0,99,0,0,0,81,0,94,0,176,0,0,0,0,0,0,0,244,0,0,0,0,0,0,0,219,0,181,0,9,0,88,0,0,0,87,0,55,0,105,0,0,0,94,0,197,0,255,0,23,0,0,0,144,0,0,0,123,0,6,0,16,0,192,0,94,0,248,0,230,0,208,0,0,0,79,0,196,0,69,0,100,0,195,0,0,0,167,0,236,0,0,0,0,0,112,0,104,0,183,0,148,0,67,0,31,0,178,0,170,0,2,0,183,0,74,0,101,0,0,0,0,0,138,0,180,0,203,0,168,0,102,0,169,0,95,0,0,0,189,0,132,0,0,0,0,0,65,0,134,0,170,0,31,0,0,0,0,0,0,0,75,0,47,0,75,0,83,0,99,0,51,0,242,0,74,0,135,0,79,0,223,0,138,0,0,0,218,0,236,0,217,0,200,0,101,0,224,0,65,0,80,0,6,0,145,0,212,0,53,0,0,0,222,0,231,0,85,0,217,0,33,0,0,0,24,0,141,0,127,0,221,0,190,0,64,0,93,0,233,0,0,0,213,0,109,0,19,0,0,0,0,0,62,0,114,0,73,0,218,0,202,0,0,0,66,0,31,0,0,0,0,0,89,0,59,0,137,0,218,0,27,0,123,0,218,0,154,0,192,0,236,0,169,0,129,0,2,0,106,0,251,0,185,0,0,0,92,0,200,0,157,0,12,0,192,0,195,0,0,0,21,0,97,0,80,0,0,0,60,0,8,0,127,0,250,0,211,0,148,0,77,0,244,0,0,0,206,0,0,0,232,0,224,0,113,0,23,0,166,0,53,0,72,0,206,0,36,0,0,0,0,0,224,0,0,0,0,0,159,0,116,0,0,0,106,0,152,0,210,0,181,0,150,0,185,0,57,0,8,0,0,0,0,0,0,0,232,0,7,0,32,0,253,0,185,0,96,0,61,0,202,0,113,0,218,0,148,0,86,0,0,0,0,0,230,0,42,0,201,0,86,0,45,0,0,0,88,0,85,0,0,0,109,0,155,0,206,0,126,0,0,0,80,0,125,0,160,0,0,0,175,0,112,0,108,0,14,0,1,0,43,0,58,0,93,0,240,0,61,0,221,0,108,0,0,0,90,0,205,0,0,0,178,0,0,0,251,0,2,0,219,0,197,0,0,0,176,0,248,0,90,0,205,0,0,0,0,0,67,0,164,0,0,0,63,0,85,0,195,0,7,0,117,0,0,0,195,0,159,0,102,0,88,0,26,0,2,0,0,0,111,0,171,0,117,0,0,0,114,0,0,0,240,0,132,0,202,0,126,0,110,0,0,0,197,0,206,0,0,0,214,0,85,0,42,0,194,0,242,0,152,0,118,0,243,0,173,0,224,0,160,0,79,0,56,0,139,0,21,0,245,0,72,0,0,0,190,0,159,0,53,0,78,0,0,0,11,0,204,0,139,0,0,0,205,0,0,0,86,0,191,0,81,0,0,0,224,0,26,0,94,0,0,0,27,0,209,0,71,0,100,0,38,0,207,0,177,0,85,0,177,0,158,0,74,0,0,0,93,0,123,0,161,0,20,0,118,0,240,0,214,0,66,0,188,0,45,0,0,0,114,0,229,0,225,0,197,0,151,0,82,0,195,0,71,0,182,0,0,0,0,0,61,0,148,0,67,0,0,0,32,0,230,0,0,0,249,0,201,0,0,0,82,0,0,0,40,0,77,0,0,0,0,0,91,0,180,0,125,0,254,0,166,0,148,0,202,0,237,0,61,0,230,0,186,0,0,0,46,0,229,0,173,0,0,0,173,0,197,0,238,0,45,0,245,0,83,0,99,0,88,0,34,0,74,0,0,0,195,0,0,0,225,0,101,0,0,0,140,0,119,0,206,0,177,0,0,0,88,0,48,0,247,0,98,0,200,0,0,0,0,0,0,0,158,0,140,0,150,0,24,0,6,0,244,0,122,0,0,0,0,0,204,0,0,0,25,0,0,0,158,0,225,0,66,0,139,0,0,0,0,0,74,0,66,0,182,0,30,0,62,0,75,0,225,0,0,0,0,0,0,0);
signal scenario_full  : scenario_type := (0,0,59,31,101,31,209,31,1,31,1,30,22,31,22,31,205,31,205,30,60,31,122,31,211,31,198,31,112,31,118,31,109,31,109,30,109,29,251,31,182,31,144,31,119,31,75,31,72,31,23,31,75,31,74,31,203,31,203,30,213,31,235,31,65,31,65,31,65,30,195,31,17,31,205,31,45,31,98,31,146,31,158,31,133,31,133,30,175,31,135,31,241,31,73,31,139,31,139,30,183,31,37,31,76,31,61,31,61,30,249,31,86,31,86,30,233,31,233,30,17,31,127,31,45,31,45,30,62,31,74,31,238,31,238,30,89,31,18,31,18,30,183,31,236,31,143,31,43,31,190,31,125,31,43,31,187,31,23,31,240,31,43,31,206,31,213,31,213,30,47,31,182,31,182,30,216,31,126,31,126,30,5,31,101,31,75,31,151,31,47,31,135,31,96,31,94,31,94,30,172,31,33,31,139,31,96,31,211,31,120,31,177,31,225,31,115,31,115,30,115,29,9,31,203,31,144,31,144,30,144,29,44,31,58,31,58,30,58,29,103,31,102,31,27,31,251,31,134,31,156,31,198,31,81,31,81,30,250,31,47,31,178,31,178,30,201,31,221,31,22,31,19,31,247,31,186,31,219,31,211,31,14,31,210,31,121,31,29,31,29,30,200,31,66,31,58,31,123,31,254,31,85,31,5,31,235,31,25,31,238,31,238,30,96,31,194,31,194,30,246,31,158,31,26,31,158,31,13,31,138,31,169,31,97,31,40,31,108,31,87,31,71,31,71,30,71,29,170,31,226,31,226,31,158,31,158,30,185,31,66,31,153,31,127,31,105,31,80,31,80,30,80,29,49,31,141,31,37,31,54,31,87,31,176,31,58,31,149,31,27,31,97,31,48,31,191,31,210,31,141,31,137,31,93,31,14,31,14,30,227,31,101,31,166,31,49,31,86,31,65,31,65,30,140,31,134,31,202,31,204,31,141,31,251,31,214,31,33,31,175,31,176,31,20,31,95,31,95,30,100,31,186,31,186,30,173,31,175,31,28,31,91,31,17,31,84,31,141,31,54,31,104,31,105,31,60,31,158,31,234,31,42,31,108,31,209,31,148,31,190,31,190,30,190,29,124,31,234,31,221,31,138,31,131,31,222,31,222,30,222,29,48,31,77,31,207,31,207,30,217,31,205,31,146,31,118,31,171,31,171,30,84,31,84,30,84,29,187,31,188,31,84,31,249,31,249,30,97,31,251,31,164,31,96,31,188,31,148,31,67,31,145,31,13,31,133,31,149,31,53,31,53,30,37,31,216,31,70,31,36,31,212,31,192,31,170,31,115,31,31,31,2,31,21,31,21,30,74,31,98,31,92,31,92,31,212,31,212,30,5,31,140,31,221,31,182,31,166,31,117,31,131,31,32,31,108,31,75,31,75,30,60,31,219,31,219,30,219,29,71,31,252,31,28,31,13,31,128,31,249,31,255,31,164,31,111,31,82,31,248,31,26,31,26,30,53,31,134,31,232,31,187,31,101,31,101,30,20,31,54,31,36,31,158,31,204,31,83,31,130,31,130,30,138,31,240,31,242,31,104,31,139,31,137,31,218,31,60,31,60,30,172,31,172,30,172,29,148,31,148,30,148,29,158,31,80,31,80,30,180,31,180,30,99,31,206,31,206,30,37,31,37,30,37,29,20,31,166,31,115,31,211,31,142,31,232,31,152,31,132,31,194,31,223,31,223,30,143,31,143,30,80,31,125,31,58,31,58,30,72,31,159,31,159,30,239,31,172,31,229,31,48,31,48,30,111,31,164,31,164,30,39,31,155,31,210,31,92,31,65,31,200,31,64,31,205,31,77,31,77,30,99,31,99,30,81,31,94,31,176,31,176,30,176,29,176,28,244,31,244,30,244,29,244,28,219,31,181,31,9,31,88,31,88,30,87,31,55,31,105,31,105,30,94,31,197,31,255,31,23,31,23,30,144,31,144,30,123,31,6,31,16,31,192,31,94,31,248,31,230,31,208,31,208,30,79,31,196,31,69,31,100,31,195,31,195,30,167,31,236,31,236,30,236,29,112,31,104,31,183,31,148,31,67,31,31,31,178,31,170,31,2,31,183,31,74,31,101,31,101,30,101,29,138,31,180,31,203,31,168,31,102,31,169,31,95,31,95,30,189,31,132,31,132,30,132,29,65,31,134,31,170,31,31,31,31,30,31,29,31,28,75,31,47,31,75,31,83,31,99,31,51,31,242,31,74,31,135,31,79,31,223,31,138,31,138,30,218,31,236,31,217,31,200,31,101,31,224,31,65,31,80,31,6,31,145,31,212,31,53,31,53,30,222,31,231,31,85,31,217,31,33,31,33,30,24,31,141,31,127,31,221,31,190,31,64,31,93,31,233,31,233,30,213,31,109,31,19,31,19,30,19,29,62,31,114,31,73,31,218,31,202,31,202,30,66,31,31,31,31,30,31,29,89,31,59,31,137,31,218,31,27,31,123,31,218,31,154,31,192,31,236,31,169,31,129,31,2,31,106,31,251,31,185,31,185,30,92,31,200,31,157,31,12,31,192,31,195,31,195,30,21,31,97,31,80,31,80,30,60,31,8,31,127,31,250,31,211,31,148,31,77,31,244,31,244,30,206,31,206,30,232,31,224,31,113,31,23,31,166,31,53,31,72,31,206,31,36,31,36,30,36,29,224,31,224,30,224,29,159,31,116,31,116,30,106,31,152,31,210,31,181,31,150,31,185,31,57,31,8,31,8,30,8,29,8,28,232,31,7,31,32,31,253,31,185,31,96,31,61,31,202,31,113,31,218,31,148,31,86,31,86,30,86,29,230,31,42,31,201,31,86,31,45,31,45,30,88,31,85,31,85,30,109,31,155,31,206,31,126,31,126,30,80,31,125,31,160,31,160,30,175,31,112,31,108,31,14,31,1,31,43,31,58,31,93,31,240,31,61,31,221,31,108,31,108,30,90,31,205,31,205,30,178,31,178,30,251,31,2,31,219,31,197,31,197,30,176,31,248,31,90,31,205,31,205,30,205,29,67,31,164,31,164,30,63,31,85,31,195,31,7,31,117,31,117,30,195,31,159,31,102,31,88,31,26,31,2,31,2,30,111,31,171,31,117,31,117,30,114,31,114,30,240,31,132,31,202,31,126,31,110,31,110,30,197,31,206,31,206,30,214,31,85,31,42,31,194,31,242,31,152,31,118,31,243,31,173,31,224,31,160,31,79,31,56,31,139,31,21,31,245,31,72,31,72,30,190,31,159,31,53,31,78,31,78,30,11,31,204,31,139,31,139,30,205,31,205,30,86,31,191,31,81,31,81,30,224,31,26,31,94,31,94,30,27,31,209,31,71,31,100,31,38,31,207,31,177,31,85,31,177,31,158,31,74,31,74,30,93,31,123,31,161,31,20,31,118,31,240,31,214,31,66,31,188,31,45,31,45,30,114,31,229,31,225,31,197,31,151,31,82,31,195,31,71,31,182,31,182,30,182,29,61,31,148,31,67,31,67,30,32,31,230,31,230,30,249,31,201,31,201,30,82,31,82,30,40,31,77,31,77,30,77,29,91,31,180,31,125,31,254,31,166,31,148,31,202,31,237,31,61,31,230,31,186,31,186,30,46,31,229,31,173,31,173,30,173,31,197,31,238,31,45,31,245,31,83,31,99,31,88,31,34,31,74,31,74,30,195,31,195,30,225,31,101,31,101,30,140,31,119,31,206,31,177,31,177,30,88,31,48,31,247,31,98,31,200,31,200,30,200,29,200,28,158,31,140,31,150,31,24,31,6,31,244,31,122,31,122,30,122,29,204,31,204,30,25,31,25,30,158,31,225,31,66,31,139,31,139,30,139,29,74,31,66,31,182,31,30,31,62,31,75,31,225,31,225,30,225,29,225,28);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
