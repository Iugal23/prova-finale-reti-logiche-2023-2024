-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_129 is
end project_tb_129;

architecture project_tb_arch_129 of project_tb_129 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 762;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,203,0,63,0,15,0,9,0,97,0,0,0,0,0,241,0,184,0,254,0,191,0,0,0,38,0,0,0,0,0,231,0,63,0,0,0,227,0,65,0,0,0,176,0,0,0,210,0,120,0,149,0,227,0,84,0,220,0,14,0,0,0,71,0,228,0,0,0,81,0,0,0,98,0,110,0,137,0,161,0,0,0,199,0,0,0,234,0,0,0,139,0,0,0,19,0,81,0,0,0,137,0,249,0,0,0,118,0,12,0,0,0,22,0,52,0,154,0,150,0,105,0,0,0,35,0,43,0,88,0,76,0,126,0,124,0,151,0,114,0,93,0,183,0,118,0,0,0,47,0,122,0,204,0,45,0,0,0,0,0,21,0,175,0,59,0,0,0,0,0,174,0,0,0,0,0,215,0,94,0,170,0,104,0,17,0,0,0,89,0,126,0,101,0,42,0,0,0,225,0,105,0,0,0,158,0,61,0,181,0,101,0,222,0,0,0,142,0,99,0,248,0,171,0,49,0,199,0,0,0,116,0,244,0,0,0,42,0,68,0,104,0,3,0,0,0,0,0,21,0,174,0,0,0,55,0,161,0,242,0,124,0,0,0,37,0,231,0,0,0,0,0,184,0,98,0,251,0,198,0,54,0,0,0,215,0,0,0,184,0,65,0,128,0,204,0,253,0,0,0,8,0,131,0,43,0,232,0,173,0,153,0,22,0,20,0,200,0,39,0,0,0,106,0,164,0,53,0,206,0,52,0,0,0,74,0,125,0,58,0,138,0,151,0,113,0,160,0,114,0,181,0,239,0,104,0,129,0,247,0,178,0,16,0,81,0,72,0,146,0,145,0,131,0,237,0,216,0,219,0,49,0,177,0,154,0,0,0,104,0,0,0,167,0,73,0,21,0,41,0,33,0,236,0,0,0,227,0,29,0,0,0,140,0,168,0,123,0,126,0,223,0,129,0,58,0,159,0,213,0,255,0,0,0,137,0,12,0,31,0,18,0,17,0,0,0,149,0,198,0,92,0,169,0,0,0,0,0,96,0,4,0,27,0,249,0,85,0,0,0,105,0,24,0,0,0,0,0,54,0,160,0,0,0,2,0,148,0,57,0,36,0,0,0,237,0,52,0,57,0,229,0,0,0,236,0,182,0,92,0,244,0,0,0,112,0,234,0,163,0,0,0,64,0,96,0,70,0,204,0,41,0,216,0,191,0,147,0,201,0,222,0,245,0,78,0,156,0,38,0,235,0,165,0,23,0,72,0,0,0,0,0,0,0,217,0,172,0,66,0,56,0,0,0,219,0,225,0,119,0,138,0,30,0,143,0,0,0,121,0,0,0,229,0,31,0,0,0,86,0,0,0,84,0,34,0,17,0,163,0,27,0,38,0,150,0,96,0,210,0,153,0,2,0,183,0,99,0,106,0,0,0,0,0,218,0,70,0,215,0,169,0,66,0,42,0,25,0,0,0,247,0,115,0,157,0,150,0,0,0,226,0,0,0,161,0,0,0,98,0,221,0,23,0,0,0,0,0,168,0,159,0,135,0,119,0,135,0,137,0,0,0,209,0,130,0,43,0,99,0,232,0,61,0,4,0,0,0,0,0,208,0,42,0,32,0,147,0,146,0,150,0,159,0,25,0,223,0,31,0,235,0,0,0,219,0,240,0,5,0,128,0,69,0,0,0,82,0,0,0,0,0,204,0,106,0,64,0,200,0,60,0,61,0,0,0,49,0,0,0,22,0,129,0,216,0,184,0,114,0,0,0,139,0,68,0,161,0,0,0,24,0,185,0,171,0,44,0,16,0,206,0,142,0,128,0,72,0,201,0,229,0,242,0,0,0,0,0,211,0,232,0,231,0,161,0,94,0,137,0,126,0,19,0,57,0,206,0,140,0,91,0,22,0,157,0,0,0,99,0,0,0,189,0,0,0,181,0,164,0,69,0,248,0,128,0,0,0,38,0,0,0,55,0,47,0,20,0,56,0,248,0,167,0,141,0,137,0,5,0,205,0,0,0,0,0,69,0,124,0,167,0,0,0,0,0,70,0,0,0,0,0,0,0,8,0,178,0,131,0,34,0,0,0,81,0,0,0,110,0,0,0,229,0,99,0,0,0,27,0,225,0,16,0,83,0,0,0,17,0,189,0,0,0,190,0,0,0,8,0,93,0,0,0,162,0,172,0,234,0,56,0,89,0,44,0,113,0,193,0,0,0,0,0,166,0,86,0,69,0,83,0,123,0,177,0,24,0,107,0,182,0,245,0,217,0,160,0,245,0,6,0,0,0,156,0,181,0,66,0,249,0,163,0,30,0,50,0,236,0,59,0,0,0,75,0,143,0,226,0,145,0,251,0,124,0,102,0,100,0,76,0,0,0,114,0,103,0,162,0,17,0,80,0,204,0,84,0,112,0,0,0,0,0,184,0,148,0,195,0,3,0,195,0,76,0,0,0,0,0,172,0,117,0,195,0,49,0,50,0,211,0,108,0,100,0,114,0,120,0,0,0,0,0,175,0,50,0,0,0,205,0,196,0,15,0,168,0,236,0,245,0,1,0,109,0,0,0,50,0,2,0,0,0,200,0,0,0,72,0,30,0,0,0,74,0,0,0,0,0,151,0,158,0,0,0,147,0,56,0,149,0,67,0,24,0,142,0,0,0,188,0,213,0,169,0,32,0,0,0,144,0,254,0,130,0,66,0,131,0,209,0,0,0,0,0,0,0,108,0,0,0,112,0,55,0,113,0,205,0,44,0,202,0,93,0,0,0,54,0,79,0,136,0,0,0,205,0,242,0,245,0,166,0,140,0,0,0,75,0,115,0,252,0,78,0,2,0,176,0,4,0,118,0,0,0,121,0,0,0,184,0,0,0,210,0,210,0,60,0,233,0,75,0,14,0,141,0,89,0,87,0,0,0,243,0,27,0,250,0,8,0,103,0,0,0,183,0,35,0,109,0,0,0,161,0,125,0,0,0,18,0,0,0,145,0,92,0,0,0,141,0,47,0,15,0,250,0,69,0,95,0,166,0,35,0,111,0,118,0,230,0,0,0,13,0,186,0,244,0,248,0,89,0,0,0,169,0,86,0,145,0,65,0,45,0,0,0,216,0,0,0,186,0,0,0,144,0,148,0,247,0,62,0,207,0,160,0,177,0,0,0,60,0,192,0,43,0,228,0,65,0,246,0,169,0,123,0,114,0,80,0,231,0,47,0,0,0,71,0,17,0,0,0,103,0,46,0,130,0,135,0,5,0,80,0,0,0,107,0,68,0,19,0,0,0,127,0,226,0,80,0,157,0,226,0,137,0,49,0,208,0,219,0,0,0,128,0,17,0,0,0,241,0,21,0,0,0,12,0,104,0,0,0,0,0,76,0,99,0,197,0,126,0,0,0,156,0,85,0,38,0,25,0,198,0,241,0,0,0,53,0);
signal scenario_full  : scenario_type := (0,0,203,31,63,31,15,31,9,31,97,31,97,30,97,29,241,31,184,31,254,31,191,31,191,30,38,31,38,30,38,29,231,31,63,31,63,30,227,31,65,31,65,30,176,31,176,30,210,31,120,31,149,31,227,31,84,31,220,31,14,31,14,30,71,31,228,31,228,30,81,31,81,30,98,31,110,31,137,31,161,31,161,30,199,31,199,30,234,31,234,30,139,31,139,30,19,31,81,31,81,30,137,31,249,31,249,30,118,31,12,31,12,30,22,31,52,31,154,31,150,31,105,31,105,30,35,31,43,31,88,31,76,31,126,31,124,31,151,31,114,31,93,31,183,31,118,31,118,30,47,31,122,31,204,31,45,31,45,30,45,29,21,31,175,31,59,31,59,30,59,29,174,31,174,30,174,29,215,31,94,31,170,31,104,31,17,31,17,30,89,31,126,31,101,31,42,31,42,30,225,31,105,31,105,30,158,31,61,31,181,31,101,31,222,31,222,30,142,31,99,31,248,31,171,31,49,31,199,31,199,30,116,31,244,31,244,30,42,31,68,31,104,31,3,31,3,30,3,29,21,31,174,31,174,30,55,31,161,31,242,31,124,31,124,30,37,31,231,31,231,30,231,29,184,31,98,31,251,31,198,31,54,31,54,30,215,31,215,30,184,31,65,31,128,31,204,31,253,31,253,30,8,31,131,31,43,31,232,31,173,31,153,31,22,31,20,31,200,31,39,31,39,30,106,31,164,31,53,31,206,31,52,31,52,30,74,31,125,31,58,31,138,31,151,31,113,31,160,31,114,31,181,31,239,31,104,31,129,31,247,31,178,31,16,31,81,31,72,31,146,31,145,31,131,31,237,31,216,31,219,31,49,31,177,31,154,31,154,30,104,31,104,30,167,31,73,31,21,31,41,31,33,31,236,31,236,30,227,31,29,31,29,30,140,31,168,31,123,31,126,31,223,31,129,31,58,31,159,31,213,31,255,31,255,30,137,31,12,31,31,31,18,31,17,31,17,30,149,31,198,31,92,31,169,31,169,30,169,29,96,31,4,31,27,31,249,31,85,31,85,30,105,31,24,31,24,30,24,29,54,31,160,31,160,30,2,31,148,31,57,31,36,31,36,30,237,31,52,31,57,31,229,31,229,30,236,31,182,31,92,31,244,31,244,30,112,31,234,31,163,31,163,30,64,31,96,31,70,31,204,31,41,31,216,31,191,31,147,31,201,31,222,31,245,31,78,31,156,31,38,31,235,31,165,31,23,31,72,31,72,30,72,29,72,28,217,31,172,31,66,31,56,31,56,30,219,31,225,31,119,31,138,31,30,31,143,31,143,30,121,31,121,30,229,31,31,31,31,30,86,31,86,30,84,31,34,31,17,31,163,31,27,31,38,31,150,31,96,31,210,31,153,31,2,31,183,31,99,31,106,31,106,30,106,29,218,31,70,31,215,31,169,31,66,31,42,31,25,31,25,30,247,31,115,31,157,31,150,31,150,30,226,31,226,30,161,31,161,30,98,31,221,31,23,31,23,30,23,29,168,31,159,31,135,31,119,31,135,31,137,31,137,30,209,31,130,31,43,31,99,31,232,31,61,31,4,31,4,30,4,29,208,31,42,31,32,31,147,31,146,31,150,31,159,31,25,31,223,31,31,31,235,31,235,30,219,31,240,31,5,31,128,31,69,31,69,30,82,31,82,30,82,29,204,31,106,31,64,31,200,31,60,31,61,31,61,30,49,31,49,30,22,31,129,31,216,31,184,31,114,31,114,30,139,31,68,31,161,31,161,30,24,31,185,31,171,31,44,31,16,31,206,31,142,31,128,31,72,31,201,31,229,31,242,31,242,30,242,29,211,31,232,31,231,31,161,31,94,31,137,31,126,31,19,31,57,31,206,31,140,31,91,31,22,31,157,31,157,30,99,31,99,30,189,31,189,30,181,31,164,31,69,31,248,31,128,31,128,30,38,31,38,30,55,31,47,31,20,31,56,31,248,31,167,31,141,31,137,31,5,31,205,31,205,30,205,29,69,31,124,31,167,31,167,30,167,29,70,31,70,30,70,29,70,28,8,31,178,31,131,31,34,31,34,30,81,31,81,30,110,31,110,30,229,31,99,31,99,30,27,31,225,31,16,31,83,31,83,30,17,31,189,31,189,30,190,31,190,30,8,31,93,31,93,30,162,31,172,31,234,31,56,31,89,31,44,31,113,31,193,31,193,30,193,29,166,31,86,31,69,31,83,31,123,31,177,31,24,31,107,31,182,31,245,31,217,31,160,31,245,31,6,31,6,30,156,31,181,31,66,31,249,31,163,31,30,31,50,31,236,31,59,31,59,30,75,31,143,31,226,31,145,31,251,31,124,31,102,31,100,31,76,31,76,30,114,31,103,31,162,31,17,31,80,31,204,31,84,31,112,31,112,30,112,29,184,31,148,31,195,31,3,31,195,31,76,31,76,30,76,29,172,31,117,31,195,31,49,31,50,31,211,31,108,31,100,31,114,31,120,31,120,30,120,29,175,31,50,31,50,30,205,31,196,31,15,31,168,31,236,31,245,31,1,31,109,31,109,30,50,31,2,31,2,30,200,31,200,30,72,31,30,31,30,30,74,31,74,30,74,29,151,31,158,31,158,30,147,31,56,31,149,31,67,31,24,31,142,31,142,30,188,31,213,31,169,31,32,31,32,30,144,31,254,31,130,31,66,31,131,31,209,31,209,30,209,29,209,28,108,31,108,30,112,31,55,31,113,31,205,31,44,31,202,31,93,31,93,30,54,31,79,31,136,31,136,30,205,31,242,31,245,31,166,31,140,31,140,30,75,31,115,31,252,31,78,31,2,31,176,31,4,31,118,31,118,30,121,31,121,30,184,31,184,30,210,31,210,31,60,31,233,31,75,31,14,31,141,31,89,31,87,31,87,30,243,31,27,31,250,31,8,31,103,31,103,30,183,31,35,31,109,31,109,30,161,31,125,31,125,30,18,31,18,30,145,31,92,31,92,30,141,31,47,31,15,31,250,31,69,31,95,31,166,31,35,31,111,31,118,31,230,31,230,30,13,31,186,31,244,31,248,31,89,31,89,30,169,31,86,31,145,31,65,31,45,31,45,30,216,31,216,30,186,31,186,30,144,31,148,31,247,31,62,31,207,31,160,31,177,31,177,30,60,31,192,31,43,31,228,31,65,31,246,31,169,31,123,31,114,31,80,31,231,31,47,31,47,30,71,31,17,31,17,30,103,31,46,31,130,31,135,31,5,31,80,31,80,30,107,31,68,31,19,31,19,30,127,31,226,31,80,31,157,31,226,31,137,31,49,31,208,31,219,31,219,30,128,31,17,31,17,30,241,31,21,31,21,30,12,31,104,31,104,30,104,29,76,31,99,31,197,31,126,31,126,30,156,31,85,31,38,31,25,31,198,31,241,31,241,30,53,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
