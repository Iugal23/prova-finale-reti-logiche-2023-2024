-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_333 is
end project_tb_333;

architecture project_tb_arch_333 of project_tb_333 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 856;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (109,0,255,0,133,0,0,0,53,0,44,0,71,0,0,0,149,0,231,0,215,0,0,0,236,0,53,0,169,0,0,0,0,0,20,0,116,0,0,0,0,0,50,0,209,0,0,0,246,0,0,0,0,0,187,0,218,0,135,0,229,0,231,0,0,0,113,0,78,0,0,0,151,0,147,0,0,0,228,0,0,0,123,0,0,0,0,0,0,0,0,0,19,0,141,0,0,0,192,0,0,0,52,0,28,0,240,0,171,0,133,0,106,0,244,0,33,0,190,0,109,0,201,0,30,0,91,0,18,0,245,0,174,0,0,0,222,0,10,0,19,0,162,0,175,0,156,0,249,0,203,0,44,0,234,0,0,0,0,0,25,0,211,0,3,0,0,0,98,0,115,0,206,0,30,0,207,0,40,0,204,0,124,0,67,0,59,0,114,0,0,0,76,0,165,0,84,0,234,0,0,0,156,0,102,0,119,0,0,0,233,0,145,0,123,0,54,0,146,0,0,0,253,0,0,0,50,0,53,0,135,0,144,0,0,0,0,0,0,0,0,0,12,0,0,0,192,0,108,0,111,0,37,0,57,0,96,0,58,0,111,0,255,0,135,0,0,0,72,0,70,0,0,0,239,0,169,0,170,0,0,0,104,0,202,0,166,0,4,0,32,0,121,0,131,0,139,0,9,0,54,0,0,0,164,0,82,0,0,0,93,0,120,0,0,0,179,0,217,0,59,0,254,0,234,0,57,0,139,0,181,0,0,0,65,0,0,0,151,0,6,0,142,0,5,0,17,0,0,0,206,0,220,0,0,0,113,0,213,0,144,0,89,0,225,0,64,0,177,0,142,0,0,0,145,0,159,0,196,0,231,0,167,0,118,0,186,0,143,0,97,0,136,0,177,0,115,0,0,0,0,0,36,0,37,0,208,0,12,0,23,0,47,0,92,0,0,0,253,0,227,0,0,0,111,0,56,0,56,0,67,0,156,0,0,0,2,0,103,0,77,0,0,0,79,0,166,0,73,0,0,0,84,0,188,0,70,0,180,0,52,0,221,0,62,0,0,0,41,0,135,0,73,0,153,0,36,0,148,0,164,0,240,0,145,0,101,0,236,0,85,0,0,0,31,0,100,0,224,0,47,0,0,0,146,0,0,0,0,0,169,0,210,0,130,0,129,0,0,0,43,0,229,0,157,0,62,0,0,0,97,0,0,0,55,0,65,0,162,0,142,0,0,0,44,0,0,0,81,0,0,0,117,0,195,0,0,0,0,0,20,0,68,0,0,0,38,0,62,0,121,0,242,0,0,0,0,0,0,0,179,0,230,0,178,0,167,0,86,0,162,0,170,0,52,0,10,0,0,0,202,0,216,0,55,0,178,0,60,0,62,0,244,0,232,0,35,0,0,0,248,0,196,0,0,0,116,0,76,0,54,0,12,0,134,0,153,0,108,0,196,0,109,0,232,0,0,0,40,0,88,0,122,0,109,0,189,0,58,0,238,0,180,0,143,0,248,0,38,0,221,0,15,0,120,0,193,0,0,0,159,0,81,0,161,0,0,0,0,0,117,0,174,0,11,0,145,0,12,0,0,0,0,0,217,0,19,0,0,0,0,0,101,0,114,0,127,0,0,0,56,0,89,0,0,0,0,0,106,0,174,0,138,0,21,0,228,0,89,0,67,0,0,0,40,0,0,0,0,0,240,0,167,0,0,0,131,0,0,0,0,0,159,0,98,0,0,0,0,0,154,0,101,0,32,0,83,0,0,0,0,0,218,0,0,0,140,0,156,0,154,0,11,0,204,0,95,0,0,0,0,0,173,0,24,0,44,0,109,0,155,0,0,0,104,0,9,0,0,0,27,0,160,0,203,0,0,0,74,0,58,0,164,0,6,0,199,0,132,0,0,0,6,0,128,0,195,0,7,0,58,0,197,0,0,0,200,0,145,0,60,0,52,0,32,0,0,0,0,0,43,0,6,0,130,0,92,0,154,0,0,0,231,0,238,0,129,0,129,0,90,0,151,0,159,0,73,0,232,0,0,0,14,0,153,0,237,0,51,0,22,0,0,0,210,0,247,0,196,0,0,0,234,0,0,0,71,0,218,0,106,0,171,0,0,0,97,0,63,0,244,0,166,0,29,0,226,0,0,0,0,0,58,0,161,0,99,0,198,0,35,0,0,0,159,0,44,0,101,0,0,0,204,0,0,0,0,0,58,0,116,0,0,0,191,0,88,0,33,0,232,0,62,0,245,0,126,0,125,0,25,0,158,0,154,0,0,0,31,0,5,0,199,0,199,0,67,0,160,0,132,0,96,0,231,0,109,0,0,0,0,0,123,0,115,0,33,0,0,0,0,0,101,0,221,0,116,0,0,0,184,0,70,0,128,0,86,0,53,0,254,0,0,0,5,0,140,0,106,0,72,0,28,0,70,0,230,0,194,0,138,0,0,0,129,0,248,0,163,0,85,0,160,0,0,0,121,0,121,0,204,0,53,0,76,0,86,0,212,0,80,0,251,0,125,0,58,0,233,0,0,0,152,0,164,0,58,0,190,0,0,0,0,0,0,0,122,0,210,0,40,0,114,0,169,0,104,0,170,0,247,0,0,0,88,0,24,0,0,0,0,0,0,0,199,0,226,0,178,0,83,0,84,0,0,0,0,0,34,0,0,0,133,0,201,0,35,0,186,0,82,0,129,0,1,0,0,0,246,0,165,0,146,0,7,0,245,0,112,0,30,0,140,0,0,0,17,0,0,0,45,0,78,0,57,0,157,0,86,0,134,0,213,0,57,0,8,0,66,0,0,0,0,0,220,0,186,0,167,0,157,0,169,0,99,0,249,0,114,0,233,0,144,0,0,0,0,0,146,0,235,0,75,0,237,0,243,0,122,0,0,0,0,0,4,0,0,0,62,0,105,0,197,0,246,0,0,0,44,0,229,0,249,0,31,0,27,0,0,0,14,0,190,0,16,0,0,0,87,0,0,0,79,0,123,0,0,0,160,0,54,0,11,0,227,0,0,0,111,0,144,0,145,0,190,0,130,0,23,0,67,0,82,0,209,0,163,0,86,0,190,0,190,0,0,0,186,0,145,0,144,0,0,0,113,0,23,0,164,0,0,0,64,0,234,0,123,0,18,0,145,0,25,0,92,0,112,0,5,0,0,0,155,0,178,0,63,0,243,0,16,0,131,0,195,0,164,0,143,0,60,0,5,0,146,0,46,0,181,0,248,0,133,0,117,0,0,0,210,0,243,0,71,0,78,0,47,0,80,0,0,0,217,0,47,0,60,0,194,0,220,0,0,0,2,0,193,0,214,0,93,0,141,0,109,0,217,0,6,0,210,0,0,0,0,0,216,0,191,0,243,0,0,0,66,0,139,0,83,0,104,0,135,0,220,0,16,0,178,0,0,0,4,0,6,0,241,0,0,0,0,0,231,0,167,0,79,0,142,0,237,0,0,0,0,0,34,0,134,0,130,0,67,0,0,0,201,0,54,0,191,0,44,0,0,0,28,0,241,0,0,0,46,0,169,0,226,0,64,0,252,0,5,0,0,0,158,0,86,0,189,0,98,0,52,0,92,0,82,0,26,0,1,0,75,0,48,0,218,0,83,0,125,0,0,0,110,0,0,0,111,0,67,0,252,0,0,0,0,0,0,0,0,0,112,0,165,0,28,0,6,0,0,0,167,0,189,0,100,0,141,0,34,0,1,0,116,0,0,0,164,0,177,0,55,0,0,0,33,0,92,0,44,0,101,0,163,0,193,0,153,0,136,0,100,0,206,0,228,0,0,0,19,0,222,0,37,0,159,0,0,0,237,0,0,0,214,0,147,0,0,0,238,0,96,0,0,0,20,0,0,0);
signal scenario_full  : scenario_type := (109,31,255,31,133,31,133,30,53,31,44,31,71,31,71,30,149,31,231,31,215,31,215,30,236,31,53,31,169,31,169,30,169,29,20,31,116,31,116,30,116,29,50,31,209,31,209,30,246,31,246,30,246,29,187,31,218,31,135,31,229,31,231,31,231,30,113,31,78,31,78,30,151,31,147,31,147,30,228,31,228,30,123,31,123,30,123,29,123,28,123,27,19,31,141,31,141,30,192,31,192,30,52,31,28,31,240,31,171,31,133,31,106,31,244,31,33,31,190,31,109,31,201,31,30,31,91,31,18,31,245,31,174,31,174,30,222,31,10,31,19,31,162,31,175,31,156,31,249,31,203,31,44,31,234,31,234,30,234,29,25,31,211,31,3,31,3,30,98,31,115,31,206,31,30,31,207,31,40,31,204,31,124,31,67,31,59,31,114,31,114,30,76,31,165,31,84,31,234,31,234,30,156,31,102,31,119,31,119,30,233,31,145,31,123,31,54,31,146,31,146,30,253,31,253,30,50,31,53,31,135,31,144,31,144,30,144,29,144,28,144,27,12,31,12,30,192,31,108,31,111,31,37,31,57,31,96,31,58,31,111,31,255,31,135,31,135,30,72,31,70,31,70,30,239,31,169,31,170,31,170,30,104,31,202,31,166,31,4,31,32,31,121,31,131,31,139,31,9,31,54,31,54,30,164,31,82,31,82,30,93,31,120,31,120,30,179,31,217,31,59,31,254,31,234,31,57,31,139,31,181,31,181,30,65,31,65,30,151,31,6,31,142,31,5,31,17,31,17,30,206,31,220,31,220,30,113,31,213,31,144,31,89,31,225,31,64,31,177,31,142,31,142,30,145,31,159,31,196,31,231,31,167,31,118,31,186,31,143,31,97,31,136,31,177,31,115,31,115,30,115,29,36,31,37,31,208,31,12,31,23,31,47,31,92,31,92,30,253,31,227,31,227,30,111,31,56,31,56,31,67,31,156,31,156,30,2,31,103,31,77,31,77,30,79,31,166,31,73,31,73,30,84,31,188,31,70,31,180,31,52,31,221,31,62,31,62,30,41,31,135,31,73,31,153,31,36,31,148,31,164,31,240,31,145,31,101,31,236,31,85,31,85,30,31,31,100,31,224,31,47,31,47,30,146,31,146,30,146,29,169,31,210,31,130,31,129,31,129,30,43,31,229,31,157,31,62,31,62,30,97,31,97,30,55,31,65,31,162,31,142,31,142,30,44,31,44,30,81,31,81,30,117,31,195,31,195,30,195,29,20,31,68,31,68,30,38,31,62,31,121,31,242,31,242,30,242,29,242,28,179,31,230,31,178,31,167,31,86,31,162,31,170,31,52,31,10,31,10,30,202,31,216,31,55,31,178,31,60,31,62,31,244,31,232,31,35,31,35,30,248,31,196,31,196,30,116,31,76,31,54,31,12,31,134,31,153,31,108,31,196,31,109,31,232,31,232,30,40,31,88,31,122,31,109,31,189,31,58,31,238,31,180,31,143,31,248,31,38,31,221,31,15,31,120,31,193,31,193,30,159,31,81,31,161,31,161,30,161,29,117,31,174,31,11,31,145,31,12,31,12,30,12,29,217,31,19,31,19,30,19,29,101,31,114,31,127,31,127,30,56,31,89,31,89,30,89,29,106,31,174,31,138,31,21,31,228,31,89,31,67,31,67,30,40,31,40,30,40,29,240,31,167,31,167,30,131,31,131,30,131,29,159,31,98,31,98,30,98,29,154,31,101,31,32,31,83,31,83,30,83,29,218,31,218,30,140,31,156,31,154,31,11,31,204,31,95,31,95,30,95,29,173,31,24,31,44,31,109,31,155,31,155,30,104,31,9,31,9,30,27,31,160,31,203,31,203,30,74,31,58,31,164,31,6,31,199,31,132,31,132,30,6,31,128,31,195,31,7,31,58,31,197,31,197,30,200,31,145,31,60,31,52,31,32,31,32,30,32,29,43,31,6,31,130,31,92,31,154,31,154,30,231,31,238,31,129,31,129,31,90,31,151,31,159,31,73,31,232,31,232,30,14,31,153,31,237,31,51,31,22,31,22,30,210,31,247,31,196,31,196,30,234,31,234,30,71,31,218,31,106,31,171,31,171,30,97,31,63,31,244,31,166,31,29,31,226,31,226,30,226,29,58,31,161,31,99,31,198,31,35,31,35,30,159,31,44,31,101,31,101,30,204,31,204,30,204,29,58,31,116,31,116,30,191,31,88,31,33,31,232,31,62,31,245,31,126,31,125,31,25,31,158,31,154,31,154,30,31,31,5,31,199,31,199,31,67,31,160,31,132,31,96,31,231,31,109,31,109,30,109,29,123,31,115,31,33,31,33,30,33,29,101,31,221,31,116,31,116,30,184,31,70,31,128,31,86,31,53,31,254,31,254,30,5,31,140,31,106,31,72,31,28,31,70,31,230,31,194,31,138,31,138,30,129,31,248,31,163,31,85,31,160,31,160,30,121,31,121,31,204,31,53,31,76,31,86,31,212,31,80,31,251,31,125,31,58,31,233,31,233,30,152,31,164,31,58,31,190,31,190,30,190,29,190,28,122,31,210,31,40,31,114,31,169,31,104,31,170,31,247,31,247,30,88,31,24,31,24,30,24,29,24,28,199,31,226,31,178,31,83,31,84,31,84,30,84,29,34,31,34,30,133,31,201,31,35,31,186,31,82,31,129,31,1,31,1,30,246,31,165,31,146,31,7,31,245,31,112,31,30,31,140,31,140,30,17,31,17,30,45,31,78,31,57,31,157,31,86,31,134,31,213,31,57,31,8,31,66,31,66,30,66,29,220,31,186,31,167,31,157,31,169,31,99,31,249,31,114,31,233,31,144,31,144,30,144,29,146,31,235,31,75,31,237,31,243,31,122,31,122,30,122,29,4,31,4,30,62,31,105,31,197,31,246,31,246,30,44,31,229,31,249,31,31,31,27,31,27,30,14,31,190,31,16,31,16,30,87,31,87,30,79,31,123,31,123,30,160,31,54,31,11,31,227,31,227,30,111,31,144,31,145,31,190,31,130,31,23,31,67,31,82,31,209,31,163,31,86,31,190,31,190,31,190,30,186,31,145,31,144,31,144,30,113,31,23,31,164,31,164,30,64,31,234,31,123,31,18,31,145,31,25,31,92,31,112,31,5,31,5,30,155,31,178,31,63,31,243,31,16,31,131,31,195,31,164,31,143,31,60,31,5,31,146,31,46,31,181,31,248,31,133,31,117,31,117,30,210,31,243,31,71,31,78,31,47,31,80,31,80,30,217,31,47,31,60,31,194,31,220,31,220,30,2,31,193,31,214,31,93,31,141,31,109,31,217,31,6,31,210,31,210,30,210,29,216,31,191,31,243,31,243,30,66,31,139,31,83,31,104,31,135,31,220,31,16,31,178,31,178,30,4,31,6,31,241,31,241,30,241,29,231,31,167,31,79,31,142,31,237,31,237,30,237,29,34,31,134,31,130,31,67,31,67,30,201,31,54,31,191,31,44,31,44,30,28,31,241,31,241,30,46,31,169,31,226,31,64,31,252,31,5,31,5,30,158,31,86,31,189,31,98,31,52,31,92,31,82,31,26,31,1,31,75,31,48,31,218,31,83,31,125,31,125,30,110,31,110,30,111,31,67,31,252,31,252,30,252,29,252,28,252,27,112,31,165,31,28,31,6,31,6,30,167,31,189,31,100,31,141,31,34,31,1,31,116,31,116,30,164,31,177,31,55,31,55,30,33,31,92,31,44,31,101,31,163,31,193,31,153,31,136,31,100,31,206,31,228,31,228,30,19,31,222,31,37,31,159,31,159,30,237,31,237,30,214,31,147,31,147,30,238,31,96,31,96,30,20,31,20,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
