-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_825 is
end project_tb_825;

architecture project_tb_arch_825 of project_tb_825 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 858;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (223,0,254,0,0,0,164,0,117,0,81,0,215,0,0,0,75,0,0,0,130,0,198,0,175,0,130,0,124,0,0,0,7,0,102,0,154,0,147,0,184,0,213,0,236,0,119,0,29,0,70,0,80,0,77,0,0,0,44,0,60,0,100,0,201,0,216,0,205,0,116,0,0,0,148,0,173,0,23,0,184,0,21,0,146,0,0,0,195,0,110,0,7,0,229,0,0,0,110,0,179,0,195,0,0,0,0,0,110,0,0,0,154,0,130,0,0,0,0,0,229,0,0,0,59,0,115,0,183,0,125,0,184,0,93,0,114,0,66,0,20,0,3,0,69,0,34,0,169,0,157,0,131,0,160,0,192,0,57,0,0,0,199,0,161,0,166,0,58,0,47,0,14,0,0,0,124,0,40,0,48,0,94,0,22,0,203,0,129,0,142,0,0,0,58,0,216,0,0,0,205,0,203,0,59,0,232,0,34,0,0,0,230,0,53,0,0,0,46,0,0,0,0,0,86,0,0,0,82,0,161,0,126,0,113,0,205,0,85,0,62,0,149,0,108,0,31,0,124,0,0,0,48,0,61,0,208,0,0,0,132,0,37,0,0,0,174,0,0,0,60,0,86,0,211,0,35,0,0,0,77,0,245,0,254,0,75,0,221,0,123,0,0,0,154,0,0,0,167,0,250,0,86,0,14,0,4,0,233,0,0,0,203,0,0,0,0,0,0,0,232,0,195,0,229,0,2,0,128,0,214,0,76,0,99,0,213,0,151,0,18,0,130,0,144,0,78,0,201,0,94,0,158,0,52,0,173,0,157,0,191,0,235,0,72,0,128,0,39,0,0,0,138,0,236,0,251,0,91,0,126,0,50,0,11,0,60,0,0,0,108,0,19,0,0,0,161,0,226,0,219,0,0,0,144,0,106,0,193,0,159,0,150,0,156,0,140,0,207,0,44,0,189,0,0,0,0,0,211,0,4,0,0,0,0,0,101,0,16,0,0,0,0,0,239,0,247,0,176,0,152,0,25,0,13,0,140,0,11,0,194,0,0,0,230,0,118,0,0,0,0,0,0,0,208,0,30,0,27,0,243,0,31,0,140,0,191,0,86,0,59,0,176,0,196,0,169,0,25,0,126,0,60,0,143,0,0,0,0,0,62,0,0,0,0,0,0,0,221,0,212,0,17,0,143,0,0,0,241,0,0,0,116,0,247,0,168,0,76,0,0,0,237,0,201,0,198,0,233,0,0,0,0,0,106,0,110,0,200,0,0,0,186,0,169,0,102,0,125,0,66,0,241,0,198,0,0,0,0,0,225,0,137,0,170,0,0,0,116,0,253,0,0,0,0,0,229,0,56,0,46,0,57,0,198,0,206,0,87,0,71,0,166,0,13,0,58,0,0,0,233,0,131,0,240,0,240,0,73,0,178,0,39,0,204,0,42,0,144,0,51,0,200,0,87,0,139,0,215,0,111,0,180,0,3,0,74,0,50,0,14,0,72,0,185,0,146,0,181,0,55,0,131,0,0,0,119,0,106,0,207,0,138,0,28,0,15,0,193,0,68,0,73,0,77,0,0,0,69,0,46,0,57,0,0,0,43,0,199,0,137,0,70,0,246,0,0,0,83,0,47,0,124,0,229,0,0,0,0,0,57,0,91,0,235,0,110,0,0,0,0,0,0,0,110,0,147,0,5,0,0,0,153,0,58,0,247,0,162,0,38,0,242,0,152,0,0,0,207,0,0,0,0,0,114,0,227,0,0,0,122,0,0,0,222,0,152,0,109,0,212,0,120,0,210,0,214,0,144,0,0,0,0,0,90,0,242,0,183,0,0,0,228,0,187,0,0,0,0,0,125,0,70,0,174,0,0,0,0,0,133,0,205,0,69,0,153,0,176,0,148,0,59,0,99,0,0,0,0,0,242,0,40,0,0,0,143,0,190,0,80,0,203,0,168,0,8,0,155,0,47,0,105,0,23,0,130,0,149,0,0,0,196,0,138,0,122,0,130,0,0,0,0,0,211,0,191,0,86,0,162,0,232,0,123,0,72,0,87,0,0,0,154,0,98,0,36,0,255,0,125,0,0,0,0,0,151,0,0,0,108,0,0,0,231,0,134,0,119,0,103,0,0,0,30,0,95,0,12,0,135,0,0,0,207,0,40,0,17,0,99,0,5,0,94,0,172,0,182,0,126,0,0,0,225,0,166,0,9,0,0,0,0,0,36,0,204,0,237,0,182,0,152,0,236,0,197,0,0,0,79,0,191,0,10,0,32,0,0,0,165,0,35,0,163,0,217,0,210,0,142,0,132,0,0,0,189,0,0,0,124,0,221,0,127,0,8,0,110,0,202,0,1,0,164,0,0,0,127,0,0,0,110,0,146,0,0,0,208,0,249,0,146,0,201,0,210,0,0,0,237,0,58,0,239,0,0,0,62,0,0,0,0,0,242,0,46,0,199,0,0,0,3,0,135,0,66,0,91,0,79,0,25,0,203,0,195,0,59,0,0,0,0,0,79,0,230,0,77,0,186,0,254,0,0,0,241,0,0,0,58,0,49,0,37,0,0,0,87,0,109,0,47,0,27,0,85,0,0,0,0,0,0,0,70,0,166,0,109,0,97,0,48,0,254,0,150,0,0,0,208,0,0,0,62,0,188,0,164,0,0,0,193,0,43,0,193,0,155,0,0,0,198,0,207,0,89,0,64,0,4,0,141,0,152,0,3,0,40,0,194,0,0,0,0,0,0,0,251,0,158,0,189,0,136,0,198,0,0,0,204,0,0,0,43,0,175,0,255,0,40,0,121,0,215,0,155,0,31,0,52,0,134,0,187,0,237,0,111,0,0,0,0,0,0,0,203,0,0,0,223,0,111,0,60,0,220,0,16,0,2,0,0,0,81,0,0,0,138,0,243,0,0,0,182,0,0,0,185,0,220,0,205,0,15,0,214,0,177,0,78,0,0,0,161,0,42,0,72,0,31,0,60,0,125,0,156,0,206,0,54,0,0,0,161,0,119,0,29,0,107,0,0,0,63,0,36,0,61,0,0,0,63,0,0,0,13,0,90,0,116,0,106,0,240,0,222,0,122,0,131,0,77,0,217,0,0,0,12,0,106,0,123,0,47,0,136,0,109,0,230,0,0,0,229,0,148,0,95,0,81,0,38,0,0,0,139,0,135,0,139,0,38,0,123,0,79,0,125,0,222,0,130,0,241,0,18,0,175,0,98,0,142,0,71,0,145,0,187,0,0,0,0,0,42,0,225,0,26,0,253,0,131,0,0,0,209,0,28,0,175,0,81,0,0,0,0,0,151,0,30,0,204,0,151,0,247,0,199,0,66,0,136,0,150,0,25,0,0,0,162,0,82,0,127,0,222,0,0,0,236,0,237,0,0,0,147,0,0,0,198,0,0,0,0,0,25,0,0,0,243,0,0,0,78,0,138,0,0,0,0,0,0,0,102,0,246,0,154,0,71,0,1,0,76,0,188,0,202,0,161,0,191,0,246,0,124,0,104,0,0,0,200,0,0,0,218,0,238,0,245,0,169,0,52,0,188,0,13,0,123,0,0,0,192,0,0,0,2,0,221,0,89,0,101,0,113,0,119,0,178,0,104,0,122,0,128,0,163,0,219,0,141,0,140,0,249,0,123,0,0,0,125,0,239,0,142,0,235,0,59,0,183,0,23,0,180,0,172,0,73,0,0,0,121,0,113,0,80,0,46,0,235,0,0,0,178,0,52,0,231,0,0,0,196,0,24,0,46,0,62,0,50,0,108,0,84,0,132,0,61,0,237,0,0,0,252,0,226,0,32,0,220,0,52,0,43,0,155,0,148,0,168,0,0,0,158,0,0,0,0,0,202,0,10,0);
signal scenario_full  : scenario_type := (223,31,254,31,254,30,164,31,117,31,81,31,215,31,215,30,75,31,75,30,130,31,198,31,175,31,130,31,124,31,124,30,7,31,102,31,154,31,147,31,184,31,213,31,236,31,119,31,29,31,70,31,80,31,77,31,77,30,44,31,60,31,100,31,201,31,216,31,205,31,116,31,116,30,148,31,173,31,23,31,184,31,21,31,146,31,146,30,195,31,110,31,7,31,229,31,229,30,110,31,179,31,195,31,195,30,195,29,110,31,110,30,154,31,130,31,130,30,130,29,229,31,229,30,59,31,115,31,183,31,125,31,184,31,93,31,114,31,66,31,20,31,3,31,69,31,34,31,169,31,157,31,131,31,160,31,192,31,57,31,57,30,199,31,161,31,166,31,58,31,47,31,14,31,14,30,124,31,40,31,48,31,94,31,22,31,203,31,129,31,142,31,142,30,58,31,216,31,216,30,205,31,203,31,59,31,232,31,34,31,34,30,230,31,53,31,53,30,46,31,46,30,46,29,86,31,86,30,82,31,161,31,126,31,113,31,205,31,85,31,62,31,149,31,108,31,31,31,124,31,124,30,48,31,61,31,208,31,208,30,132,31,37,31,37,30,174,31,174,30,60,31,86,31,211,31,35,31,35,30,77,31,245,31,254,31,75,31,221,31,123,31,123,30,154,31,154,30,167,31,250,31,86,31,14,31,4,31,233,31,233,30,203,31,203,30,203,29,203,28,232,31,195,31,229,31,2,31,128,31,214,31,76,31,99,31,213,31,151,31,18,31,130,31,144,31,78,31,201,31,94,31,158,31,52,31,173,31,157,31,191,31,235,31,72,31,128,31,39,31,39,30,138,31,236,31,251,31,91,31,126,31,50,31,11,31,60,31,60,30,108,31,19,31,19,30,161,31,226,31,219,31,219,30,144,31,106,31,193,31,159,31,150,31,156,31,140,31,207,31,44,31,189,31,189,30,189,29,211,31,4,31,4,30,4,29,101,31,16,31,16,30,16,29,239,31,247,31,176,31,152,31,25,31,13,31,140,31,11,31,194,31,194,30,230,31,118,31,118,30,118,29,118,28,208,31,30,31,27,31,243,31,31,31,140,31,191,31,86,31,59,31,176,31,196,31,169,31,25,31,126,31,60,31,143,31,143,30,143,29,62,31,62,30,62,29,62,28,221,31,212,31,17,31,143,31,143,30,241,31,241,30,116,31,247,31,168,31,76,31,76,30,237,31,201,31,198,31,233,31,233,30,233,29,106,31,110,31,200,31,200,30,186,31,169,31,102,31,125,31,66,31,241,31,198,31,198,30,198,29,225,31,137,31,170,31,170,30,116,31,253,31,253,30,253,29,229,31,56,31,46,31,57,31,198,31,206,31,87,31,71,31,166,31,13,31,58,31,58,30,233,31,131,31,240,31,240,31,73,31,178,31,39,31,204,31,42,31,144,31,51,31,200,31,87,31,139,31,215,31,111,31,180,31,3,31,74,31,50,31,14,31,72,31,185,31,146,31,181,31,55,31,131,31,131,30,119,31,106,31,207,31,138,31,28,31,15,31,193,31,68,31,73,31,77,31,77,30,69,31,46,31,57,31,57,30,43,31,199,31,137,31,70,31,246,31,246,30,83,31,47,31,124,31,229,31,229,30,229,29,57,31,91,31,235,31,110,31,110,30,110,29,110,28,110,31,147,31,5,31,5,30,153,31,58,31,247,31,162,31,38,31,242,31,152,31,152,30,207,31,207,30,207,29,114,31,227,31,227,30,122,31,122,30,222,31,152,31,109,31,212,31,120,31,210,31,214,31,144,31,144,30,144,29,90,31,242,31,183,31,183,30,228,31,187,31,187,30,187,29,125,31,70,31,174,31,174,30,174,29,133,31,205,31,69,31,153,31,176,31,148,31,59,31,99,31,99,30,99,29,242,31,40,31,40,30,143,31,190,31,80,31,203,31,168,31,8,31,155,31,47,31,105,31,23,31,130,31,149,31,149,30,196,31,138,31,122,31,130,31,130,30,130,29,211,31,191,31,86,31,162,31,232,31,123,31,72,31,87,31,87,30,154,31,98,31,36,31,255,31,125,31,125,30,125,29,151,31,151,30,108,31,108,30,231,31,134,31,119,31,103,31,103,30,30,31,95,31,12,31,135,31,135,30,207,31,40,31,17,31,99,31,5,31,94,31,172,31,182,31,126,31,126,30,225,31,166,31,9,31,9,30,9,29,36,31,204,31,237,31,182,31,152,31,236,31,197,31,197,30,79,31,191,31,10,31,32,31,32,30,165,31,35,31,163,31,217,31,210,31,142,31,132,31,132,30,189,31,189,30,124,31,221,31,127,31,8,31,110,31,202,31,1,31,164,31,164,30,127,31,127,30,110,31,146,31,146,30,208,31,249,31,146,31,201,31,210,31,210,30,237,31,58,31,239,31,239,30,62,31,62,30,62,29,242,31,46,31,199,31,199,30,3,31,135,31,66,31,91,31,79,31,25,31,203,31,195,31,59,31,59,30,59,29,79,31,230,31,77,31,186,31,254,31,254,30,241,31,241,30,58,31,49,31,37,31,37,30,87,31,109,31,47,31,27,31,85,31,85,30,85,29,85,28,70,31,166,31,109,31,97,31,48,31,254,31,150,31,150,30,208,31,208,30,62,31,188,31,164,31,164,30,193,31,43,31,193,31,155,31,155,30,198,31,207,31,89,31,64,31,4,31,141,31,152,31,3,31,40,31,194,31,194,30,194,29,194,28,251,31,158,31,189,31,136,31,198,31,198,30,204,31,204,30,43,31,175,31,255,31,40,31,121,31,215,31,155,31,31,31,52,31,134,31,187,31,237,31,111,31,111,30,111,29,111,28,203,31,203,30,223,31,111,31,60,31,220,31,16,31,2,31,2,30,81,31,81,30,138,31,243,31,243,30,182,31,182,30,185,31,220,31,205,31,15,31,214,31,177,31,78,31,78,30,161,31,42,31,72,31,31,31,60,31,125,31,156,31,206,31,54,31,54,30,161,31,119,31,29,31,107,31,107,30,63,31,36,31,61,31,61,30,63,31,63,30,13,31,90,31,116,31,106,31,240,31,222,31,122,31,131,31,77,31,217,31,217,30,12,31,106,31,123,31,47,31,136,31,109,31,230,31,230,30,229,31,148,31,95,31,81,31,38,31,38,30,139,31,135,31,139,31,38,31,123,31,79,31,125,31,222,31,130,31,241,31,18,31,175,31,98,31,142,31,71,31,145,31,187,31,187,30,187,29,42,31,225,31,26,31,253,31,131,31,131,30,209,31,28,31,175,31,81,31,81,30,81,29,151,31,30,31,204,31,151,31,247,31,199,31,66,31,136,31,150,31,25,31,25,30,162,31,82,31,127,31,222,31,222,30,236,31,237,31,237,30,147,31,147,30,198,31,198,30,198,29,25,31,25,30,243,31,243,30,78,31,138,31,138,30,138,29,138,28,102,31,246,31,154,31,71,31,1,31,76,31,188,31,202,31,161,31,191,31,246,31,124,31,104,31,104,30,200,31,200,30,218,31,238,31,245,31,169,31,52,31,188,31,13,31,123,31,123,30,192,31,192,30,2,31,221,31,89,31,101,31,113,31,119,31,178,31,104,31,122,31,128,31,163,31,219,31,141,31,140,31,249,31,123,31,123,30,125,31,239,31,142,31,235,31,59,31,183,31,23,31,180,31,172,31,73,31,73,30,121,31,113,31,80,31,46,31,235,31,235,30,178,31,52,31,231,31,231,30,196,31,24,31,46,31,62,31,50,31,108,31,84,31,132,31,61,31,237,31,237,30,252,31,226,31,32,31,220,31,52,31,43,31,155,31,148,31,168,31,168,30,158,31,158,30,158,29,202,31,10,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
