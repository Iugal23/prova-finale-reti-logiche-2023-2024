-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_904 is
end project_tb_904;

architecture project_tb_arch_904 of project_tb_904 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 247;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,29,0,0,0,106,0,127,0,23,0,8,0,0,0,145,0,195,0,193,0,200,0,190,0,75,0,71,0,0,0,177,0,253,0,157,0,132,0,7,0,0,0,38,0,0,0,253,0,240,0,128,0,0,0,83,0,128,0,156,0,138,0,138,0,83,0,218,0,222,0,0,0,0,0,31,0,217,0,204,0,83,0,247,0,148,0,170,0,232,0,197,0,195,0,108,0,0,0,209,0,204,0,0,0,63,0,195,0,180,0,48,0,250,0,93,0,239,0,103,0,239,0,31,0,67,0,52,0,199,0,224,0,34,0,10,0,37,0,0,0,116,0,96,0,0,0,21,0,89,0,18,0,42,0,17,0,183,0,0,0,248,0,46,0,107,0,150,0,114,0,133,0,76,0,83,0,27,0,179,0,48,0,114,0,200,0,0,0,0,0,198,0,204,0,219,0,2,0,0,0,0,0,194,0,35,0,107,0,222,0,205,0,99,0,116,0,89,0,0,0,51,0,231,0,159,0,92,0,107,0,0,0,0,0,0,0,194,0,0,0,104,0,204,0,87,0,0,0,118,0,205,0,197,0,66,0,251,0,0,0,80,0,216,0,0,0,113,0,0,0,196,0,49,0,124,0,39,0,153,0,149,0,128,0,249,0,119,0,110,0,62,0,14,0,22,0,97,0,26,0,89,0,0,0,0,0,120,0,49,0,141,0,123,0,146,0,205,0,20,0,157,0,139,0,174,0,246,0,0,0,202,0,89,0,40,0,204,0,130,0,101,0,184,0,198,0,16,0,216,0,146,0,159,0,0,0,105,0,134,0,145,0,170,0,198,0,0,0,125,0,213,0,0,0,112,0,32,0,118,0,0,0,224,0,30,0,47,0,58,0,0,0,197,0,170,0,0,0,222,0,117,0,87,0,0,0,127,0,49,0,130,0,78,0,0,0,19,0,199,0,13,0,0,0,118,0,221,0,94,0,67,0,66,0,188,0,228,0,48,0,0,0,194,0,0,0,3,0,168,0,166,0,0,0,0,0,130,0,150,0,0,0,104,0,68,0,64,0,229,0,223,0,0,0,212,0,56,0,0,0,136,0,54,0,0,0,67,0,241,0,0,0);
signal scenario_full  : scenario_type := (0,0,29,31,29,30,106,31,127,31,23,31,8,31,8,30,145,31,195,31,193,31,200,31,190,31,75,31,71,31,71,30,177,31,253,31,157,31,132,31,7,31,7,30,38,31,38,30,253,31,240,31,128,31,128,30,83,31,128,31,156,31,138,31,138,31,83,31,218,31,222,31,222,30,222,29,31,31,217,31,204,31,83,31,247,31,148,31,170,31,232,31,197,31,195,31,108,31,108,30,209,31,204,31,204,30,63,31,195,31,180,31,48,31,250,31,93,31,239,31,103,31,239,31,31,31,67,31,52,31,199,31,224,31,34,31,10,31,37,31,37,30,116,31,96,31,96,30,21,31,89,31,18,31,42,31,17,31,183,31,183,30,248,31,46,31,107,31,150,31,114,31,133,31,76,31,83,31,27,31,179,31,48,31,114,31,200,31,200,30,200,29,198,31,204,31,219,31,2,31,2,30,2,29,194,31,35,31,107,31,222,31,205,31,99,31,116,31,89,31,89,30,51,31,231,31,159,31,92,31,107,31,107,30,107,29,107,28,194,31,194,30,104,31,204,31,87,31,87,30,118,31,205,31,197,31,66,31,251,31,251,30,80,31,216,31,216,30,113,31,113,30,196,31,49,31,124,31,39,31,153,31,149,31,128,31,249,31,119,31,110,31,62,31,14,31,22,31,97,31,26,31,89,31,89,30,89,29,120,31,49,31,141,31,123,31,146,31,205,31,20,31,157,31,139,31,174,31,246,31,246,30,202,31,89,31,40,31,204,31,130,31,101,31,184,31,198,31,16,31,216,31,146,31,159,31,159,30,105,31,134,31,145,31,170,31,198,31,198,30,125,31,213,31,213,30,112,31,32,31,118,31,118,30,224,31,30,31,47,31,58,31,58,30,197,31,170,31,170,30,222,31,117,31,87,31,87,30,127,31,49,31,130,31,78,31,78,30,19,31,199,31,13,31,13,30,118,31,221,31,94,31,67,31,66,31,188,31,228,31,48,31,48,30,194,31,194,30,3,31,168,31,166,31,166,30,166,29,130,31,150,31,150,30,104,31,68,31,64,31,229,31,223,31,223,30,212,31,56,31,56,30,136,31,54,31,54,30,67,31,241,31,241,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
