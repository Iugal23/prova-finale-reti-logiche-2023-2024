-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_774 is
end project_tb_774;

architecture project_tb_arch_774 of project_tb_774 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 750;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,29,0,134,0,170,0,81,0,0,0,199,0,8,0,135,0,149,0,254,0,28,0,16,0,0,0,24,0,0,0,216,0,149,0,129,0,129,0,0,0,128,0,0,0,20,0,0,0,177,0,76,0,52,0,74,0,118,0,144,0,138,0,0,0,120,0,192,0,192,0,209,0,193,0,236,0,61,0,142,0,207,0,0,0,234,0,152,0,121,0,0,0,0,0,0,0,0,0,0,0,69,0,241,0,78,0,156,0,164,0,204,0,165,0,172,0,169,0,138,0,2,0,129,0,195,0,212,0,13,0,164,0,137,0,71,0,126,0,225,0,189,0,228,0,203,0,215,0,0,0,98,0,54,0,0,0,185,0,76,0,0,0,26,0,242,0,233,0,195,0,171,0,77,0,89,0,49,0,130,0,226,0,84,0,0,0,32,0,137,0,222,0,209,0,197,0,102,0,2,0,240,0,0,0,0,0,58,0,205,0,60,0,177,0,74,0,109,0,153,0,77,0,178,0,242,0,39,0,146,0,159,0,96,0,115,0,90,0,0,0,55,0,140,0,6,0,86,0,39,0,237,0,0,0,120,0,0,0,59,0,0,0,50,0,58,0,35,0,0,0,0,0,224,0,0,0,86,0,157,0,0,0,0,0,102,0,39,0,0,0,169,0,165,0,45,0,229,0,48,0,27,0,0,0,0,0,0,0,71,0,136,0,250,0,0,0,54,0,98,0,46,0,0,0,0,0,122,0,145,0,108,0,16,0,75,0,227,0,35,0,59,0,11,0,0,0,0,0,0,0,216,0,0,0,0,0,38,0,70,0,0,0,0,0,45,0,184,0,77,0,43,0,0,0,228,0,134,0,168,0,209,0,0,0,112,0,0,0,29,0,82,0,210,0,166,0,0,0,60,0,0,0,16,0,18,0,37,0,173,0,0,0,212,0,0,0,200,0,0,0,0,0,130,0,0,0,183,0,206,0,0,0,229,0,188,0,29,0,35,0,156,0,167,0,112,0,52,0,133,0,178,0,38,0,138,0,246,0,10,0,67,0,0,0,4,0,64,0,103,0,189,0,144,0,14,0,67,0,0,0,193,0,0,0,48,0,100,0,0,0,0,0,64,0,0,0,0,0,51,0,0,0,73,0,101,0,0,0,186,0,59,0,205,0,85,0,0,0,183,0,225,0,57,0,73,0,192,0,161,0,144,0,42,0,207,0,0,0,0,0,0,0,46,0,121,0,209,0,0,0,95,0,231,0,42,0,64,0,0,0,0,0,188,0,81,0,92,0,64,0,87,0,247,0,52,0,127,0,189,0,158,0,37,0,254,0,120,0,160,0,48,0,124,0,47,0,249,0,232,0,243,0,196,0,62,0,127,0,49,0,23,0,53,0,12,0,210,0,28,0,5,0,110,0,0,0,233,0,1,0,101,0,1,0,232,0,165,0,127,0,37,0,83,0,13,0,250,0,0,0,46,0,147,0,197,0,81,0,194,0,0,0,9,0,68,0,0,0,0,0,0,0,209,0,0,0,10,0,38,0,63,0,211,0,17,0,252,0,2,0,242,0,0,0,136,0,57,0,247,0,79,0,237,0,249,0,180,0,9,0,161,0,48,0,42,0,72,0,132,0,54,0,220,0,31,0,172,0,253,0,0,0,243,0,197,0,195,0,57,0,182,0,236,0,0,0,27,0,169,0,61,0,0,0,127,0,126,0,0,0,245,0,22,0,0,0,195,0,0,0,46,0,178,0,130,0,11,0,171,0,146,0,248,0,178,0,117,0,5,0,143,0,60,0,0,0,0,0,97,0,18,0,248,0,1,0,226,0,0,0,56,0,183,0,221,0,230,0,22,0,162,0,48,0,142,0,87,0,0,0,0,0,135,0,180,0,0,0,15,0,164,0,12,0,110,0,166,0,206,0,114,0,37,0,206,0,0,0,172,0,116,0,184,0,33,0,218,0,156,0,212,0,54,0,34,0,0,0,125,0,152,0,0,0,166,0,0,0,18,0,187,0,0,0,253,0,251,0,129,0,77,0,121,0,0,0,11,0,0,0,47,0,237,0,20,0,0,0,95,0,0,0,233,0,72,0,51,0,118,0,250,0,197,0,213,0,124,0,58,0,204,0,198,0,78,0,118,0,54,0,0,0,104,0,51,0,0,0,13,0,194,0,0,0,61,0,180,0,0,0,126,0,94,0,160,0,0,0,118,0,0,0,149,0,0,0,175,0,132,0,169,0,62,0,0,0,215,0,0,0,191,0,205,0,122,0,80,0,0,0,164,0,115,0,234,0,0,0,22,0,153,0,240,0,240,0,156,0,135,0,122,0,204,0,168,0,149,0,88,0,245,0,0,0,127,0,224,0,164,0,78,0,0,0,249,0,0,0,23,0,165,0,253,0,131,0,0,0,129,0,142,0,217,0,210,0,0,0,0,0,223,0,0,0,133,0,184,0,65,0,19,0,169,0,170,0,66,0,23,0,31,0,232,0,93,0,2,0,143,0,196,0,7,0,213,0,0,0,0,0,0,0,21,0,54,0,194,0,76,0,151,0,228,0,37,0,213,0,26,0,53,0,116,0,206,0,39,0,98,0,50,0,131,0,147,0,94,0,243,0,0,0,252,0,193,0,210,0,48,0,184,0,71,0,19,0,180,0,219,0,93,0,66,0,158,0,177,0,33,0,91,0,34,0,0,0,0,0,51,0,0,0,185,0,71,0,245,0,178,0,139,0,0,0,0,0,0,0,203,0,0,0,192,0,0,0,135,0,79,0,254,0,0,0,101,0,57,0,136,0,0,0,189,0,209,0,146,0,117,0,28,0,109,0,110,0,0,0,93,0,167,0,15,0,107,0,0,0,90,0,137,0,0,0,159,0,123,0,83,0,133,0,206,0,171,0,0,0,0,0,245,0,56,0,207,0,108,0,202,0,240,0,94,0,172,0,151,0,17,0,0,0,165,0,28,0,0,0,0,0,53,0,108,0,41,0,156,0,239,0,13,0,73,0,157,0,245,0,93,0,245,0,0,0,76,0,0,0,42,0,123,0,0,0,132,0,225,0,0,0,0,0,45,0,33,0,188,0,25,0,64,0,0,0,17,0,252,0,128,0,0,0,248,0,61,0,41,0,188,0,198,0,108,0,0,0,101,0,222,0,132,0,201,0,16,0,138,0,121,0,0,0,219,0,85,0,0,0,64,0,146,0,200,0,36,0,50,0,0,0,185,0,114,0,208,0,251,0,0,0,21,0,202,0,73,0,155,0,0,0,215,0,69,0,0,0,251,0,60,0,120,0,179,0,205,0,222,0,111,0,193,0,226,0,0,0,4,0,0,0,0,0,230,0,0,0,0,0,189,0,20,0,34,0,0,0,121,0);
signal scenario_full  : scenario_type := (0,0,29,31,134,31,170,31,81,31,81,30,199,31,8,31,135,31,149,31,254,31,28,31,16,31,16,30,24,31,24,30,216,31,149,31,129,31,129,31,129,30,128,31,128,30,20,31,20,30,177,31,76,31,52,31,74,31,118,31,144,31,138,31,138,30,120,31,192,31,192,31,209,31,193,31,236,31,61,31,142,31,207,31,207,30,234,31,152,31,121,31,121,30,121,29,121,28,121,27,121,26,69,31,241,31,78,31,156,31,164,31,204,31,165,31,172,31,169,31,138,31,2,31,129,31,195,31,212,31,13,31,164,31,137,31,71,31,126,31,225,31,189,31,228,31,203,31,215,31,215,30,98,31,54,31,54,30,185,31,76,31,76,30,26,31,242,31,233,31,195,31,171,31,77,31,89,31,49,31,130,31,226,31,84,31,84,30,32,31,137,31,222,31,209,31,197,31,102,31,2,31,240,31,240,30,240,29,58,31,205,31,60,31,177,31,74,31,109,31,153,31,77,31,178,31,242,31,39,31,146,31,159,31,96,31,115,31,90,31,90,30,55,31,140,31,6,31,86,31,39,31,237,31,237,30,120,31,120,30,59,31,59,30,50,31,58,31,35,31,35,30,35,29,224,31,224,30,86,31,157,31,157,30,157,29,102,31,39,31,39,30,169,31,165,31,45,31,229,31,48,31,27,31,27,30,27,29,27,28,71,31,136,31,250,31,250,30,54,31,98,31,46,31,46,30,46,29,122,31,145,31,108,31,16,31,75,31,227,31,35,31,59,31,11,31,11,30,11,29,11,28,216,31,216,30,216,29,38,31,70,31,70,30,70,29,45,31,184,31,77,31,43,31,43,30,228,31,134,31,168,31,209,31,209,30,112,31,112,30,29,31,82,31,210,31,166,31,166,30,60,31,60,30,16,31,18,31,37,31,173,31,173,30,212,31,212,30,200,31,200,30,200,29,130,31,130,30,183,31,206,31,206,30,229,31,188,31,29,31,35,31,156,31,167,31,112,31,52,31,133,31,178,31,38,31,138,31,246,31,10,31,67,31,67,30,4,31,64,31,103,31,189,31,144,31,14,31,67,31,67,30,193,31,193,30,48,31,100,31,100,30,100,29,64,31,64,30,64,29,51,31,51,30,73,31,101,31,101,30,186,31,59,31,205,31,85,31,85,30,183,31,225,31,57,31,73,31,192,31,161,31,144,31,42,31,207,31,207,30,207,29,207,28,46,31,121,31,209,31,209,30,95,31,231,31,42,31,64,31,64,30,64,29,188,31,81,31,92,31,64,31,87,31,247,31,52,31,127,31,189,31,158,31,37,31,254,31,120,31,160,31,48,31,124,31,47,31,249,31,232,31,243,31,196,31,62,31,127,31,49,31,23,31,53,31,12,31,210,31,28,31,5,31,110,31,110,30,233,31,1,31,101,31,1,31,232,31,165,31,127,31,37,31,83,31,13,31,250,31,250,30,46,31,147,31,197,31,81,31,194,31,194,30,9,31,68,31,68,30,68,29,68,28,209,31,209,30,10,31,38,31,63,31,211,31,17,31,252,31,2,31,242,31,242,30,136,31,57,31,247,31,79,31,237,31,249,31,180,31,9,31,161,31,48,31,42,31,72,31,132,31,54,31,220,31,31,31,172,31,253,31,253,30,243,31,197,31,195,31,57,31,182,31,236,31,236,30,27,31,169,31,61,31,61,30,127,31,126,31,126,30,245,31,22,31,22,30,195,31,195,30,46,31,178,31,130,31,11,31,171,31,146,31,248,31,178,31,117,31,5,31,143,31,60,31,60,30,60,29,97,31,18,31,248,31,1,31,226,31,226,30,56,31,183,31,221,31,230,31,22,31,162,31,48,31,142,31,87,31,87,30,87,29,135,31,180,31,180,30,15,31,164,31,12,31,110,31,166,31,206,31,114,31,37,31,206,31,206,30,172,31,116,31,184,31,33,31,218,31,156,31,212,31,54,31,34,31,34,30,125,31,152,31,152,30,166,31,166,30,18,31,187,31,187,30,253,31,251,31,129,31,77,31,121,31,121,30,11,31,11,30,47,31,237,31,20,31,20,30,95,31,95,30,233,31,72,31,51,31,118,31,250,31,197,31,213,31,124,31,58,31,204,31,198,31,78,31,118,31,54,31,54,30,104,31,51,31,51,30,13,31,194,31,194,30,61,31,180,31,180,30,126,31,94,31,160,31,160,30,118,31,118,30,149,31,149,30,175,31,132,31,169,31,62,31,62,30,215,31,215,30,191,31,205,31,122,31,80,31,80,30,164,31,115,31,234,31,234,30,22,31,153,31,240,31,240,31,156,31,135,31,122,31,204,31,168,31,149,31,88,31,245,31,245,30,127,31,224,31,164,31,78,31,78,30,249,31,249,30,23,31,165,31,253,31,131,31,131,30,129,31,142,31,217,31,210,31,210,30,210,29,223,31,223,30,133,31,184,31,65,31,19,31,169,31,170,31,66,31,23,31,31,31,232,31,93,31,2,31,143,31,196,31,7,31,213,31,213,30,213,29,213,28,21,31,54,31,194,31,76,31,151,31,228,31,37,31,213,31,26,31,53,31,116,31,206,31,39,31,98,31,50,31,131,31,147,31,94,31,243,31,243,30,252,31,193,31,210,31,48,31,184,31,71,31,19,31,180,31,219,31,93,31,66,31,158,31,177,31,33,31,91,31,34,31,34,30,34,29,51,31,51,30,185,31,71,31,245,31,178,31,139,31,139,30,139,29,139,28,203,31,203,30,192,31,192,30,135,31,79,31,254,31,254,30,101,31,57,31,136,31,136,30,189,31,209,31,146,31,117,31,28,31,109,31,110,31,110,30,93,31,167,31,15,31,107,31,107,30,90,31,137,31,137,30,159,31,123,31,83,31,133,31,206,31,171,31,171,30,171,29,245,31,56,31,207,31,108,31,202,31,240,31,94,31,172,31,151,31,17,31,17,30,165,31,28,31,28,30,28,29,53,31,108,31,41,31,156,31,239,31,13,31,73,31,157,31,245,31,93,31,245,31,245,30,76,31,76,30,42,31,123,31,123,30,132,31,225,31,225,30,225,29,45,31,33,31,188,31,25,31,64,31,64,30,17,31,252,31,128,31,128,30,248,31,61,31,41,31,188,31,198,31,108,31,108,30,101,31,222,31,132,31,201,31,16,31,138,31,121,31,121,30,219,31,85,31,85,30,64,31,146,31,200,31,36,31,50,31,50,30,185,31,114,31,208,31,251,31,251,30,21,31,202,31,73,31,155,31,155,30,215,31,69,31,69,30,251,31,60,31,120,31,179,31,205,31,222,31,111,31,193,31,226,31,226,30,4,31,4,30,4,29,230,31,230,30,230,29,189,31,20,31,34,31,34,30,121,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
