-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 407;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,31,0,32,0,0,0,201,0,174,0,211,0,101,0,6,0,224,0,148,0,0,0,48,0,25,0,10,0,217,0,208,0,0,0,128,0,179,0,0,0,138,0,189,0,242,0,207,0,113,0,157,0,0,0,39,0,71,0,51,0,215,0,155,0,119,0,94,0,54,0,13,0,0,0,27,0,0,0,151,0,93,0,0,0,104,0,85,0,132,0,32,0,86,0,54,0,0,0,0,0,68,0,213,0,222,0,78,0,87,0,216,0,84,0,107,0,100,0,0,0,128,0,9,0,0,0,96,0,0,0,2,0,0,0,171,0,181,0,93,0,0,0,74,0,102,0,49,0,213,0,249,0,0,0,5,0,236,0,121,0,29,0,165,0,121,0,210,0,122,0,252,0,0,0,118,0,11,0,23,0,232,0,16,0,244,0,141,0,245,0,212,0,96,0,115,0,27,0,119,0,196,0,112,0,180,0,66,0,169,0,175,0,116,0,0,0,131,0,173,0,115,0,253,0,19,0,106,0,246,0,145,0,206,0,179,0,0,0,29,0,0,0,73,0,168,0,37,0,149,0,0,0,152,0,12,0,37,0,0,0,2,0,103,0,178,0,0,0,112,0,0,0,15,0,0,0,0,0,0,0,30,0,0,0,0,0,36,0,0,0,132,0,119,0,96,0,243,0,121,0,204,0,24,0,149,0,250,0,167,0,68,0,0,0,152,0,118,0,163,0,42,0,75,0,154,0,155,0,10,0,0,0,23,0,176,0,194,0,235,0,0,0,0,0,241,0,0,0,67,0,99,0,231,0,0,0,0,0,34,0,186,0,222,0,176,0,6,0,128,0,23,0,139,0,0,0,219,0,74,0,157,0,109,0,167,0,148,0,143,0,85,0,21,0,208,0,54,0,104,0,228,0,63,0,39,0,230,0,163,0,145,0,246,0,51,0,0,0,0,0,68,0,103,0,32,0,51,0,166,0,62,0,92,0,26,0,50,0,85,0,85,0,190,0,251,0,0,0,75,0,97,0,209,0,0,0,0,0,179,0,209,0,10,0,213,0,165,0,12,0,194,0,50,0,160,0,172,0,204,0,0,0,244,0,239,0,74,0,0,0,0,0,41,0,114,0,0,0,8,0,247,0,60,0,17,0,95,0,132,0,0,0,0,0,53,0,130,0,182,0,199,0,19,0,0,0,8,0,128,0,0,0,0,0,68,0,253,0,30,0,4,0,0,0,208,0,192,0,161,0,40,0,0,0,249,0,6,0,47,0,246,0,59,0,190,0,152,0,111,0,0,0,0,0,0,0,234,0,197,0,0,0,45,0,0,0,253,0,26,0,63,0,254,0,0,0,174,0,51,0,250,0,83,0,182,0,62,0,111,0,125,0,191,0,75,0,68,0,23,0,199,0,215,0,181,0,3,0,0,0,0,0,117,0,44,0,31,0,35,0,207,0,0,0,199,0,0,0,0,0,188,0,202,0,0,0,0,0,0,0,69,0,11,0,18,0,117,0,148,0,253,0,217,0,211,0,14,0,161,0,16,0,56,0,191,0,0,0,18,0,180,0,175,0,0,0,209,0,183,0,0,0,35,0,0,0,0,0,0,0,0,0,4,0,220,0,18,0,0,0,247,0,245,0,161,0,121,0,4,0,10,0,196,0,196,0,0,0,13,0,130,0,25,0,225,0,0,0,26,0,166,0,0,0,165,0,0,0,0,0,124,0,134,0,159,0,0,0,32,0,137,0,222,0,83,0,95,0,213,0,6,0,170,0,129,0,147,0,3,0,246,0,42,0,0,0,214,0,53,0,0,0,8,0,3,0,31,0,176,0,106,0);
signal scenario_full  : scenario_type := (0,0,31,31,32,31,32,30,201,31,174,31,211,31,101,31,6,31,224,31,148,31,148,30,48,31,25,31,10,31,217,31,208,31,208,30,128,31,179,31,179,30,138,31,189,31,242,31,207,31,113,31,157,31,157,30,39,31,71,31,51,31,215,31,155,31,119,31,94,31,54,31,13,31,13,30,27,31,27,30,151,31,93,31,93,30,104,31,85,31,132,31,32,31,86,31,54,31,54,30,54,29,68,31,213,31,222,31,78,31,87,31,216,31,84,31,107,31,100,31,100,30,128,31,9,31,9,30,96,31,96,30,2,31,2,30,171,31,181,31,93,31,93,30,74,31,102,31,49,31,213,31,249,31,249,30,5,31,236,31,121,31,29,31,165,31,121,31,210,31,122,31,252,31,252,30,118,31,11,31,23,31,232,31,16,31,244,31,141,31,245,31,212,31,96,31,115,31,27,31,119,31,196,31,112,31,180,31,66,31,169,31,175,31,116,31,116,30,131,31,173,31,115,31,253,31,19,31,106,31,246,31,145,31,206,31,179,31,179,30,29,31,29,30,73,31,168,31,37,31,149,31,149,30,152,31,12,31,37,31,37,30,2,31,103,31,178,31,178,30,112,31,112,30,15,31,15,30,15,29,15,28,30,31,30,30,30,29,36,31,36,30,132,31,119,31,96,31,243,31,121,31,204,31,24,31,149,31,250,31,167,31,68,31,68,30,152,31,118,31,163,31,42,31,75,31,154,31,155,31,10,31,10,30,23,31,176,31,194,31,235,31,235,30,235,29,241,31,241,30,67,31,99,31,231,31,231,30,231,29,34,31,186,31,222,31,176,31,6,31,128,31,23,31,139,31,139,30,219,31,74,31,157,31,109,31,167,31,148,31,143,31,85,31,21,31,208,31,54,31,104,31,228,31,63,31,39,31,230,31,163,31,145,31,246,31,51,31,51,30,51,29,68,31,103,31,32,31,51,31,166,31,62,31,92,31,26,31,50,31,85,31,85,31,190,31,251,31,251,30,75,31,97,31,209,31,209,30,209,29,179,31,209,31,10,31,213,31,165,31,12,31,194,31,50,31,160,31,172,31,204,31,204,30,244,31,239,31,74,31,74,30,74,29,41,31,114,31,114,30,8,31,247,31,60,31,17,31,95,31,132,31,132,30,132,29,53,31,130,31,182,31,199,31,19,31,19,30,8,31,128,31,128,30,128,29,68,31,253,31,30,31,4,31,4,30,208,31,192,31,161,31,40,31,40,30,249,31,6,31,47,31,246,31,59,31,190,31,152,31,111,31,111,30,111,29,111,28,234,31,197,31,197,30,45,31,45,30,253,31,26,31,63,31,254,31,254,30,174,31,51,31,250,31,83,31,182,31,62,31,111,31,125,31,191,31,75,31,68,31,23,31,199,31,215,31,181,31,3,31,3,30,3,29,117,31,44,31,31,31,35,31,207,31,207,30,199,31,199,30,199,29,188,31,202,31,202,30,202,29,202,28,69,31,11,31,18,31,117,31,148,31,253,31,217,31,211,31,14,31,161,31,16,31,56,31,191,31,191,30,18,31,180,31,175,31,175,30,209,31,183,31,183,30,35,31,35,30,35,29,35,28,35,27,4,31,220,31,18,31,18,30,247,31,245,31,161,31,121,31,4,31,10,31,196,31,196,31,196,30,13,31,130,31,25,31,225,31,225,30,26,31,166,31,166,30,165,31,165,30,165,29,124,31,134,31,159,31,159,30,32,31,137,31,222,31,83,31,95,31,213,31,6,31,170,31,129,31,147,31,3,31,246,31,42,31,42,30,214,31,53,31,53,30,8,31,3,31,31,31,176,31,106,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
