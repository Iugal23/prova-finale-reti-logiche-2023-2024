-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 699;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (169,0,0,0,91,0,73,0,58,0,187,0,0,0,156,0,188,0,248,0,0,0,93,0,228,0,124,0,4,0,64,0,0,0,0,0,15,0,92,0,194,0,8,0,63,0,0,0,28,0,17,0,181,0,16,0,227,0,162,0,117,0,16,0,196,0,82,0,46,0,132,0,186,0,175,0,173,0,0,0,205,0,230,0,0,0,86,0,100,0,247,0,240,0,115,0,0,0,0,0,0,0,209,0,78,0,247,0,177,0,91,0,191,0,227,0,52,0,177,0,3,0,17,0,16,0,0,0,156,0,117,0,144,0,40,0,130,0,129,0,127,0,138,0,162,0,49,0,49,0,39,0,136,0,116,0,0,0,51,0,138,0,189,0,87,0,0,0,106,0,180,0,229,0,0,0,0,0,0,0,0,0,59,0,76,0,78,0,79,0,0,0,0,0,147,0,188,0,181,0,0,0,197,0,93,0,145,0,75,0,0,0,0,0,0,0,119,0,5,0,13,0,21,0,62,0,185,0,125,0,0,0,4,0,61,0,93,0,235,0,19,0,234,0,0,0,58,0,0,0,29,0,228,0,105,0,231,0,75,0,186,0,53,0,190,0,90,0,121,0,0,0,52,0,0,0,165,0,181,0,232,0,0,0,95,0,119,0,0,0,0,0,32,0,9,0,85,0,239,0,214,0,184,0,137,0,0,0,75,0,0,0,142,0,206,0,0,0,0,0,10,0,0,0,183,0,46,0,0,0,184,0,223,0,198,0,0,0,0,0,0,0,201,0,117,0,0,0,253,0,204,0,88,0,112,0,238,0,0,0,219,0,10,0,182,0,26,0,0,0,68,0,121,0,165,0,33,0,56,0,255,0,92,0,134,0,25,0,22,0,0,0,234,0,149,0,239,0,91,0,235,0,229,0,60,0,143,0,182,0,0,0,73,0,77,0,136,0,148,0,194,0,44,0,185,0,211,0,49,0,44,0,201,0,0,0,118,0,149,0,0,0,250,0,18,0,0,0,125,0,230,0,93,0,135,0,50,0,95,0,83,0,0,0,13,0,72,0,16,0,171,0,204,0,0,0,85,0,17,0,204,0,232,0,0,0,103,0,1,0,40,0,118,0,236,0,0,0,228,0,71,0,149,0,217,0,63,0,65,0,0,0,186,0,29,0,0,0,98,0,0,0,7,0,202,0,0,0,97,0,0,0,58,0,226,0,184,0,76,0,144,0,0,0,24,0,190,0,0,0,210,0,113,0,194,0,46,0,157,0,168,0,9,0,134,0,100,0,193,0,8,0,44,0,0,0,94,0,103,0,187,0,137,0,0,0,0,0,28,0,116,0,198,0,0,0,0,0,159,0,12,0,147,0,69,0,174,0,0,0,0,0,2,0,36,0,0,0,105,0,135,0,0,0,81,0,97,0,163,0,0,0,68,0,87,0,96,0,40,0,56,0,78,0,126,0,196,0,158,0,0,0,23,0,59,0,199,0,219,0,0,0,247,0,26,0,127,0,207,0,0,0,240,0,245,0,130,0,160,0,31,0,6,0,18,0,115,0,0,0,31,0,72,0,69,0,7,0,223,0,197,0,192,0,200,0,181,0,227,0,7,0,0,0,163,0,209,0,248,0,0,0,33,0,132,0,220,0,134,0,251,0,39,0,227,0,0,0,0,0,175,0,61,0,116,0,188,0,149,0,73,0,136,0,179,0,213,0,0,0,17,0,0,0,180,0,232,0,9,0,60,0,87,0,84,0,227,0,0,0,0,0,60,0,223,0,115,0,104,0,161,0,0,0,11,0,138,0,31,0,211,0,0,0,0,0,169,0,130,0,66,0,204,0,0,0,110,0,202,0,160,0,0,0,205,0,212,0,60,0,54,0,227,0,229,0,22,0,33,0,0,0,67,0,115,0,0,0,26,0,0,0,136,0,213,0,3,0,169,0,65,0,67,0,100,0,0,0,0,0,164,0,0,0,190,0,252,0,173,0,219,0,37,0,7,0,232,0,108,0,78,0,0,0,70,0,61,0,205,0,75,0,183,0,179,0,0,0,176,0,236,0,173,0,233,0,229,0,217,0,175,0,221,0,49,0,0,0,135,0,0,0,185,0,201,0,133,0,65,0,146,0,210,0,236,0,0,0,0,0,249,0,91,0,72,0,152,0,97,0,199,0,125,0,246,0,234,0,0,0,208,0,117,0,86,0,137,0,173,0,164,0,59,0,0,0,250,0,237,0,0,0,71,0,193,0,57,0,62,0,0,0,131,0,48,0,252,0,199,0,2,0,28,0,113,0,189,0,50,0,22,0,138,0,115,0,182,0,213,0,63,0,105,0,205,0,247,0,11,0,0,0,81,0,245,0,91,0,83,0,117,0,0,0,82,0,189,0,102,0,47,0,168,0,135,0,98,0,188,0,251,0,177,0,0,0,43,0,152,0,0,0,110,0,0,0,78,0,165,0,189,0,19,0,217,0,92,0,106,0,123,0,61,0,0,0,113,0,26,0,74,0,0,0,40,0,110,0,13,0,71,0,49,0,0,0,247,0,169,0,0,0,77,0,121,0,227,0,0,0,207,0,177,0,200,0,232,0,177,0,58,0,17,0,97,0,197,0,28,0,0,0,18,0,155,0,220,0,148,0,96,0,240,0,15,0,199,0,42,0,0,0,210,0,223,0,83,0,0,0,133,0,127,0,127,0,238,0,119,0,55,0,149,0,3,0,242,0,82,0,104,0,81,0,40,0,250,0,0,0,46,0,239,0,73,0,185,0,184,0,3,0,218,0,96,0,253,0,137,0,184,0,213,0,0,0,0,0,0,0,232,0,201,0,0,0,62,0,164,0,169,0,229,0,164,0,132,0,217,0,221,0,16,0,126,0,0,0,135,0,182,0,133,0,45,0,115,0,0,0,4,0,0,0,28,0,238,0,46,0,51,0,108,0,173,0,121,0,149,0,0,0,57,0,0,0,230,0,214,0,206,0,0,0,115,0,172,0,203,0,0,0,212,0,97,0,131,0,0,0,0,0,150,0,255,0,88,0,193,0,174,0,194,0,131,0,213,0,155,0,208,0,26,0,0,0,246,0,163,0,28,0,192,0,69,0,242,0,0,0,0,0,217,0,8,0,220,0,53,0,221,0,0,0,170,0,0,0);
signal scenario_full  : scenario_type := (169,31,169,30,91,31,73,31,58,31,187,31,187,30,156,31,188,31,248,31,248,30,93,31,228,31,124,31,4,31,64,31,64,30,64,29,15,31,92,31,194,31,8,31,63,31,63,30,28,31,17,31,181,31,16,31,227,31,162,31,117,31,16,31,196,31,82,31,46,31,132,31,186,31,175,31,173,31,173,30,205,31,230,31,230,30,86,31,100,31,247,31,240,31,115,31,115,30,115,29,115,28,209,31,78,31,247,31,177,31,91,31,191,31,227,31,52,31,177,31,3,31,17,31,16,31,16,30,156,31,117,31,144,31,40,31,130,31,129,31,127,31,138,31,162,31,49,31,49,31,39,31,136,31,116,31,116,30,51,31,138,31,189,31,87,31,87,30,106,31,180,31,229,31,229,30,229,29,229,28,229,27,59,31,76,31,78,31,79,31,79,30,79,29,147,31,188,31,181,31,181,30,197,31,93,31,145,31,75,31,75,30,75,29,75,28,119,31,5,31,13,31,21,31,62,31,185,31,125,31,125,30,4,31,61,31,93,31,235,31,19,31,234,31,234,30,58,31,58,30,29,31,228,31,105,31,231,31,75,31,186,31,53,31,190,31,90,31,121,31,121,30,52,31,52,30,165,31,181,31,232,31,232,30,95,31,119,31,119,30,119,29,32,31,9,31,85,31,239,31,214,31,184,31,137,31,137,30,75,31,75,30,142,31,206,31,206,30,206,29,10,31,10,30,183,31,46,31,46,30,184,31,223,31,198,31,198,30,198,29,198,28,201,31,117,31,117,30,253,31,204,31,88,31,112,31,238,31,238,30,219,31,10,31,182,31,26,31,26,30,68,31,121,31,165,31,33,31,56,31,255,31,92,31,134,31,25,31,22,31,22,30,234,31,149,31,239,31,91,31,235,31,229,31,60,31,143,31,182,31,182,30,73,31,77,31,136,31,148,31,194,31,44,31,185,31,211,31,49,31,44,31,201,31,201,30,118,31,149,31,149,30,250,31,18,31,18,30,125,31,230,31,93,31,135,31,50,31,95,31,83,31,83,30,13,31,72,31,16,31,171,31,204,31,204,30,85,31,17,31,204,31,232,31,232,30,103,31,1,31,40,31,118,31,236,31,236,30,228,31,71,31,149,31,217,31,63,31,65,31,65,30,186,31,29,31,29,30,98,31,98,30,7,31,202,31,202,30,97,31,97,30,58,31,226,31,184,31,76,31,144,31,144,30,24,31,190,31,190,30,210,31,113,31,194,31,46,31,157,31,168,31,9,31,134,31,100,31,193,31,8,31,44,31,44,30,94,31,103,31,187,31,137,31,137,30,137,29,28,31,116,31,198,31,198,30,198,29,159,31,12,31,147,31,69,31,174,31,174,30,174,29,2,31,36,31,36,30,105,31,135,31,135,30,81,31,97,31,163,31,163,30,68,31,87,31,96,31,40,31,56,31,78,31,126,31,196,31,158,31,158,30,23,31,59,31,199,31,219,31,219,30,247,31,26,31,127,31,207,31,207,30,240,31,245,31,130,31,160,31,31,31,6,31,18,31,115,31,115,30,31,31,72,31,69,31,7,31,223,31,197,31,192,31,200,31,181,31,227,31,7,31,7,30,163,31,209,31,248,31,248,30,33,31,132,31,220,31,134,31,251,31,39,31,227,31,227,30,227,29,175,31,61,31,116,31,188,31,149,31,73,31,136,31,179,31,213,31,213,30,17,31,17,30,180,31,232,31,9,31,60,31,87,31,84,31,227,31,227,30,227,29,60,31,223,31,115,31,104,31,161,31,161,30,11,31,138,31,31,31,211,31,211,30,211,29,169,31,130,31,66,31,204,31,204,30,110,31,202,31,160,31,160,30,205,31,212,31,60,31,54,31,227,31,229,31,22,31,33,31,33,30,67,31,115,31,115,30,26,31,26,30,136,31,213,31,3,31,169,31,65,31,67,31,100,31,100,30,100,29,164,31,164,30,190,31,252,31,173,31,219,31,37,31,7,31,232,31,108,31,78,31,78,30,70,31,61,31,205,31,75,31,183,31,179,31,179,30,176,31,236,31,173,31,233,31,229,31,217,31,175,31,221,31,49,31,49,30,135,31,135,30,185,31,201,31,133,31,65,31,146,31,210,31,236,31,236,30,236,29,249,31,91,31,72,31,152,31,97,31,199,31,125,31,246,31,234,31,234,30,208,31,117,31,86,31,137,31,173,31,164,31,59,31,59,30,250,31,237,31,237,30,71,31,193,31,57,31,62,31,62,30,131,31,48,31,252,31,199,31,2,31,28,31,113,31,189,31,50,31,22,31,138,31,115,31,182,31,213,31,63,31,105,31,205,31,247,31,11,31,11,30,81,31,245,31,91,31,83,31,117,31,117,30,82,31,189,31,102,31,47,31,168,31,135,31,98,31,188,31,251,31,177,31,177,30,43,31,152,31,152,30,110,31,110,30,78,31,165,31,189,31,19,31,217,31,92,31,106,31,123,31,61,31,61,30,113,31,26,31,74,31,74,30,40,31,110,31,13,31,71,31,49,31,49,30,247,31,169,31,169,30,77,31,121,31,227,31,227,30,207,31,177,31,200,31,232,31,177,31,58,31,17,31,97,31,197,31,28,31,28,30,18,31,155,31,220,31,148,31,96,31,240,31,15,31,199,31,42,31,42,30,210,31,223,31,83,31,83,30,133,31,127,31,127,31,238,31,119,31,55,31,149,31,3,31,242,31,82,31,104,31,81,31,40,31,250,31,250,30,46,31,239,31,73,31,185,31,184,31,3,31,218,31,96,31,253,31,137,31,184,31,213,31,213,30,213,29,213,28,232,31,201,31,201,30,62,31,164,31,169,31,229,31,164,31,132,31,217,31,221,31,16,31,126,31,126,30,135,31,182,31,133,31,45,31,115,31,115,30,4,31,4,30,28,31,238,31,46,31,51,31,108,31,173,31,121,31,149,31,149,30,57,31,57,30,230,31,214,31,206,31,206,30,115,31,172,31,203,31,203,30,212,31,97,31,131,31,131,30,131,29,150,31,255,31,88,31,193,31,174,31,194,31,131,31,213,31,155,31,208,31,26,31,26,30,246,31,163,31,28,31,192,31,69,31,242,31,242,30,242,29,217,31,8,31,220,31,53,31,221,31,221,30,170,31,170,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
