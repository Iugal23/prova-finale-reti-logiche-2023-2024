-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 614;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,136,0,0,0,62,0,223,0,0,0,0,0,90,0,33,0,88,0,117,0,234,0,122,0,140,0,40,0,6,0,233,0,60,0,244,0,203,0,121,0,44,0,0,0,128,0,250,0,44,0,30,0,0,0,154,0,84,0,226,0,219,0,187,0,209,0,6,0,176,0,161,0,57,0,146,0,196,0,219,0,117,0,98,0,230,0,208,0,228,0,57,0,182,0,86,0,0,0,36,0,10,0,0,0,37,0,226,0,213,0,246,0,18,0,203,0,0,0,155,0,98,0,65,0,17,0,0,0,162,0,141,0,242,0,118,0,0,0,0,0,0,0,234,0,0,0,114,0,197,0,120,0,124,0,39,0,91,0,110,0,128,0,251,0,0,0,101,0,204,0,173,0,251,0,165,0,233,0,30,0,45,0,43,0,0,0,177,0,87,0,88,0,201,0,168,0,0,0,34,0,0,0,189,0,2,0,0,0,92,0,0,0,0,0,93,0,247,0,170,0,226,0,237,0,75,0,0,0,232,0,175,0,32,0,199,0,213,0,47,0,210,0,52,0,13,0,20,0,88,0,0,0,42,0,46,0,138,0,97,0,6,0,223,0,175,0,100,0,46,0,29,0,51,0,16,0,0,0,110,0,109,0,91,0,216,0,80,0,0,0,39,0,0,0,89,0,0,0,90,0,111,0,207,0,0,0,0,0,48,0,132,0,0,0,0,0,0,0,105,0,227,0,246,0,0,0,47,0,84,0,0,0,0,0,182,0,248,0,221,0,148,0,243,0,250,0,0,0,169,0,98,0,169,0,121,0,53,0,87,0,0,0,109,0,0,0,161,0,46,0,0,0,0,0,175,0,34,0,228,0,33,0,7,0,28,0,0,0,125,0,91,0,192,0,239,0,0,0,206,0,0,0,139,0,138,0,14,0,183,0,119,0,164,0,211,0,173,0,90,0,44,0,43,0,6,0,3,0,162,0,198,0,122,0,88,0,0,0,41,0,110,0,0,0,245,0,105,0,0,0,130,0,15,0,66,0,135,0,154,0,0,0,138,0,0,0,51,0,76,0,94,0,25,0,0,0,81,0,15,0,236,0,167,0,66,0,82,0,0,0,213,0,255,0,104,0,0,0,78,0,72,0,170,0,146,0,0,0,230,0,10,0,0,0,0,0,124,0,0,0,0,0,0,0,222,0,178,0,202,0,0,0,230,0,199,0,0,0,0,0,51,0,24,0,55,0,0,0,0,0,0,0,88,0,8,0,212,0,11,0,170,0,155,0,167,0,162,0,96,0,154,0,235,0,0,0,8,0,13,0,125,0,129,0,209,0,0,0,128,0,208,0,0,0,0,0,0,0,85,0,100,0,0,0,133,0,161,0,107,0,161,0,221,0,0,0,140,0,154,0,0,0,48,0,207,0,186,0,103,0,70,0,0,0,31,0,66,0,214,0,202,0,226,0,96,0,106,0,85,0,121,0,200,0,43,0,30,0,137,0,182,0,4,0,0,0,30,0,31,0,77,0,119,0,154,0,35,0,113,0,0,0,157,0,187,0,191,0,0,0,0,0,203,0,202,0,249,0,41,0,59,0,215,0,152,0,151,0,163,0,98,0,46,0,244,0,29,0,254,0,23,0,122,0,0,0,173,0,117,0,158,0,43,0,190,0,27,0,0,0,164,0,149,0,223,0,183,0,103,0,63,0,122,0,27,0,0,0,63,0,160,0,177,0,27,0,63,0,182,0,0,0,160,0,0,0,232,0,222,0,63,0,51,0,0,0,217,0,24,0,128,0,243,0,97,0,23,0,88,0,0,0,105,0,99,0,198,0,0,0,187,0,8,0,0,0,254,0,216,0,191,0,168,0,0,0,8,0,227,0,0,0,249,0,116,0,0,0,254,0,102,0,153,0,97,0,0,0,150,0,14,0,202,0,80,0,5,0,181,0,55,0,5,0,1,0,0,0,68,0,0,0,195,0,0,0,142,0,196,0,22,0,0,0,0,0,9,0,42,0,20,0,140,0,128,0,17,0,0,0,10,0,52,0,191,0,69,0,0,0,37,0,122,0,0,0,193,0,106,0,0,0,241,0,229,0,122,0,4,0,167,0,252,0,107,0,142,0,173,0,0,0,137,0,232,0,0,0,31,0,186,0,114,0,8,0,0,0,174,0,226,0,0,0,0,0,174,0,156,0,0,0,158,0,24,0,103,0,13,0,202,0,10,0,76,0,5,0,0,0,73,0,19,0,204,0,195,0,190,0,186,0,108,0,231,0,109,0,0,0,0,0,148,0,66,0,0,0,230,0,206,0,66,0,104,0,0,0,125,0,247,0,107,0,166,0,125,0,42,0,178,0,36,0,180,0,230,0,137,0,0,0,157,0,162,0,103,0,5,0,212,0,199,0,227,0,30,0,59,0,0,0,28,0,26,0,11,0,24,0,153,0,45,0,182,0,0,0,0,0,210,0,33,0,67,0,0,0,165,0,70,0,0,0,228,0,60,0,235,0,216,0,225,0,0,0,51,0,46,0,193,0,59,0,167,0,204,0,4,0,179,0,142,0,110,0,243,0,116,0,18,0,0,0,79,0,118,0,105,0,0,0,19,0,171,0,0,0,0,0,94,0,147,0,254,0,247,0,0,0,121,0,146,0,220,0,150,0,250,0,220,0,201,0,0,0,116,0,81,0,105,0,66,0,121,0,1,0,70,0,0,0,218,0,204,0,5,0,196,0,91,0,233,0,255,0,0,0,119,0,255,0,134,0,149,0);
signal scenario_full  : scenario_type := (0,0,136,31,136,30,62,31,223,31,223,30,223,29,90,31,33,31,88,31,117,31,234,31,122,31,140,31,40,31,6,31,233,31,60,31,244,31,203,31,121,31,44,31,44,30,128,31,250,31,44,31,30,31,30,30,154,31,84,31,226,31,219,31,187,31,209,31,6,31,176,31,161,31,57,31,146,31,196,31,219,31,117,31,98,31,230,31,208,31,228,31,57,31,182,31,86,31,86,30,36,31,10,31,10,30,37,31,226,31,213,31,246,31,18,31,203,31,203,30,155,31,98,31,65,31,17,31,17,30,162,31,141,31,242,31,118,31,118,30,118,29,118,28,234,31,234,30,114,31,197,31,120,31,124,31,39,31,91,31,110,31,128,31,251,31,251,30,101,31,204,31,173,31,251,31,165,31,233,31,30,31,45,31,43,31,43,30,177,31,87,31,88,31,201,31,168,31,168,30,34,31,34,30,189,31,2,31,2,30,92,31,92,30,92,29,93,31,247,31,170,31,226,31,237,31,75,31,75,30,232,31,175,31,32,31,199,31,213,31,47,31,210,31,52,31,13,31,20,31,88,31,88,30,42,31,46,31,138,31,97,31,6,31,223,31,175,31,100,31,46,31,29,31,51,31,16,31,16,30,110,31,109,31,91,31,216,31,80,31,80,30,39,31,39,30,89,31,89,30,90,31,111,31,207,31,207,30,207,29,48,31,132,31,132,30,132,29,132,28,105,31,227,31,246,31,246,30,47,31,84,31,84,30,84,29,182,31,248,31,221,31,148,31,243,31,250,31,250,30,169,31,98,31,169,31,121,31,53,31,87,31,87,30,109,31,109,30,161,31,46,31,46,30,46,29,175,31,34,31,228,31,33,31,7,31,28,31,28,30,125,31,91,31,192,31,239,31,239,30,206,31,206,30,139,31,138,31,14,31,183,31,119,31,164,31,211,31,173,31,90,31,44,31,43,31,6,31,3,31,162,31,198,31,122,31,88,31,88,30,41,31,110,31,110,30,245,31,105,31,105,30,130,31,15,31,66,31,135,31,154,31,154,30,138,31,138,30,51,31,76,31,94,31,25,31,25,30,81,31,15,31,236,31,167,31,66,31,82,31,82,30,213,31,255,31,104,31,104,30,78,31,72,31,170,31,146,31,146,30,230,31,10,31,10,30,10,29,124,31,124,30,124,29,124,28,222,31,178,31,202,31,202,30,230,31,199,31,199,30,199,29,51,31,24,31,55,31,55,30,55,29,55,28,88,31,8,31,212,31,11,31,170,31,155,31,167,31,162,31,96,31,154,31,235,31,235,30,8,31,13,31,125,31,129,31,209,31,209,30,128,31,208,31,208,30,208,29,208,28,85,31,100,31,100,30,133,31,161,31,107,31,161,31,221,31,221,30,140,31,154,31,154,30,48,31,207,31,186,31,103,31,70,31,70,30,31,31,66,31,214,31,202,31,226,31,96,31,106,31,85,31,121,31,200,31,43,31,30,31,137,31,182,31,4,31,4,30,30,31,31,31,77,31,119,31,154,31,35,31,113,31,113,30,157,31,187,31,191,31,191,30,191,29,203,31,202,31,249,31,41,31,59,31,215,31,152,31,151,31,163,31,98,31,46,31,244,31,29,31,254,31,23,31,122,31,122,30,173,31,117,31,158,31,43,31,190,31,27,31,27,30,164,31,149,31,223,31,183,31,103,31,63,31,122,31,27,31,27,30,63,31,160,31,177,31,27,31,63,31,182,31,182,30,160,31,160,30,232,31,222,31,63,31,51,31,51,30,217,31,24,31,128,31,243,31,97,31,23,31,88,31,88,30,105,31,99,31,198,31,198,30,187,31,8,31,8,30,254,31,216,31,191,31,168,31,168,30,8,31,227,31,227,30,249,31,116,31,116,30,254,31,102,31,153,31,97,31,97,30,150,31,14,31,202,31,80,31,5,31,181,31,55,31,5,31,1,31,1,30,68,31,68,30,195,31,195,30,142,31,196,31,22,31,22,30,22,29,9,31,42,31,20,31,140,31,128,31,17,31,17,30,10,31,52,31,191,31,69,31,69,30,37,31,122,31,122,30,193,31,106,31,106,30,241,31,229,31,122,31,4,31,167,31,252,31,107,31,142,31,173,31,173,30,137,31,232,31,232,30,31,31,186,31,114,31,8,31,8,30,174,31,226,31,226,30,226,29,174,31,156,31,156,30,158,31,24,31,103,31,13,31,202,31,10,31,76,31,5,31,5,30,73,31,19,31,204,31,195,31,190,31,186,31,108,31,231,31,109,31,109,30,109,29,148,31,66,31,66,30,230,31,206,31,66,31,104,31,104,30,125,31,247,31,107,31,166,31,125,31,42,31,178,31,36,31,180,31,230,31,137,31,137,30,157,31,162,31,103,31,5,31,212,31,199,31,227,31,30,31,59,31,59,30,28,31,26,31,11,31,24,31,153,31,45,31,182,31,182,30,182,29,210,31,33,31,67,31,67,30,165,31,70,31,70,30,228,31,60,31,235,31,216,31,225,31,225,30,51,31,46,31,193,31,59,31,167,31,204,31,4,31,179,31,142,31,110,31,243,31,116,31,18,31,18,30,79,31,118,31,105,31,105,30,19,31,171,31,171,30,171,29,94,31,147,31,254,31,247,31,247,30,121,31,146,31,220,31,150,31,250,31,220,31,201,31,201,30,116,31,81,31,105,31,66,31,121,31,1,31,70,31,70,30,218,31,204,31,5,31,196,31,91,31,233,31,255,31,255,30,119,31,255,31,134,31,149,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
