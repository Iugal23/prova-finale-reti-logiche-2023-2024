-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_541 is
end project_tb_541;

architecture project_tb_arch_541 of project_tb_541 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 796;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (172,0,33,0,186,0,186,0,112,0,106,0,0,0,16,0,27,0,78,0,177,0,211,0,125,0,0,0,96,0,205,0,99,0,113,0,241,0,43,0,102,0,29,0,98,0,0,0,93,0,176,0,203,0,174,0,0,0,202,0,215,0,81,0,236,0,148,0,86,0,248,0,137,0,53,0,16,0,74,0,0,0,19,0,0,0,0,0,253,0,175,0,0,0,0,0,191,0,0,0,195,0,70,0,210,0,5,0,70,0,8,0,176,0,45,0,4,0,0,0,243,0,164,0,102,0,188,0,149,0,193,0,76,0,27,0,0,0,92,0,123,0,109,0,1,0,253,0,202,0,132,0,204,0,80,0,214,0,230,0,53,0,221,0,31,0,0,0,100,0,144,0,27,0,20,0,53,0,0,0,150,0,0,0,117,0,195,0,149,0,13,0,0,0,64,0,0,0,58,0,148,0,179,0,22,0,165,0,0,0,141,0,38,0,70,0,254,0,53,0,78,0,169,0,0,0,0,0,4,0,241,0,75,0,187,0,121,0,169,0,0,0,148,0,32,0,0,0,238,0,0,0,210,0,63,0,81,0,0,0,0,0,143,0,76,0,182,0,0,0,113,0,111,0,198,0,61,0,218,0,151,0,154,0,49,0,142,0,10,0,0,0,199,0,50,0,143,0,48,0,85,0,63,0,206,0,46,0,214,0,95,0,0,0,118,0,0,0,125,0,161,0,226,0,224,0,0,0,201,0,189,0,60,0,0,0,15,0,89,0,0,0,102,0,0,0,0,0,224,0,0,0,0,0,73,0,145,0,0,0,59,0,0,0,113,0,30,0,41,0,31,0,122,0,159,0,0,0,230,0,98,0,232,0,186,0,43,0,118,0,57,0,0,0,0,0,151,0,0,0,243,0,77,0,223,0,87,0,16,0,150,0,86,0,0,0,101,0,20,0,0,0,224,0,0,0,192,0,0,0,0,0,38,0,22,0,223,0,254,0,0,0,123,0,134,0,0,0,150,0,67,0,0,0,140,0,0,0,188,0,125,0,151,0,216,0,60,0,0,0,138,0,191,0,147,0,61,0,190,0,4,0,35,0,229,0,112,0,111,0,218,0,0,0,174,0,229,0,206,0,179,0,23,0,129,0,0,0,90,0,155,0,70,0,85,0,248,0,45,0,117,0,92,0,210,0,187,0,212,0,199,0,124,0,202,0,112,0,52,0,231,0,229,0,211,0,4,0,0,0,80,0,115,0,113,0,20,0,145,0,211,0,130,0,126,0,6,0,12,0,0,0,137,0,0,0,25,0,54,0,127,0,0,0,0,0,55,0,121,0,0,0,157,0,21,0,25,0,84,0,191,0,57,0,16,0,27,0,50,0,0,0,185,0,0,0,227,0,21,0,246,0,167,0,96,0,232,0,65,0,194,0,218,0,199,0,0,0,0,0,135,0,214,0,119,0,165,0,0,0,86,0,117,0,19,0,34,0,0,0,164,0,217,0,28,0,148,0,24,0,156,0,148,0,233,0,252,0,253,0,189,0,0,0,43,0,44,0,15,0,0,0,147,0,48,0,172,0,226,0,170,0,0,0,0,0,0,0,51,0,147,0,25,0,209,0,67,0,0,0,147,0,88,0,192,0,0,0,169,0,177,0,154,0,198,0,0,0,170,0,94,0,65,0,131,0,0,0,67,0,237,0,228,0,0,0,253,0,218,0,197,0,135,0,7,0,0,0,196,0,68,0,120,0,0,0,98,0,51,0,236,0,0,0,202,0,102,0,55,0,178,0,0,0,34,0,0,0,207,0,233,0,227,0,32,0,0,0,39,0,46,0,168,0,141,0,130,0,25,0,168,0,0,0,39,0,62,0,84,0,121,0,0,0,38,0,145,0,197,0,12,0,51,0,0,0,221,0,0,0,47,0,0,0,0,0,0,0,100,0,112,0,209,0,136,0,6,0,92,0,215,0,178,0,41,0,3,0,77,0,164,0,73,0,80,0,150,0,242,0,0,0,197,0,21,0,71,0,148,0,237,0,80,0,95,0,180,0,0,0,0,0,117,0,182,0,226,0,184,0,177,0,204,0,177,0,23,0,93,0,217,0,246,0,126,0,38,0,144,0,108,0,140,0,113,0,0,0,214,0,197,0,22,0,72,0,0,0,15,0,76,0,0,0,231,0,0,0,239,0,149,0,71,0,246,0,49,0,112,0,0,0,0,0,91,0,245,0,0,0,28,0,231,0,247,0,81,0,1,0,0,0,25,0,0,0,0,0,117,0,13,0,90,0,3,0,38,0,202,0,139,0,0,0,0,0,209,0,0,0,241,0,57,0,45,0,55,0,63,0,173,0,0,0,115,0,0,0,64,0,233,0,61,0,250,0,0,0,90,0,145,0,195,0,4,0,0,0,154,0,0,0,239,0,105,0,74,0,154,0,112,0,0,0,105,0,88,0,47,0,206,0,128,0,0,0,154,0,199,0,34,0,142,0,0,0,92,0,47,0,170,0,0,0,26,0,79,0,20,0,0,0,182,0,224,0,177,0,235,0,79,0,187,0,2,0,50,0,0,0,0,0,0,0,60,0,59,0,0,0,182,0,119,0,17,0,0,0,219,0,78,0,14,0,198,0,91,0,199,0,0,0,0,0,58,0,128,0,130,0,240,0,13,0,0,0,182,0,109,0,14,0,200,0,0,0,62,0,208,0,93,0,235,0,12,0,242,0,22,0,48,0,212,0,0,0,82,0,40,0,54,0,122,0,0,0,0,0,76,0,16,0,171,0,192,0,0,0,251,0,80,0,140,0,39,0,216,0,0,0,226,0,164,0,64,0,0,0,214,0,162,0,0,0,173,0,72,0,54,0,90,0,28,0,81,0,27,0,0,0,252,0,32,0,191,0,50,0,105,0,0,0,5,0,10,0,28,0,94,0,106,0,67,0,0,0,237,0,184,0,45,0,224,0,12,0,29,0,0,0,0,0,23,0,107,0,185,0,0,0,149,0,46,0,127,0,251,0,167,0,166,0,0,0,0,0,162,0,142,0,237,0,193,0,197,0,187,0,0,0,104,0,139,0,0,0,0,0,212,0,90,0,0,0,151,0,95,0,252,0,128,0,0,0,28,0,206,0,244,0,83,0,108,0,0,0,37,0,66,0,160,0,100,0,76,0,252,0,236,0,95,0,70,0,0,0,3,0,0,0,0,0,0,0,225,0,218,0,0,0,84,0,17,0,0,0,193,0,16,0,0,0,36,0,0,0,83,0,0,0,236,0,64,0,114,0,175,0,0,0,96,0,91,0,0,0,44,0,87,0,92,0,253,0,165,0,203,0,8,0,19,0,96,0,112,0,244,0,177,0,185,0,140,0,148,0,200,0,161,0,218,0,155,0,97,0,88,0,211,0,35,0,0,0,152,0,194,0,106,0,157,0,0,0,194,0,161,0,62,0,135,0,189,0,71,0,251,0,95,0,28,0,59,0,192,0,151,0,246,0,199,0,111,0,65,0,80,0,140,0,249,0,168,0,193,0,213,0,104,0,0,0,224,0,0,0,87,0,0,0,19,0,0,0,175,0,0,0,30,0,217,0);
signal scenario_full  : scenario_type := (172,31,33,31,186,31,186,31,112,31,106,31,106,30,16,31,27,31,78,31,177,31,211,31,125,31,125,30,96,31,205,31,99,31,113,31,241,31,43,31,102,31,29,31,98,31,98,30,93,31,176,31,203,31,174,31,174,30,202,31,215,31,81,31,236,31,148,31,86,31,248,31,137,31,53,31,16,31,74,31,74,30,19,31,19,30,19,29,253,31,175,31,175,30,175,29,191,31,191,30,195,31,70,31,210,31,5,31,70,31,8,31,176,31,45,31,4,31,4,30,243,31,164,31,102,31,188,31,149,31,193,31,76,31,27,31,27,30,92,31,123,31,109,31,1,31,253,31,202,31,132,31,204,31,80,31,214,31,230,31,53,31,221,31,31,31,31,30,100,31,144,31,27,31,20,31,53,31,53,30,150,31,150,30,117,31,195,31,149,31,13,31,13,30,64,31,64,30,58,31,148,31,179,31,22,31,165,31,165,30,141,31,38,31,70,31,254,31,53,31,78,31,169,31,169,30,169,29,4,31,241,31,75,31,187,31,121,31,169,31,169,30,148,31,32,31,32,30,238,31,238,30,210,31,63,31,81,31,81,30,81,29,143,31,76,31,182,31,182,30,113,31,111,31,198,31,61,31,218,31,151,31,154,31,49,31,142,31,10,31,10,30,199,31,50,31,143,31,48,31,85,31,63,31,206,31,46,31,214,31,95,31,95,30,118,31,118,30,125,31,161,31,226,31,224,31,224,30,201,31,189,31,60,31,60,30,15,31,89,31,89,30,102,31,102,30,102,29,224,31,224,30,224,29,73,31,145,31,145,30,59,31,59,30,113,31,30,31,41,31,31,31,122,31,159,31,159,30,230,31,98,31,232,31,186,31,43,31,118,31,57,31,57,30,57,29,151,31,151,30,243,31,77,31,223,31,87,31,16,31,150,31,86,31,86,30,101,31,20,31,20,30,224,31,224,30,192,31,192,30,192,29,38,31,22,31,223,31,254,31,254,30,123,31,134,31,134,30,150,31,67,31,67,30,140,31,140,30,188,31,125,31,151,31,216,31,60,31,60,30,138,31,191,31,147,31,61,31,190,31,4,31,35,31,229,31,112,31,111,31,218,31,218,30,174,31,229,31,206,31,179,31,23,31,129,31,129,30,90,31,155,31,70,31,85,31,248,31,45,31,117,31,92,31,210,31,187,31,212,31,199,31,124,31,202,31,112,31,52,31,231,31,229,31,211,31,4,31,4,30,80,31,115,31,113,31,20,31,145,31,211,31,130,31,126,31,6,31,12,31,12,30,137,31,137,30,25,31,54,31,127,31,127,30,127,29,55,31,121,31,121,30,157,31,21,31,25,31,84,31,191,31,57,31,16,31,27,31,50,31,50,30,185,31,185,30,227,31,21,31,246,31,167,31,96,31,232,31,65,31,194,31,218,31,199,31,199,30,199,29,135,31,214,31,119,31,165,31,165,30,86,31,117,31,19,31,34,31,34,30,164,31,217,31,28,31,148,31,24,31,156,31,148,31,233,31,252,31,253,31,189,31,189,30,43,31,44,31,15,31,15,30,147,31,48,31,172,31,226,31,170,31,170,30,170,29,170,28,51,31,147,31,25,31,209,31,67,31,67,30,147,31,88,31,192,31,192,30,169,31,177,31,154,31,198,31,198,30,170,31,94,31,65,31,131,31,131,30,67,31,237,31,228,31,228,30,253,31,218,31,197,31,135,31,7,31,7,30,196,31,68,31,120,31,120,30,98,31,51,31,236,31,236,30,202,31,102,31,55,31,178,31,178,30,34,31,34,30,207,31,233,31,227,31,32,31,32,30,39,31,46,31,168,31,141,31,130,31,25,31,168,31,168,30,39,31,62,31,84,31,121,31,121,30,38,31,145,31,197,31,12,31,51,31,51,30,221,31,221,30,47,31,47,30,47,29,47,28,100,31,112,31,209,31,136,31,6,31,92,31,215,31,178,31,41,31,3,31,77,31,164,31,73,31,80,31,150,31,242,31,242,30,197,31,21,31,71,31,148,31,237,31,80,31,95,31,180,31,180,30,180,29,117,31,182,31,226,31,184,31,177,31,204,31,177,31,23,31,93,31,217,31,246,31,126,31,38,31,144,31,108,31,140,31,113,31,113,30,214,31,197,31,22,31,72,31,72,30,15,31,76,31,76,30,231,31,231,30,239,31,149,31,71,31,246,31,49,31,112,31,112,30,112,29,91,31,245,31,245,30,28,31,231,31,247,31,81,31,1,31,1,30,25,31,25,30,25,29,117,31,13,31,90,31,3,31,38,31,202,31,139,31,139,30,139,29,209,31,209,30,241,31,57,31,45,31,55,31,63,31,173,31,173,30,115,31,115,30,64,31,233,31,61,31,250,31,250,30,90,31,145,31,195,31,4,31,4,30,154,31,154,30,239,31,105,31,74,31,154,31,112,31,112,30,105,31,88,31,47,31,206,31,128,31,128,30,154,31,199,31,34,31,142,31,142,30,92,31,47,31,170,31,170,30,26,31,79,31,20,31,20,30,182,31,224,31,177,31,235,31,79,31,187,31,2,31,50,31,50,30,50,29,50,28,60,31,59,31,59,30,182,31,119,31,17,31,17,30,219,31,78,31,14,31,198,31,91,31,199,31,199,30,199,29,58,31,128,31,130,31,240,31,13,31,13,30,182,31,109,31,14,31,200,31,200,30,62,31,208,31,93,31,235,31,12,31,242,31,22,31,48,31,212,31,212,30,82,31,40,31,54,31,122,31,122,30,122,29,76,31,16,31,171,31,192,31,192,30,251,31,80,31,140,31,39,31,216,31,216,30,226,31,164,31,64,31,64,30,214,31,162,31,162,30,173,31,72,31,54,31,90,31,28,31,81,31,27,31,27,30,252,31,32,31,191,31,50,31,105,31,105,30,5,31,10,31,28,31,94,31,106,31,67,31,67,30,237,31,184,31,45,31,224,31,12,31,29,31,29,30,29,29,23,31,107,31,185,31,185,30,149,31,46,31,127,31,251,31,167,31,166,31,166,30,166,29,162,31,142,31,237,31,193,31,197,31,187,31,187,30,104,31,139,31,139,30,139,29,212,31,90,31,90,30,151,31,95,31,252,31,128,31,128,30,28,31,206,31,244,31,83,31,108,31,108,30,37,31,66,31,160,31,100,31,76,31,252,31,236,31,95,31,70,31,70,30,3,31,3,30,3,29,3,28,225,31,218,31,218,30,84,31,17,31,17,30,193,31,16,31,16,30,36,31,36,30,83,31,83,30,236,31,64,31,114,31,175,31,175,30,96,31,91,31,91,30,44,31,87,31,92,31,253,31,165,31,203,31,8,31,19,31,96,31,112,31,244,31,177,31,185,31,140,31,148,31,200,31,161,31,218,31,155,31,97,31,88,31,211,31,35,31,35,30,152,31,194,31,106,31,157,31,157,30,194,31,161,31,62,31,135,31,189,31,71,31,251,31,95,31,28,31,59,31,192,31,151,31,246,31,199,31,111,31,65,31,80,31,140,31,249,31,168,31,193,31,213,31,104,31,104,30,224,31,224,30,87,31,87,30,19,31,19,30,175,31,175,30,30,31,217,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
