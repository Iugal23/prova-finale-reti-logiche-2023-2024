-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 251;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (7,0,239,0,0,0,74,0,35,0,56,0,227,0,188,0,0,0,0,0,115,0,243,0,7,0,32,0,96,0,207,0,9,0,164,0,88,0,0,0,0,0,0,0,6,0,191,0,253,0,5,0,15,0,90,0,155,0,146,0,169,0,192,0,237,0,128,0,0,0,155,0,0,0,14,0,0,0,0,0,90,0,142,0,228,0,115,0,230,0,170,0,43,0,0,0,29,0,18,0,162,0,0,0,232,0,177,0,221,0,188,0,244,0,57,0,0,0,50,0,154,0,241,0,0,0,81,0,156,0,0,0,78,0,36,0,187,0,228,0,117,0,204,0,20,0,134,0,111,0,249,0,13,0,81,0,71,0,161,0,38,0,1,0,88,0,0,0,252,0,3,0,0,0,20,0,104,0,51,0,0,0,0,0,83,0,44,0,40,0,226,0,179,0,45,0,189,0,91,0,144,0,199,0,177,0,171,0,155,0,0,0,103,0,0,0,31,0,190,0,0,0,120,0,115,0,99,0,206,0,152,0,0,0,244,0,235,0,20,0,146,0,0,0,0,0,100,0,0,0,242,0,172,0,189,0,157,0,242,0,0,0,124,0,0,0,135,0,0,0,0,0,147,0,104,0,196,0,0,0,0,0,0,0,224,0,155,0,0,0,34,0,89,0,26,0,225,0,34,0,8,0,132,0,0,0,157,0,112,0,65,0,157,0,90,0,0,0,29,0,232,0,167,0,230,0,215,0,22,0,168,0,181,0,199,0,221,0,64,0,240,0,108,0,233,0,171,0,173,0,0,0,0,0,174,0,167,0,144,0,0,0,105,0,61,0,77,0,13,0,134,0,245,0,253,0,0,0,159,0,172,0,153,0,126,0,43,0,4,0,210,0,39,0,20,0,94,0,36,0,151,0,192,0,198,0,207,0,96,0,234,0,53,0,3,0,173,0,255,0,185,0,142,0,231,0,133,0,150,0,0,0,106,0,0,0,197,0,248,0,212,0,56,0,223,0,108,0,78,0,107,0,0,0,249,0,97,0,0,0,0,0,132,0,0,0,205,0,166,0,166,0,0,0,42,0,58,0,0,0,1,0,0,0,27,0,0,0,36,0,80,0,116,0,12,0,0,0,114,0,0,0);
signal scenario_full  : scenario_type := (7,31,239,31,239,30,74,31,35,31,56,31,227,31,188,31,188,30,188,29,115,31,243,31,7,31,32,31,96,31,207,31,9,31,164,31,88,31,88,30,88,29,88,28,6,31,191,31,253,31,5,31,15,31,90,31,155,31,146,31,169,31,192,31,237,31,128,31,128,30,155,31,155,30,14,31,14,30,14,29,90,31,142,31,228,31,115,31,230,31,170,31,43,31,43,30,29,31,18,31,162,31,162,30,232,31,177,31,221,31,188,31,244,31,57,31,57,30,50,31,154,31,241,31,241,30,81,31,156,31,156,30,78,31,36,31,187,31,228,31,117,31,204,31,20,31,134,31,111,31,249,31,13,31,81,31,71,31,161,31,38,31,1,31,88,31,88,30,252,31,3,31,3,30,20,31,104,31,51,31,51,30,51,29,83,31,44,31,40,31,226,31,179,31,45,31,189,31,91,31,144,31,199,31,177,31,171,31,155,31,155,30,103,31,103,30,31,31,190,31,190,30,120,31,115,31,99,31,206,31,152,31,152,30,244,31,235,31,20,31,146,31,146,30,146,29,100,31,100,30,242,31,172,31,189,31,157,31,242,31,242,30,124,31,124,30,135,31,135,30,135,29,147,31,104,31,196,31,196,30,196,29,196,28,224,31,155,31,155,30,34,31,89,31,26,31,225,31,34,31,8,31,132,31,132,30,157,31,112,31,65,31,157,31,90,31,90,30,29,31,232,31,167,31,230,31,215,31,22,31,168,31,181,31,199,31,221,31,64,31,240,31,108,31,233,31,171,31,173,31,173,30,173,29,174,31,167,31,144,31,144,30,105,31,61,31,77,31,13,31,134,31,245,31,253,31,253,30,159,31,172,31,153,31,126,31,43,31,4,31,210,31,39,31,20,31,94,31,36,31,151,31,192,31,198,31,207,31,96,31,234,31,53,31,3,31,173,31,255,31,185,31,142,31,231,31,133,31,150,31,150,30,106,31,106,30,197,31,248,31,212,31,56,31,223,31,108,31,78,31,107,31,107,30,249,31,97,31,97,30,97,29,132,31,132,30,205,31,166,31,166,31,166,30,42,31,58,31,58,30,1,31,1,30,27,31,27,30,36,31,80,31,116,31,12,31,12,30,114,31,114,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
