-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_963 is
end project_tb_963;

architecture project_tb_arch_963 of project_tb_963 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 422;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (179,0,222,0,0,0,26,0,39,0,0,0,109,0,0,0,227,0,63,0,0,0,0,0,0,0,18,0,0,0,230,0,0,0,212,0,249,0,87,0,0,0,27,0,170,0,0,0,0,0,141,0,44,0,0,0,75,0,249,0,117,0,188,0,179,0,201,0,215,0,38,0,0,0,0,0,0,0,173,0,134,0,73,0,73,0,229,0,156,0,225,0,6,0,0,0,0,0,116,0,52,0,0,0,0,0,206,0,175,0,94,0,111,0,115,0,238,0,161,0,48,0,52,0,241,0,137,0,204,0,249,0,224,0,0,0,21,0,0,0,0,0,233,0,0,0,0,0,149,0,199,0,146,0,0,0,157,0,0,0,244,0,149,0,64,0,136,0,0,0,215,0,97,0,0,0,226,0,0,0,78,0,117,0,0,0,106,0,0,0,0,0,185,0,0,0,152,0,30,0,13,0,183,0,116,0,58,0,12,0,14,0,228,0,143,0,111,0,88,0,236,0,115,0,0,0,0,0,199,0,66,0,46,0,21,0,172,0,133,0,189,0,80,0,196,0,1,0,46,0,0,0,217,0,39,0,170,0,138,0,105,0,64,0,13,0,194,0,150,0,33,0,93,0,8,0,148,0,59,0,79,0,0,0,145,0,159,0,76,0,48,0,190,0,46,0,196,0,173,0,123,0,180,0,140,0,15,0,63,0,73,0,134,0,0,0,245,0,124,0,154,0,167,0,0,0,165,0,0,0,0,0,217,0,152,0,252,0,134,0,80,0,41,0,103,0,99,0,0,0,5,0,98,0,165,0,44,0,0,0,3,0,130,0,113,0,126,0,21,0,192,0,132,0,15,0,113,0,0,0,190,0,11,0,40,0,187,0,255,0,146,0,225,0,147,0,154,0,101,0,10,0,198,0,165,0,2,0,91,0,202,0,180,0,71,0,8,0,121,0,186,0,129,0,166,0,96,0,122,0,132,0,136,0,0,0,167,0,136,0,176,0,0,0,0,0,5,0,0,0,176,0,105,0,195,0,165,0,229,0,0,0,0,0,76,0,170,0,0,0,209,0,0,0,89,0,238,0,51,0,93,0,171,0,249,0,238,0,90,0,73,0,238,0,207,0,90,0,41,0,44,0,102,0,149,0,13,0,87,0,73,0,0,0,58,0,30,0,235,0,9,0,0,0,0,0,113,0,0,0,114,0,161,0,0,0,8,0,213,0,0,0,213,0,53,0,106,0,155,0,11,0,154,0,201,0,101,0,202,0,197,0,198,0,55,0,170,0,34,0,124,0,128,0,13,0,88,0,85,0,0,0,140,0,101,0,64,0,12,0,55,0,250,0,166,0,0,0,48,0,0,0,221,0,37,0,68,0,160,0,185,0,174,0,0,0,237,0,78,0,115,0,9,0,177,0,67,0,0,0,61,0,0,0,106,0,154,0,63,0,0,0,40,0,84,0,11,0,201,0,36,0,150,0,211,0,182,0,47,0,55,0,152,0,216,0,0,0,152,0,61,0,145,0,0,0,175,0,0,0,232,0,194,0,221,0,0,0,245,0,214,0,160,0,50,0,0,0,0,0,0,0,172,0,48,0,185,0,232,0,198,0,221,0,175,0,132,0,202,0,57,0,184,0,0,0,0,0,13,0,0,0,142,0,11,0,0,0,50,0,138,0,215,0,242,0,0,0,181,0,0,0,147,0,245,0,45,0,215,0,20,0,216,0,228,0,0,0,99,0,5,0,130,0,45,0,172,0,156,0,140,0,186,0,96,0,0,0,231,0,21,0,115,0,77,0,100,0,0,0,227,0,0,0,99,0,115,0,19,0,123,0,0,0,162,0,68,0,0,0,0,0,192,0,179,0,0,0,22,0,209,0,19,0,0,0,194,0,147,0,11,0,172,0);
signal scenario_full  : scenario_type := (179,31,222,31,222,30,26,31,39,31,39,30,109,31,109,30,227,31,63,31,63,30,63,29,63,28,18,31,18,30,230,31,230,30,212,31,249,31,87,31,87,30,27,31,170,31,170,30,170,29,141,31,44,31,44,30,75,31,249,31,117,31,188,31,179,31,201,31,215,31,38,31,38,30,38,29,38,28,173,31,134,31,73,31,73,31,229,31,156,31,225,31,6,31,6,30,6,29,116,31,52,31,52,30,52,29,206,31,175,31,94,31,111,31,115,31,238,31,161,31,48,31,52,31,241,31,137,31,204,31,249,31,224,31,224,30,21,31,21,30,21,29,233,31,233,30,233,29,149,31,199,31,146,31,146,30,157,31,157,30,244,31,149,31,64,31,136,31,136,30,215,31,97,31,97,30,226,31,226,30,78,31,117,31,117,30,106,31,106,30,106,29,185,31,185,30,152,31,30,31,13,31,183,31,116,31,58,31,12,31,14,31,228,31,143,31,111,31,88,31,236,31,115,31,115,30,115,29,199,31,66,31,46,31,21,31,172,31,133,31,189,31,80,31,196,31,1,31,46,31,46,30,217,31,39,31,170,31,138,31,105,31,64,31,13,31,194,31,150,31,33,31,93,31,8,31,148,31,59,31,79,31,79,30,145,31,159,31,76,31,48,31,190,31,46,31,196,31,173,31,123,31,180,31,140,31,15,31,63,31,73,31,134,31,134,30,245,31,124,31,154,31,167,31,167,30,165,31,165,30,165,29,217,31,152,31,252,31,134,31,80,31,41,31,103,31,99,31,99,30,5,31,98,31,165,31,44,31,44,30,3,31,130,31,113,31,126,31,21,31,192,31,132,31,15,31,113,31,113,30,190,31,11,31,40,31,187,31,255,31,146,31,225,31,147,31,154,31,101,31,10,31,198,31,165,31,2,31,91,31,202,31,180,31,71,31,8,31,121,31,186,31,129,31,166,31,96,31,122,31,132,31,136,31,136,30,167,31,136,31,176,31,176,30,176,29,5,31,5,30,176,31,105,31,195,31,165,31,229,31,229,30,229,29,76,31,170,31,170,30,209,31,209,30,89,31,238,31,51,31,93,31,171,31,249,31,238,31,90,31,73,31,238,31,207,31,90,31,41,31,44,31,102,31,149,31,13,31,87,31,73,31,73,30,58,31,30,31,235,31,9,31,9,30,9,29,113,31,113,30,114,31,161,31,161,30,8,31,213,31,213,30,213,31,53,31,106,31,155,31,11,31,154,31,201,31,101,31,202,31,197,31,198,31,55,31,170,31,34,31,124,31,128,31,13,31,88,31,85,31,85,30,140,31,101,31,64,31,12,31,55,31,250,31,166,31,166,30,48,31,48,30,221,31,37,31,68,31,160,31,185,31,174,31,174,30,237,31,78,31,115,31,9,31,177,31,67,31,67,30,61,31,61,30,106,31,154,31,63,31,63,30,40,31,84,31,11,31,201,31,36,31,150,31,211,31,182,31,47,31,55,31,152,31,216,31,216,30,152,31,61,31,145,31,145,30,175,31,175,30,232,31,194,31,221,31,221,30,245,31,214,31,160,31,50,31,50,30,50,29,50,28,172,31,48,31,185,31,232,31,198,31,221,31,175,31,132,31,202,31,57,31,184,31,184,30,184,29,13,31,13,30,142,31,11,31,11,30,50,31,138,31,215,31,242,31,242,30,181,31,181,30,147,31,245,31,45,31,215,31,20,31,216,31,228,31,228,30,99,31,5,31,130,31,45,31,172,31,156,31,140,31,186,31,96,31,96,30,231,31,21,31,115,31,77,31,100,31,100,30,227,31,227,30,99,31,115,31,19,31,123,31,123,30,162,31,68,31,68,30,68,29,192,31,179,31,179,30,22,31,209,31,19,31,19,30,194,31,147,31,11,31,172,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
