-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_972 is
end project_tb_972;

architecture project_tb_arch_972 of project_tb_972 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 746;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (48,0,0,0,90,0,0,0,125,0,172,0,216,0,170,0,67,0,161,0,41,0,224,0,3,0,0,0,3,0,210,0,0,0,129,0,0,0,193,0,226,0,0,0,0,0,0,0,0,0,196,0,213,0,0,0,21,0,0,0,252,0,60,0,39,0,163,0,123,0,0,0,195,0,110,0,131,0,184,0,28,0,108,0,61,0,194,0,209,0,251,0,116,0,179,0,224,0,37,0,244,0,236,0,188,0,191,0,45,0,181,0,117,0,3,0,65,0,152,0,33,0,0,0,143,0,101,0,0,0,75,0,154,0,0,0,0,0,0,0,125,0,0,0,142,0,196,0,52,0,0,0,122,0,190,0,128,0,124,0,137,0,0,0,165,0,173,0,123,0,176,0,0,0,114,0,0,0,125,0,142,0,91,0,165,0,241,0,0,0,21,0,160,0,251,0,177,0,48,0,148,0,240,0,18,0,38,0,0,0,77,0,252,0,138,0,212,0,67,0,253,0,118,0,0,0,125,0,227,0,55,0,60,0,163,0,92,0,0,0,19,0,0,0,190,0,2,0,226,0,84,0,112,0,116,0,0,0,25,0,0,0,195,0,21,0,0,0,49,0,229,0,24,0,19,0,109,0,15,0,12,0,209,0,0,0,222,0,21,0,71,0,0,0,200,0,33,0,0,0,0,0,0,0,140,0,0,0,0,0,168,0,0,0,65,0,95,0,224,0,0,0,0,0,204,0,115,0,210,0,13,0,27,0,0,0,1,0,219,0,245,0,0,0,164,0,147,0,170,0,76,0,225,0,21,0,118,0,209,0,190,0,53,0,54,0,202,0,0,0,60,0,110,0,85,0,6,0,113,0,27,0,93,0,6,0,179,0,52,0,68,0,86,0,222,0,194,0,52,0,254,0,169,0,1,0,177,0,56,0,198,0,136,0,0,0,104,0,167,0,53,0,186,0,23,0,83,0,179,0,69,0,91,0,16,0,0,0,112,0,83,0,40,0,157,0,90,0,0,0,7,0,110,0,103,0,93,0,165,0,224,0,15,0,241,0,0,0,182,0,166,0,67,0,224,0,0,0,177,0,126,0,0,0,37,0,0,0,207,0,158,0,108,0,39,0,173,0,209,0,218,0,217,0,90,0,184,0,54,0,235,0,20,0,94,0,106,0,101,0,128,0,76,0,17,0,88,0,0,0,14,0,177,0,19,0,176,0,21,0,235,0,247,0,123,0,0,0,171,0,1,0,238,0,49,0,62,0,101,0,138,0,229,0,0,0,176,0,200,0,0,0,0,0,176,0,124,0,0,0,4,0,246,0,46,0,121,0,183,0,14,0,243,0,119,0,113,0,87,0,0,0,0,0,92,0,82,0,183,0,0,0,0,0,123,0,239,0,183,0,235,0,130,0,163,0,123,0,53,0,0,0,105,0,120,0,119,0,188,0,88,0,157,0,197,0,227,0,232,0,0,0,0,0,165,0,0,0,63,0,245,0,124,0,25,0,45,0,169,0,0,0,55,0,240,0,214,0,68,0,116,0,0,0,237,0,184,0,186,0,0,0,61,0,226,0,0,0,37,0,37,0,164,0,0,0,190,0,207,0,228,0,198,0,0,0,183,0,81,0,0,0,0,0,148,0,157,0,112,0,173,0,16,0,108,0,0,0,0,0,63,0,62,0,169,0,36,0,54,0,0,0,162,0,239,0,54,0,86,0,98,0,31,0,71,0,20,0,164,0,0,0,65,0,0,0,124,0,0,0,185,0,166,0,0,0,7,0,0,0,0,0,53,0,0,0,59,0,75,0,0,0,0,0,11,0,0,0,144,0,119,0,172,0,223,0,0,0,251,0,177,0,243,0,164,0,101,0,69,0,205,0,159,0,251,0,48,0,131,0,30,0,6,0,166,0,189,0,78,0,158,0,0,0,0,0,176,0,0,0,228,0,114,0,0,0,253,0,0,0,114,0,148,0,0,0,134,0,171,0,14,0,90,0,0,0,170,0,0,0,0,0,103,0,206,0,139,0,0,0,0,0,211,0,140,0,64,0,235,0,176,0,112,0,39,0,88,0,219,0,235,0,72,0,7,0,0,0,121,0,171,0,0,0,188,0,49,0,0,0,100,0,80,0,212,0,218,0,243,0,113,0,76,0,73,0,87,0,231,0,170,0,27,0,140,0,13,0,62,0,69,0,102,0,110,0,243,0,55,0,0,0,145,0,59,0,65,0,193,0,116,0,73,0,223,0,54,0,244,0,232,0,216,0,140,0,62,0,0,0,134,0,180,0,54,0,146,0,150,0,101,0,123,0,0,0,58,0,63,0,0,0,0,0,204,0,207,0,179,0,129,0,212,0,158,0,168,0,0,0,30,0,0,0,134,0,0,0,224,0,103,0,240,0,105,0,0,0,54,0,131,0,79,0,187,0,67,0,8,0,168,0,96,0,5,0,134,0,98,0,0,0,0,0,31,0,222,0,191,0,14,0,18,0,196,0,247,0,0,0,51,0,191,0,38,0,137,0,147,0,226,0,0,0,0,0,96,0,250,0,180,0,232,0,24,0,169,0,19,0,225,0,95,0,0,0,221,0,205,0,16,0,158,0,138,0,119,0,191,0,246,0,183,0,209,0,151,0,0,0,0,0,0,0,0,0,224,0,245,0,30,0,15,0,128,0,242,0,214,0,255,0,129,0,223,0,1,0,181,0,60,0,227,0,0,0,43,0,4,0,208,0,83,0,230,0,165,0,245,0,105,0,171,0,56,0,0,0,220,0,124,0,121,0,0,0,253,0,128,0,162,0,0,0,0,0,0,0,161,0,0,0,17,0,195,0,110,0,27,0,0,0,71,0,56,0,127,0,98,0,156,0,107,0,0,0,0,0,0,0,8,0,162,0,92,0,19,0,164,0,190,0,39,0,176,0,250,0,56,0,0,0,43,0,88,0,135,0,85,0,70,0,37,0,153,0,63,0,95,0,193,0,122,0,118,0,0,0,131,0,159,0,152,0,131,0,120,0,173,0,161,0,39,0,246,0,90,0,233,0,182,0,149,0,77,0,0,0,0,0,123,0,6,0,0,0,64,0,129,0,169,0,8,0,9,0,159,0,187,0,5,0,0,0,25,0,28,0,103,0,36,0,28,0,171,0,45,0,0,0,223,0,79,0,39,0,0,0,21,0,219,0,0,0,93,0,30,0,252,0,128,0,202,0,0,0,207,0,46,0,119,0,9,0,185,0,144,0,43,0,74,0,18,0,213,0,124,0,253,0,84,0,0,0,201,0,55,0,86,0,56,0,45,0,246,0,39,0,39,0,72,0,0,0,119,0,0,0,209,0,222,0,200,0,113,0,172,0,0,0,147,0);
signal scenario_full  : scenario_type := (48,31,48,30,90,31,90,30,125,31,172,31,216,31,170,31,67,31,161,31,41,31,224,31,3,31,3,30,3,31,210,31,210,30,129,31,129,30,193,31,226,31,226,30,226,29,226,28,226,27,196,31,213,31,213,30,21,31,21,30,252,31,60,31,39,31,163,31,123,31,123,30,195,31,110,31,131,31,184,31,28,31,108,31,61,31,194,31,209,31,251,31,116,31,179,31,224,31,37,31,244,31,236,31,188,31,191,31,45,31,181,31,117,31,3,31,65,31,152,31,33,31,33,30,143,31,101,31,101,30,75,31,154,31,154,30,154,29,154,28,125,31,125,30,142,31,196,31,52,31,52,30,122,31,190,31,128,31,124,31,137,31,137,30,165,31,173,31,123,31,176,31,176,30,114,31,114,30,125,31,142,31,91,31,165,31,241,31,241,30,21,31,160,31,251,31,177,31,48,31,148,31,240,31,18,31,38,31,38,30,77,31,252,31,138,31,212,31,67,31,253,31,118,31,118,30,125,31,227,31,55,31,60,31,163,31,92,31,92,30,19,31,19,30,190,31,2,31,226,31,84,31,112,31,116,31,116,30,25,31,25,30,195,31,21,31,21,30,49,31,229,31,24,31,19,31,109,31,15,31,12,31,209,31,209,30,222,31,21,31,71,31,71,30,200,31,33,31,33,30,33,29,33,28,140,31,140,30,140,29,168,31,168,30,65,31,95,31,224,31,224,30,224,29,204,31,115,31,210,31,13,31,27,31,27,30,1,31,219,31,245,31,245,30,164,31,147,31,170,31,76,31,225,31,21,31,118,31,209,31,190,31,53,31,54,31,202,31,202,30,60,31,110,31,85,31,6,31,113,31,27,31,93,31,6,31,179,31,52,31,68,31,86,31,222,31,194,31,52,31,254,31,169,31,1,31,177,31,56,31,198,31,136,31,136,30,104,31,167,31,53,31,186,31,23,31,83,31,179,31,69,31,91,31,16,31,16,30,112,31,83,31,40,31,157,31,90,31,90,30,7,31,110,31,103,31,93,31,165,31,224,31,15,31,241,31,241,30,182,31,166,31,67,31,224,31,224,30,177,31,126,31,126,30,37,31,37,30,207,31,158,31,108,31,39,31,173,31,209,31,218,31,217,31,90,31,184,31,54,31,235,31,20,31,94,31,106,31,101,31,128,31,76,31,17,31,88,31,88,30,14,31,177,31,19,31,176,31,21,31,235,31,247,31,123,31,123,30,171,31,1,31,238,31,49,31,62,31,101,31,138,31,229,31,229,30,176,31,200,31,200,30,200,29,176,31,124,31,124,30,4,31,246,31,46,31,121,31,183,31,14,31,243,31,119,31,113,31,87,31,87,30,87,29,92,31,82,31,183,31,183,30,183,29,123,31,239,31,183,31,235,31,130,31,163,31,123,31,53,31,53,30,105,31,120,31,119,31,188,31,88,31,157,31,197,31,227,31,232,31,232,30,232,29,165,31,165,30,63,31,245,31,124,31,25,31,45,31,169,31,169,30,55,31,240,31,214,31,68,31,116,31,116,30,237,31,184,31,186,31,186,30,61,31,226,31,226,30,37,31,37,31,164,31,164,30,190,31,207,31,228,31,198,31,198,30,183,31,81,31,81,30,81,29,148,31,157,31,112,31,173,31,16,31,108,31,108,30,108,29,63,31,62,31,169,31,36,31,54,31,54,30,162,31,239,31,54,31,86,31,98,31,31,31,71,31,20,31,164,31,164,30,65,31,65,30,124,31,124,30,185,31,166,31,166,30,7,31,7,30,7,29,53,31,53,30,59,31,75,31,75,30,75,29,11,31,11,30,144,31,119,31,172,31,223,31,223,30,251,31,177,31,243,31,164,31,101,31,69,31,205,31,159,31,251,31,48,31,131,31,30,31,6,31,166,31,189,31,78,31,158,31,158,30,158,29,176,31,176,30,228,31,114,31,114,30,253,31,253,30,114,31,148,31,148,30,134,31,171,31,14,31,90,31,90,30,170,31,170,30,170,29,103,31,206,31,139,31,139,30,139,29,211,31,140,31,64,31,235,31,176,31,112,31,39,31,88,31,219,31,235,31,72,31,7,31,7,30,121,31,171,31,171,30,188,31,49,31,49,30,100,31,80,31,212,31,218,31,243,31,113,31,76,31,73,31,87,31,231,31,170,31,27,31,140,31,13,31,62,31,69,31,102,31,110,31,243,31,55,31,55,30,145,31,59,31,65,31,193,31,116,31,73,31,223,31,54,31,244,31,232,31,216,31,140,31,62,31,62,30,134,31,180,31,54,31,146,31,150,31,101,31,123,31,123,30,58,31,63,31,63,30,63,29,204,31,207,31,179,31,129,31,212,31,158,31,168,31,168,30,30,31,30,30,134,31,134,30,224,31,103,31,240,31,105,31,105,30,54,31,131,31,79,31,187,31,67,31,8,31,168,31,96,31,5,31,134,31,98,31,98,30,98,29,31,31,222,31,191,31,14,31,18,31,196,31,247,31,247,30,51,31,191,31,38,31,137,31,147,31,226,31,226,30,226,29,96,31,250,31,180,31,232,31,24,31,169,31,19,31,225,31,95,31,95,30,221,31,205,31,16,31,158,31,138,31,119,31,191,31,246,31,183,31,209,31,151,31,151,30,151,29,151,28,151,27,224,31,245,31,30,31,15,31,128,31,242,31,214,31,255,31,129,31,223,31,1,31,181,31,60,31,227,31,227,30,43,31,4,31,208,31,83,31,230,31,165,31,245,31,105,31,171,31,56,31,56,30,220,31,124,31,121,31,121,30,253,31,128,31,162,31,162,30,162,29,162,28,161,31,161,30,17,31,195,31,110,31,27,31,27,30,71,31,56,31,127,31,98,31,156,31,107,31,107,30,107,29,107,28,8,31,162,31,92,31,19,31,164,31,190,31,39,31,176,31,250,31,56,31,56,30,43,31,88,31,135,31,85,31,70,31,37,31,153,31,63,31,95,31,193,31,122,31,118,31,118,30,131,31,159,31,152,31,131,31,120,31,173,31,161,31,39,31,246,31,90,31,233,31,182,31,149,31,77,31,77,30,77,29,123,31,6,31,6,30,64,31,129,31,169,31,8,31,9,31,159,31,187,31,5,31,5,30,25,31,28,31,103,31,36,31,28,31,171,31,45,31,45,30,223,31,79,31,39,31,39,30,21,31,219,31,219,30,93,31,30,31,252,31,128,31,202,31,202,30,207,31,46,31,119,31,9,31,185,31,144,31,43,31,74,31,18,31,213,31,124,31,253,31,84,31,84,30,201,31,55,31,86,31,56,31,45,31,246,31,39,31,39,31,72,31,72,30,119,31,119,30,209,31,222,31,200,31,113,31,172,31,172,30,147,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
