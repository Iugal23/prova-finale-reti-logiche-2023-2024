-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 249;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (83,0,0,0,0,0,39,0,166,0,210,0,242,0,213,0,3,0,58,0,151,0,37,0,179,0,25,0,48,0,94,0,67,0,48,0,10,0,151,0,141,0,0,0,173,0,155,0,102,0,185,0,68,0,131,0,148,0,15,0,233,0,53,0,242,0,131,0,60,0,0,0,252,0,0,0,127,0,42,0,53,0,0,0,48,0,8,0,38,0,0,0,156,0,0,0,203,0,232,0,236,0,146,0,0,0,194,0,170,0,40,0,68,0,224,0,0,0,132,0,212,0,42,0,0,0,110,0,17,0,134,0,128,0,186,0,130,0,0,0,0,0,24,0,241,0,49,0,179,0,8,0,204,0,148,0,183,0,0,0,40,0,0,0,116,0,153,0,20,0,86,0,86,0,147,0,21,0,119,0,0,0,139,0,220,0,0,0,0,0,103,0,0,0,39,0,148,0,118,0,197,0,56,0,206,0,75,0,184,0,115,0,0,0,22,0,156,0,5,0,232,0,226,0,47,0,213,0,229,0,0,0,233,0,87,0,0,0,0,0,164,0,159,0,8,0,180,0,100,0,98,0,148,0,0,0,16,0,0,0,0,0,0,0,209,0,125,0,132,0,88,0,209,0,61,0,58,0,7,0,0,0,80,0,57,0,11,0,58,0,75,0,184,0,47,0,244,0,67,0,160,0,0,0,66,0,213,0,244,0,145,0,119,0,236,0,198,0,0,0,106,0,100,0,0,0,200,0,3,0,12,0,92,0,121,0,121,0,154,0,185,0,83,0,0,0,0,0,116,0,197,0,0,0,0,0,191,0,121,0,154,0,4,0,200,0,40,0,194,0,160,0,72,0,228,0,56,0,95,0,97,0,184,0,237,0,108,0,96,0,22,0,223,0,195,0,168,0,0,0,100,0,0,0,51,0,247,0,0,0,183,0,162,0,45,0,176,0,98,0,193,0,0,0,182,0,34,0,123,0,8,0,61,0,245,0,221,0,0,0,98,0,0,0,56,0,3,0,26,0,36,0,0,0,0,0,16,0,240,0,95,0,199,0,133,0,85,0,69,0,233,0,245,0,53,0,85,0,213,0,213,0,90,0,145,0,146,0,131,0,225,0,234,0,0,0,192,0);
signal scenario_full  : scenario_type := (83,31,83,30,83,29,39,31,166,31,210,31,242,31,213,31,3,31,58,31,151,31,37,31,179,31,25,31,48,31,94,31,67,31,48,31,10,31,151,31,141,31,141,30,173,31,155,31,102,31,185,31,68,31,131,31,148,31,15,31,233,31,53,31,242,31,131,31,60,31,60,30,252,31,252,30,127,31,42,31,53,31,53,30,48,31,8,31,38,31,38,30,156,31,156,30,203,31,232,31,236,31,146,31,146,30,194,31,170,31,40,31,68,31,224,31,224,30,132,31,212,31,42,31,42,30,110,31,17,31,134,31,128,31,186,31,130,31,130,30,130,29,24,31,241,31,49,31,179,31,8,31,204,31,148,31,183,31,183,30,40,31,40,30,116,31,153,31,20,31,86,31,86,31,147,31,21,31,119,31,119,30,139,31,220,31,220,30,220,29,103,31,103,30,39,31,148,31,118,31,197,31,56,31,206,31,75,31,184,31,115,31,115,30,22,31,156,31,5,31,232,31,226,31,47,31,213,31,229,31,229,30,233,31,87,31,87,30,87,29,164,31,159,31,8,31,180,31,100,31,98,31,148,31,148,30,16,31,16,30,16,29,16,28,209,31,125,31,132,31,88,31,209,31,61,31,58,31,7,31,7,30,80,31,57,31,11,31,58,31,75,31,184,31,47,31,244,31,67,31,160,31,160,30,66,31,213,31,244,31,145,31,119,31,236,31,198,31,198,30,106,31,100,31,100,30,200,31,3,31,12,31,92,31,121,31,121,31,154,31,185,31,83,31,83,30,83,29,116,31,197,31,197,30,197,29,191,31,121,31,154,31,4,31,200,31,40,31,194,31,160,31,72,31,228,31,56,31,95,31,97,31,184,31,237,31,108,31,96,31,22,31,223,31,195,31,168,31,168,30,100,31,100,30,51,31,247,31,247,30,183,31,162,31,45,31,176,31,98,31,193,31,193,30,182,31,34,31,123,31,8,31,61,31,245,31,221,31,221,30,98,31,98,30,56,31,3,31,26,31,36,31,36,30,36,29,16,31,240,31,95,31,199,31,133,31,85,31,69,31,233,31,245,31,53,31,85,31,213,31,213,31,90,31,145,31,146,31,131,31,225,31,234,31,234,30,192,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
