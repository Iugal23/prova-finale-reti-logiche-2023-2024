-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 341;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (34,0,192,0,3,0,156,0,0,0,101,0,24,0,0,0,213,0,128,0,211,0,228,0,49,0,0,0,177,0,7,0,0,0,226,0,180,0,187,0,1,0,186,0,161,0,247,0,216,0,252,0,85,0,227,0,8,0,116,0,218,0,6,0,0,0,66,0,246,0,108,0,39,0,26,0,0,0,172,0,180,0,231,0,156,0,234,0,97,0,148,0,58,0,22,0,83,0,204,0,191,0,0,0,0,0,27,0,0,0,31,0,110,0,29,0,0,0,140,0,34,0,172,0,94,0,220,0,94,0,144,0,56,0,0,0,193,0,93,0,23,0,162,0,149,0,122,0,179,0,0,0,123,0,0,0,79,0,137,0,246,0,10,0,18,0,125,0,212,0,82,0,80,0,234,0,129,0,0,0,0,0,28,0,86,0,44,0,83,0,110,0,7,0,176,0,117,0,106,0,239,0,246,0,93,0,231,0,56,0,208,0,0,0,0,0,66,0,95,0,107,0,204,0,0,0,40,0,25,0,250,0,0,0,189,0,133,0,156,0,0,0,84,0,21,0,105,0,184,0,70,0,120,0,97,0,251,0,26,0,0,0,150,0,40,0,90,0,126,0,0,0,0,0,69,0,55,0,215,0,46,0,144,0,0,0,47,0,147,0,7,0,210,0,149,0,53,0,3,0,0,0,0,0,99,0,6,0,146,0,28,0,0,0,0,0,50,0,12,0,0,0,71,0,50,0,205,0,41,0,94,0,202,0,121,0,0,0,0,0,95,0,217,0,186,0,167,0,160,0,24,0,245,0,74,0,9,0,248,0,173,0,234,0,96,0,102,0,33,0,82,0,0,0,0,0,102,0,11,0,175,0,226,0,144,0,177,0,248,0,173,0,0,0,0,0,231,0,165,0,86,0,219,0,145,0,0,0,49,0,25,0,15,0,27,0,159,0,253,0,103,0,191,0,0,0,124,0,42,0,216,0,66,0,203,0,166,0,221,0,0,0,24,0,217,0,229,0,0,0,0,0,127,0,26,0,6,0,183,0,10,0,194,0,62,0,134,0,75,0,106,0,54,0,66,0,144,0,0,0,18,0,193,0,134,0,0,0,63,0,0,0,0,0,234,0,229,0,251,0,57,0,71,0,22,0,0,0,0,0,30,0,0,0,113,0,192,0,15,0,153,0,182,0,115,0,174,0,198,0,223,0,0,0,69,0,215,0,154,0,58,0,42,0,4,0,0,0,206,0,0,0,0,0,0,0,106,0,111,0,0,0,155,0,233,0,205,0,111,0,0,0,74,0,103,0,0,0,0,0,187,0,171,0,108,0,0,0,4,0,250,0,190,0,140,0,239,0,222,0,248,0,0,0,214,0,45,0,0,0,0,0,129,0,0,0,0,0,86,0,137,0,72,0,120,0,195,0,49,0,182,0,230,0,147,0,119,0,147,0,95,0,147,0,109,0,201,0,131,0,168,0,0,0,43,0,53,0,101,0,35,0,0,0,87,0,27,0,0,0,0,0,177,0,0,0,0,0,95,0,174,0);
signal scenario_full  : scenario_type := (34,31,192,31,3,31,156,31,156,30,101,31,24,31,24,30,213,31,128,31,211,31,228,31,49,31,49,30,177,31,7,31,7,30,226,31,180,31,187,31,1,31,186,31,161,31,247,31,216,31,252,31,85,31,227,31,8,31,116,31,218,31,6,31,6,30,66,31,246,31,108,31,39,31,26,31,26,30,172,31,180,31,231,31,156,31,234,31,97,31,148,31,58,31,22,31,83,31,204,31,191,31,191,30,191,29,27,31,27,30,31,31,110,31,29,31,29,30,140,31,34,31,172,31,94,31,220,31,94,31,144,31,56,31,56,30,193,31,93,31,23,31,162,31,149,31,122,31,179,31,179,30,123,31,123,30,79,31,137,31,246,31,10,31,18,31,125,31,212,31,82,31,80,31,234,31,129,31,129,30,129,29,28,31,86,31,44,31,83,31,110,31,7,31,176,31,117,31,106,31,239,31,246,31,93,31,231,31,56,31,208,31,208,30,208,29,66,31,95,31,107,31,204,31,204,30,40,31,25,31,250,31,250,30,189,31,133,31,156,31,156,30,84,31,21,31,105,31,184,31,70,31,120,31,97,31,251,31,26,31,26,30,150,31,40,31,90,31,126,31,126,30,126,29,69,31,55,31,215,31,46,31,144,31,144,30,47,31,147,31,7,31,210,31,149,31,53,31,3,31,3,30,3,29,99,31,6,31,146,31,28,31,28,30,28,29,50,31,12,31,12,30,71,31,50,31,205,31,41,31,94,31,202,31,121,31,121,30,121,29,95,31,217,31,186,31,167,31,160,31,24,31,245,31,74,31,9,31,248,31,173,31,234,31,96,31,102,31,33,31,82,31,82,30,82,29,102,31,11,31,175,31,226,31,144,31,177,31,248,31,173,31,173,30,173,29,231,31,165,31,86,31,219,31,145,31,145,30,49,31,25,31,15,31,27,31,159,31,253,31,103,31,191,31,191,30,124,31,42,31,216,31,66,31,203,31,166,31,221,31,221,30,24,31,217,31,229,31,229,30,229,29,127,31,26,31,6,31,183,31,10,31,194,31,62,31,134,31,75,31,106,31,54,31,66,31,144,31,144,30,18,31,193,31,134,31,134,30,63,31,63,30,63,29,234,31,229,31,251,31,57,31,71,31,22,31,22,30,22,29,30,31,30,30,113,31,192,31,15,31,153,31,182,31,115,31,174,31,198,31,223,31,223,30,69,31,215,31,154,31,58,31,42,31,4,31,4,30,206,31,206,30,206,29,206,28,106,31,111,31,111,30,155,31,233,31,205,31,111,31,111,30,74,31,103,31,103,30,103,29,187,31,171,31,108,31,108,30,4,31,250,31,190,31,140,31,239,31,222,31,248,31,248,30,214,31,45,31,45,30,45,29,129,31,129,30,129,29,86,31,137,31,72,31,120,31,195,31,49,31,182,31,230,31,147,31,119,31,147,31,95,31,147,31,109,31,201,31,131,31,168,31,168,30,43,31,53,31,101,31,35,31,35,30,87,31,27,31,27,30,27,29,177,31,177,30,177,29,95,31,174,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
