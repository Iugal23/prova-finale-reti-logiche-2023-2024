-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 978;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (1,0,71,0,0,0,0,0,0,0,98,0,177,0,163,0,71,0,143,0,55,0,0,0,0,0,96,0,14,0,4,0,211,0,0,0,69,0,156,0,97,0,76,0,0,0,131,0,0,0,17,0,148,0,34,0,41,0,82,0,226,0,81,0,210,0,1,0,170,0,169,0,8,0,138,0,209,0,222,0,15,0,190,0,0,0,0,0,131,0,188,0,203,0,70,0,0,0,101,0,0,0,73,0,102,0,158,0,129,0,240,0,150,0,160,0,58,0,0,0,217,0,118,0,201,0,49,0,210,0,252,0,125,0,0,0,205,0,37,0,94,0,18,0,89,0,0,0,198,0,222,0,52,0,7,0,237,0,229,0,11,0,220,0,48,0,45,0,44,0,16,0,47,0,0,0,29,0,18,0,50,0,20,0,0,0,172,0,140,0,240,0,119,0,0,0,69,0,72,0,0,0,174,0,215,0,237,0,244,0,143,0,195,0,202,0,198,0,26,0,76,0,89,0,0,0,34,0,109,0,87,0,251,0,71,0,18,0,208,0,146,0,37,0,183,0,146,0,0,0,0,0,142,0,174,0,52,0,197,0,159,0,56,0,149,0,120,0,27,0,0,0,241,0,142,0,78,0,237,0,186,0,229,0,167,0,6,0,0,0,2,0,35,0,11,0,110,0,0,0,212,0,97,0,113,0,251,0,89,0,59,0,0,0,184,0,222,0,8,0,232,0,111,0,140,0,182,0,164,0,15,0,12,0,0,0,29,0,239,0,94,0,60,0,237,0,182,0,80,0,204,0,171,0,0,0,248,0,101,0,129,0,11,0,76,0,158,0,0,0,69,0,155,0,53,0,166,0,184,0,0,0,33,0,197,0,230,0,235,0,0,0,0,0,0,0,61,0,184,0,0,0,0,0,39,0,244,0,136,0,159,0,3,0,72,0,131,0,0,0,0,0,16,0,34,0,164,0,18,0,62,0,248,0,205,0,202,0,0,0,110,0,8,0,86,0,129,0,54,0,0,0,86,0,96,0,239,0,176,0,107,0,0,0,105,0,32,0,87,0,0,0,0,0,0,0,207,0,0,0,124,0,191,0,0,0,77,0,152,0,239,0,47,0,131,0,230,0,113,0,199,0,118,0,155,0,134,0,0,0,134,0,0,0,43,0,207,0,0,0,173,0,40,0,0,0,70,0,233,0,118,0,119,0,42,0,44,0,105,0,0,0,20,0,40,0,4,0,149,0,75,0,79,0,39,0,220,0,44,0,109,0,0,0,216,0,251,0,0,0,141,0,71,0,34,0,201,0,40,0,51,0,218,0,109,0,0,0,0,0,74,0,69,0,133,0,0,0,0,0,185,0,243,0,44,0,157,0,154,0,252,0,55,0,211,0,119,0,230,0,252,0,0,0,116,0,38,0,133,0,236,0,122,0,0,0,227,0,194,0,48,0,0,0,183,0,114,0,179,0,0,0,96,0,138,0,202,0,32,0,158,0,243,0,217,0,244,0,156,0,183,0,131,0,106,0,0,0,209,0,181,0,220,0,8,0,62,0,80,0,43,0,0,0,63,0,107,0,0,0,126,0,175,0,0,0,209,0,251,0,200,0,233,0,196,0,0,0,0,0,104,0,0,0,197,0,168,0,72,0,124,0,15,0,49,0,204,0,58,0,230,0,190,0,142,0,131,0,134,0,25,0,113,0,141,0,51,0,40,0,42,0,161,0,223,0,86,0,12,0,58,0,0,0,74,0,97,0,0,0,0,0,0,0,159,0,156,0,25,0,1,0,0,0,91,0,17,0,186,0,114,0,191,0,0,0,218,0,0,0,193,0,50,0,23,0,67,0,164,0,10,0,93,0,200,0,240,0,0,0,235,0,76,0,113,0,0,0,23,0,224,0,111,0,0,0,0,0,12,0,170,0,152,0,76,0,197,0,51,0,121,0,233,0,27,0,255,0,4,0,0,0,121,0,33,0,156,0,176,0,242,0,1,0,77,0,62,0,47,0,0,0,0,0,63,0,203,0,0,0,91,0,6,0,40,0,135,0,127,0,0,0,118,0,10,0,235,0,163,0,152,0,217,0,249,0,5,0,176,0,0,0,73,0,166,0,8,0,0,0,211,0,134,0,230,0,0,0,226,0,110,0,0,0,60,0,161,0,230,0,225,0,183,0,136,0,203,0,22,0,225,0,177,0,30,0,255,0,0,0,103,0,23,0,152,0,169,0,191,0,175,0,165,0,248,0,217,0,210,0,166,0,250,0,105,0,168,0,218,0,179,0,211,0,0,0,81,0,216,0,61,0,120,0,169,0,103,0,232,0,107,0,0,0,81,0,0,0,0,0,66,0,199,0,12,0,34,0,9,0,199,0,250,0,0,0,152,0,222,0,198,0,0,0,0,0,214,0,75,0,0,0,0,0,0,0,74,0,223,0,21,0,142,0,0,0,0,0,165,0,176,0,0,0,188,0,0,0,240,0,3,0,237,0,179,0,48,0,70,0,122,0,192,0,0,0,114,0,97,0,156,0,0,0,28,0,194,0,0,0,84,0,222,0,0,0,213,0,68,0,101,0,234,0,73,0,25,0,215,0,0,0,72,0,179,0,38,0,141,0,143,0,85,0,186,0,212,0,206,0,207,0,0,0,0,0,193,0,70,0,166,0,87,0,44,0,22,0,40,0,58,0,142,0,52,0,112,0,198,0,0,0,38,0,132,0,96,0,157,0,192,0,28,0,0,0,208,0,0,0,0,0,65,0,175,0,107,0,0,0,255,0,35,0,67,0,94,0,100,0,0,0,144,0,61,0,224,0,174,0,59,0,204,0,94,0,242,0,0,0,148,0,147,0,37,0,0,0,0,0,60,0,49,0,0,0,224,0,85,0,243,0,160,0,51,0,173,0,0,0,159,0,188,0,102,0,138,0,106,0,70,0,62,0,79,0,84,0,0,0,245,0,227,0,0,0,28,0,0,0,12,0,49,0,141,0,238,0,95,0,249,0,61,0,191,0,239,0,245,0,23,0,60,0,113,0,71,0,116,0,26,0,68,0,0,0,236,0,98,0,0,0,88,0,254,0,168,0,193,0,126,0,83,0,72,0,0,0,0,0,33,0,80,0,0,0,250,0,245,0,49,0,200,0,11,0,74,0,218,0,41,0,0,0,130,0,120,0,193,0,72,0,134,0,70,0,0,0,94,0,0,0,124,0,0,0,144,0,44,0,53,0,45,0,213,0,171,0,207,0,77,0,253,0,46,0,81,0,85,0,62,0,52,0,0,0,19,0,225,0,110,0,221,0,0,0,89,0,206,0,28,0,128,0,69,0,39,0,128,0,0,0,250,0,0,0,0,0,115,0,54,0,113,0,0,0,0,0,165,0,225,0,20,0,0,0,0,0,82,0,139,0,160,0,204,0,0,0,0,0,175,0,201,0,47,0,66,0,0,0,115,0,34,0,218,0,248,0,201,0,102,0,67,0,210,0,181,0,0,0,132,0,192,0,49,0,0,0,16,0,216,0,0,0,36,0,106,0,156,0,0,0,113,0,225,0,240,0,205,0,142,0,189,0,225,0,0,0,25,0,0,0,102,0,0,0,62,0,88,0,202,0,79,0,220,0,0,0,251,0,93,0,118,0,231,0,46,0,106,0,174,0,154,0,172,0,72,0,0,0,12,0,214,0,84,0,0,0,0,0,165,0,0,0,169,0,215,0,39,0,172,0,11,0,187,0,169,0,109,0,8,0,85,0,20,0,0,0,248,0,254,0,239,0,0,0,82,0,55,0,0,0,241,0,40,0,8,0,153,0,41,0,212,0,0,0,167,0,247,0,175,0,184,0,50,0,166,0,221,0,81,0,208,0,0,0,57,0,160,0,0,0,162,0,0,0,0,0,10,0,224,0,0,0,223,0,245,0,162,0,247,0,0,0,16,0,0,0,239,0,98,0,148,0,246,0,54,0,75,0,130,0,96,0,0,0,0,0,108,0,10,0,0,0,0,0,25,0,0,0,0,0,185,0,0,0,225,0,214,0,59,0,218,0,0,0,0,0,4,0,108,0,0,0,62,0,151,0,71,0,107,0,43,0,195,0,0,0,0,0,191,0,30,0,231,0,0,0,0,0,165,0,129,0,0,0,2,0,0,0,0,0,8,0,147,0,0,0,0,0,192,0,53,0,147,0,187,0,130,0,0,0,44,0,135,0,50,0,85,0,173,0,154,0,48,0,238,0,0,0,224,0,128,0,222,0,126,0,221,0,237,0,248,0,0,0,0,0,133,0,43,0,112,0,55,0,0,0,136,0,109,0,0,0,0,0,133,0,203,0,11,0,123,0,2,0,153,0,0,0,151,0,117,0,154,0,227,0,201,0,0,0,54,0,83,0,0,0,0,0,230,0,178,0,140,0);
signal scenario_full  : scenario_type := (1,31,71,31,71,30,71,29,71,28,98,31,177,31,163,31,71,31,143,31,55,31,55,30,55,29,96,31,14,31,4,31,211,31,211,30,69,31,156,31,97,31,76,31,76,30,131,31,131,30,17,31,148,31,34,31,41,31,82,31,226,31,81,31,210,31,1,31,170,31,169,31,8,31,138,31,209,31,222,31,15,31,190,31,190,30,190,29,131,31,188,31,203,31,70,31,70,30,101,31,101,30,73,31,102,31,158,31,129,31,240,31,150,31,160,31,58,31,58,30,217,31,118,31,201,31,49,31,210,31,252,31,125,31,125,30,205,31,37,31,94,31,18,31,89,31,89,30,198,31,222,31,52,31,7,31,237,31,229,31,11,31,220,31,48,31,45,31,44,31,16,31,47,31,47,30,29,31,18,31,50,31,20,31,20,30,172,31,140,31,240,31,119,31,119,30,69,31,72,31,72,30,174,31,215,31,237,31,244,31,143,31,195,31,202,31,198,31,26,31,76,31,89,31,89,30,34,31,109,31,87,31,251,31,71,31,18,31,208,31,146,31,37,31,183,31,146,31,146,30,146,29,142,31,174,31,52,31,197,31,159,31,56,31,149,31,120,31,27,31,27,30,241,31,142,31,78,31,237,31,186,31,229,31,167,31,6,31,6,30,2,31,35,31,11,31,110,31,110,30,212,31,97,31,113,31,251,31,89,31,59,31,59,30,184,31,222,31,8,31,232,31,111,31,140,31,182,31,164,31,15,31,12,31,12,30,29,31,239,31,94,31,60,31,237,31,182,31,80,31,204,31,171,31,171,30,248,31,101,31,129,31,11,31,76,31,158,31,158,30,69,31,155,31,53,31,166,31,184,31,184,30,33,31,197,31,230,31,235,31,235,30,235,29,235,28,61,31,184,31,184,30,184,29,39,31,244,31,136,31,159,31,3,31,72,31,131,31,131,30,131,29,16,31,34,31,164,31,18,31,62,31,248,31,205,31,202,31,202,30,110,31,8,31,86,31,129,31,54,31,54,30,86,31,96,31,239,31,176,31,107,31,107,30,105,31,32,31,87,31,87,30,87,29,87,28,207,31,207,30,124,31,191,31,191,30,77,31,152,31,239,31,47,31,131,31,230,31,113,31,199,31,118,31,155,31,134,31,134,30,134,31,134,30,43,31,207,31,207,30,173,31,40,31,40,30,70,31,233,31,118,31,119,31,42,31,44,31,105,31,105,30,20,31,40,31,4,31,149,31,75,31,79,31,39,31,220,31,44,31,109,31,109,30,216,31,251,31,251,30,141,31,71,31,34,31,201,31,40,31,51,31,218,31,109,31,109,30,109,29,74,31,69,31,133,31,133,30,133,29,185,31,243,31,44,31,157,31,154,31,252,31,55,31,211,31,119,31,230,31,252,31,252,30,116,31,38,31,133,31,236,31,122,31,122,30,227,31,194,31,48,31,48,30,183,31,114,31,179,31,179,30,96,31,138,31,202,31,32,31,158,31,243,31,217,31,244,31,156,31,183,31,131,31,106,31,106,30,209,31,181,31,220,31,8,31,62,31,80,31,43,31,43,30,63,31,107,31,107,30,126,31,175,31,175,30,209,31,251,31,200,31,233,31,196,31,196,30,196,29,104,31,104,30,197,31,168,31,72,31,124,31,15,31,49,31,204,31,58,31,230,31,190,31,142,31,131,31,134,31,25,31,113,31,141,31,51,31,40,31,42,31,161,31,223,31,86,31,12,31,58,31,58,30,74,31,97,31,97,30,97,29,97,28,159,31,156,31,25,31,1,31,1,30,91,31,17,31,186,31,114,31,191,31,191,30,218,31,218,30,193,31,50,31,23,31,67,31,164,31,10,31,93,31,200,31,240,31,240,30,235,31,76,31,113,31,113,30,23,31,224,31,111,31,111,30,111,29,12,31,170,31,152,31,76,31,197,31,51,31,121,31,233,31,27,31,255,31,4,31,4,30,121,31,33,31,156,31,176,31,242,31,1,31,77,31,62,31,47,31,47,30,47,29,63,31,203,31,203,30,91,31,6,31,40,31,135,31,127,31,127,30,118,31,10,31,235,31,163,31,152,31,217,31,249,31,5,31,176,31,176,30,73,31,166,31,8,31,8,30,211,31,134,31,230,31,230,30,226,31,110,31,110,30,60,31,161,31,230,31,225,31,183,31,136,31,203,31,22,31,225,31,177,31,30,31,255,31,255,30,103,31,23,31,152,31,169,31,191,31,175,31,165,31,248,31,217,31,210,31,166,31,250,31,105,31,168,31,218,31,179,31,211,31,211,30,81,31,216,31,61,31,120,31,169,31,103,31,232,31,107,31,107,30,81,31,81,30,81,29,66,31,199,31,12,31,34,31,9,31,199,31,250,31,250,30,152,31,222,31,198,31,198,30,198,29,214,31,75,31,75,30,75,29,75,28,74,31,223,31,21,31,142,31,142,30,142,29,165,31,176,31,176,30,188,31,188,30,240,31,3,31,237,31,179,31,48,31,70,31,122,31,192,31,192,30,114,31,97,31,156,31,156,30,28,31,194,31,194,30,84,31,222,31,222,30,213,31,68,31,101,31,234,31,73,31,25,31,215,31,215,30,72,31,179,31,38,31,141,31,143,31,85,31,186,31,212,31,206,31,207,31,207,30,207,29,193,31,70,31,166,31,87,31,44,31,22,31,40,31,58,31,142,31,52,31,112,31,198,31,198,30,38,31,132,31,96,31,157,31,192,31,28,31,28,30,208,31,208,30,208,29,65,31,175,31,107,31,107,30,255,31,35,31,67,31,94,31,100,31,100,30,144,31,61,31,224,31,174,31,59,31,204,31,94,31,242,31,242,30,148,31,147,31,37,31,37,30,37,29,60,31,49,31,49,30,224,31,85,31,243,31,160,31,51,31,173,31,173,30,159,31,188,31,102,31,138,31,106,31,70,31,62,31,79,31,84,31,84,30,245,31,227,31,227,30,28,31,28,30,12,31,49,31,141,31,238,31,95,31,249,31,61,31,191,31,239,31,245,31,23,31,60,31,113,31,71,31,116,31,26,31,68,31,68,30,236,31,98,31,98,30,88,31,254,31,168,31,193,31,126,31,83,31,72,31,72,30,72,29,33,31,80,31,80,30,250,31,245,31,49,31,200,31,11,31,74,31,218,31,41,31,41,30,130,31,120,31,193,31,72,31,134,31,70,31,70,30,94,31,94,30,124,31,124,30,144,31,44,31,53,31,45,31,213,31,171,31,207,31,77,31,253,31,46,31,81,31,85,31,62,31,52,31,52,30,19,31,225,31,110,31,221,31,221,30,89,31,206,31,28,31,128,31,69,31,39,31,128,31,128,30,250,31,250,30,250,29,115,31,54,31,113,31,113,30,113,29,165,31,225,31,20,31,20,30,20,29,82,31,139,31,160,31,204,31,204,30,204,29,175,31,201,31,47,31,66,31,66,30,115,31,34,31,218,31,248,31,201,31,102,31,67,31,210,31,181,31,181,30,132,31,192,31,49,31,49,30,16,31,216,31,216,30,36,31,106,31,156,31,156,30,113,31,225,31,240,31,205,31,142,31,189,31,225,31,225,30,25,31,25,30,102,31,102,30,62,31,88,31,202,31,79,31,220,31,220,30,251,31,93,31,118,31,231,31,46,31,106,31,174,31,154,31,172,31,72,31,72,30,12,31,214,31,84,31,84,30,84,29,165,31,165,30,169,31,215,31,39,31,172,31,11,31,187,31,169,31,109,31,8,31,85,31,20,31,20,30,248,31,254,31,239,31,239,30,82,31,55,31,55,30,241,31,40,31,8,31,153,31,41,31,212,31,212,30,167,31,247,31,175,31,184,31,50,31,166,31,221,31,81,31,208,31,208,30,57,31,160,31,160,30,162,31,162,30,162,29,10,31,224,31,224,30,223,31,245,31,162,31,247,31,247,30,16,31,16,30,239,31,98,31,148,31,246,31,54,31,75,31,130,31,96,31,96,30,96,29,108,31,10,31,10,30,10,29,25,31,25,30,25,29,185,31,185,30,225,31,214,31,59,31,218,31,218,30,218,29,4,31,108,31,108,30,62,31,151,31,71,31,107,31,43,31,195,31,195,30,195,29,191,31,30,31,231,31,231,30,231,29,165,31,129,31,129,30,2,31,2,30,2,29,8,31,147,31,147,30,147,29,192,31,53,31,147,31,187,31,130,31,130,30,44,31,135,31,50,31,85,31,173,31,154,31,48,31,238,31,238,30,224,31,128,31,222,31,126,31,221,31,237,31,248,31,248,30,248,29,133,31,43,31,112,31,55,31,55,30,136,31,109,31,109,30,109,29,133,31,203,31,11,31,123,31,2,31,153,31,153,30,151,31,117,31,154,31,227,31,201,31,201,30,54,31,83,31,83,30,83,29,230,31,178,31,140,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
