-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_343 is
end project_tb_343;

architecture project_tb_arch_343 of project_tb_343 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 221;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (21,0,117,0,63,0,212,0,55,0,155,0,0,0,0,0,0,0,147,0,0,0,78,0,178,0,121,0,0,0,65,0,100,0,10,0,18,0,96,0,247,0,0,0,0,0,82,0,134,0,0,0,141,0,112,0,184,0,206,0,19,0,64,0,146,0,99,0,73,0,0,0,16,0,90,0,73,0,248,0,72,0,29,0,220,0,195,0,252,0,55,0,108,0,50,0,15,0,81,0,100,0,0,0,24,0,0,0,0,0,241,0,99,0,4,0,127,0,0,0,0,0,49,0,0,0,212,0,192,0,0,0,0,0,0,0,204,0,169,0,44,0,0,0,64,0,0,0,111,0,18,0,208,0,0,0,126,0,192,0,84,0,228,0,213,0,0,0,185,0,0,0,37,0,106,0,48,0,228,0,101,0,221,0,175,0,223,0,67,0,58,0,0,0,65,0,187,0,31,0,164,0,46,0,118,0,0,0,186,0,0,0,160,0,0,0,214,0,121,0,213,0,36,0,53,0,227,0,0,0,10,0,0,0,218,0,192,0,66,0,82,0,0,0,12,0,188,0,77,0,0,0,216,0,0,0,63,0,226,0,12,0,170,0,0,0,84,0,229,0,146,0,0,0,0,0,244,0,82,0,0,0,159,0,45,0,0,0,107,0,47,0,26,0,19,0,218,0,134,0,0,0,71,0,114,0,0,0,220,0,27,0,201,0,90,0,0,0,132,0,98,0,100,0,0,0,61,0,221,0,0,0,102,0,0,0,0,0,0,0,152,0,252,0,124,0,139,0,196,0,64,0,175,0,21,0,124,0,8,0,39,0,69,0,39,0,153,0,170,0,81,0,225,0,127,0,77,0,0,0,136,0,37,0,0,0,188,0,23,0,0,0,147,0,0,0,0,0,61,0,155,0,235,0,183,0,50,0,98,0,0,0,60,0,1,0,244,0,97,0,187,0,28,0,100,0,127,0,132,0,192,0,34,0,133,0,0,0,123,0,251,0);
signal scenario_full  : scenario_type := (21,31,117,31,63,31,212,31,55,31,155,31,155,30,155,29,155,28,147,31,147,30,78,31,178,31,121,31,121,30,65,31,100,31,10,31,18,31,96,31,247,31,247,30,247,29,82,31,134,31,134,30,141,31,112,31,184,31,206,31,19,31,64,31,146,31,99,31,73,31,73,30,16,31,90,31,73,31,248,31,72,31,29,31,220,31,195,31,252,31,55,31,108,31,50,31,15,31,81,31,100,31,100,30,24,31,24,30,24,29,241,31,99,31,4,31,127,31,127,30,127,29,49,31,49,30,212,31,192,31,192,30,192,29,192,28,204,31,169,31,44,31,44,30,64,31,64,30,111,31,18,31,208,31,208,30,126,31,192,31,84,31,228,31,213,31,213,30,185,31,185,30,37,31,106,31,48,31,228,31,101,31,221,31,175,31,223,31,67,31,58,31,58,30,65,31,187,31,31,31,164,31,46,31,118,31,118,30,186,31,186,30,160,31,160,30,214,31,121,31,213,31,36,31,53,31,227,31,227,30,10,31,10,30,218,31,192,31,66,31,82,31,82,30,12,31,188,31,77,31,77,30,216,31,216,30,63,31,226,31,12,31,170,31,170,30,84,31,229,31,146,31,146,30,146,29,244,31,82,31,82,30,159,31,45,31,45,30,107,31,47,31,26,31,19,31,218,31,134,31,134,30,71,31,114,31,114,30,220,31,27,31,201,31,90,31,90,30,132,31,98,31,100,31,100,30,61,31,221,31,221,30,102,31,102,30,102,29,102,28,152,31,252,31,124,31,139,31,196,31,64,31,175,31,21,31,124,31,8,31,39,31,69,31,39,31,153,31,170,31,81,31,225,31,127,31,77,31,77,30,136,31,37,31,37,30,188,31,23,31,23,30,147,31,147,30,147,29,61,31,155,31,235,31,183,31,50,31,98,31,98,30,60,31,1,31,244,31,97,31,187,31,28,31,100,31,127,31,132,31,192,31,34,31,133,31,133,30,123,31,251,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
