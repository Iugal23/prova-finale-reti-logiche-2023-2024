-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_131 is
end project_tb_131;

architecture project_tb_arch_131 of project_tb_131 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 695;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (198,0,0,0,66,0,115,0,163,0,118,0,0,0,0,0,43,0,165,0,11,0,47,0,121,0,0,0,148,0,153,0,147,0,89,0,7,0,142,0,249,0,255,0,0,0,0,0,158,0,0,0,76,0,219,0,0,0,144,0,0,0,193,0,163,0,219,0,249,0,34,0,64,0,18,0,255,0,32,0,222,0,133,0,226,0,17,0,0,0,175,0,0,0,0,0,244,0,0,0,68,0,130,0,58,0,0,0,245,0,150,0,36,0,8,0,203,0,247,0,178,0,0,0,80,0,130,0,0,0,147,0,223,0,5,0,201,0,56,0,0,0,187,0,230,0,198,0,222,0,212,0,201,0,213,0,174,0,33,0,23,0,108,0,17,0,210,0,0,0,0,0,0,0,76,0,128,0,149,0,120,0,172,0,43,0,104,0,0,0,0,0,152,0,0,0,0,0,163,0,0,0,5,0,25,0,99,0,42,0,39,0,0,0,128,0,0,0,35,0,224,0,0,0,147,0,148,0,45,0,179,0,141,0,176,0,82,0,204,0,79,0,0,0,121,0,231,0,235,0,6,0,161,0,11,0,28,0,95,0,0,0,245,0,126,0,0,0,0,0,0,0,1,0,207,0,0,0,249,0,5,0,126,0,130,0,0,0,159,0,78,0,0,0,113,0,155,0,158,0,49,0,138,0,128,0,118,0,0,0,4,0,0,0,101,0,184,0,0,0,130,0,230,0,0,0,204,0,201,0,0,0,150,0,128,0,128,0,79,0,15,0,243,0,171,0,189,0,200,0,0,0,24,0,118,0,102,0,157,0,0,0,0,0,3,0,47,0,0,0,164,0,64,0,0,0,190,0,0,0,1,0,0,0,130,0,0,0,0,0,224,0,0,0,209,0,140,0,29,0,55,0,53,0,184,0,244,0,174,0,133,0,184,0,0,0,205,0,46,0,25,0,184,0,148,0,243,0,0,0,128,0,78,0,75,0,138,0,107,0,11,0,174,0,116,0,128,0,0,0,0,0,244,0,0,0,0,0,24,0,69,0,116,0,0,0,166,0,186,0,183,0,76,0,200,0,240,0,107,0,5,0,19,0,88,0,133,0,183,0,241,0,199,0,113,0,91,0,87,0,40,0,154,0,40,0,66,0,97,0,175,0,208,0,0,0,190,0,0,0,89,0,127,0,214,0,168,0,199,0,87,0,38,0,169,0,1,0,13,0,0,0,0,0,0,0,208,0,255,0,215,0,86,0,244,0,43,0,2,0,151,0,119,0,50,0,68,0,56,0,90,0,186,0,0,0,0,0,0,0,208,0,0,0,143,0,53,0,94,0,149,0,0,0,182,0,61,0,107,0,255,0,117,0,224,0,0,0,0,0,0,0,0,0,104,0,0,0,249,0,0,0,14,0,50,0,27,0,0,0,0,0,250,0,162,0,6,0,204,0,250,0,134,0,232,0,105,0,142,0,39,0,93,0,180,0,131,0,106,0,226,0,167,0,36,0,177,0,81,0,115,0,63,0,40,0,69,0,131,0,145,0,146,0,170,0,210,0,0,0,173,0,246,0,174,0,203,0,0,0,152,0,207,0,153,0,41,0,107,0,243,0,230,0,189,0,189,0,166,0,212,0,135,0,33,0,182,0,129,0,141,0,89,0,126,0,61,0,70,0,0,0,194,0,173,0,10,0,0,0,0,0,0,0,198,0,39,0,143,0,9,0,163,0,0,0,17,0,119,0,190,0,0,0,180,0,0,0,2,0,228,0,0,0,0,0,12,0,236,0,240,0,0,0,0,0,68,0,48,0,0,0,19,0,0,0,41,0,0,0,99,0,239,0,78,0,4,0,68,0,251,0,255,0,0,0,198,0,0,0,13,0,149,0,199,0,213,0,17,0,248,0,0,0,0,0,183,0,203,0,0,0,178,0,138,0,114,0,0,0,23,0,0,0,27,0,46,0,129,0,226,0,85,0,0,0,0,0,161,0,192,0,89,0,0,0,151,0,126,0,37,0,158,0,175,0,43,0,38,0,0,0,60,0,216,0,0,0,116,0,228,0,205,0,14,0,127,0,158,0,250,0,169,0,122,0,0,0,253,0,84,0,129,0,62,0,183,0,82,0,134,0,35,0,212,0,188,0,142,0,34,0,138,0,0,0,79,0,206,0,162,0,42,0,1,0,143,0,39,0,234,0,123,0,69,0,12,0,0,0,37,0,250,0,0,0,149,0,10,0,142,0,159,0,0,0,69,0,37,0,104,0,0,0,0,0,240,0,78,0,13,0,76,0,60,0,78,0,247,0,16,0,0,0,68,0,16,0,249,0,240,0,45,0,103,0,168,0,182,0,177,0,0,0,207,0,93,0,166,0,160,0,255,0,0,0,241,0,0,0,255,0,63,0,0,0,203,0,163,0,0,0,144,0,0,0,0,0,229,0,9,0,130,0,49,0,165,0,62,0,21,0,85,0,61,0,210,0,95,0,32,0,117,0,0,0,176,0,116,0,40,0,146,0,226,0,72,0,225,0,82,0,9,0,27,0,0,0,0,0,188,0,0,0,104,0,0,0,194,0,215,0,0,0,234,0,66,0,98,0,115,0,0,0,253,0,146,0,14,0,212,0,49,0,151,0,18,0,129,0,100,0,105,0,233,0,169,0,137,0,219,0,80,0,74,0,195,0,71,0,0,0,0,0,140,0,209,0,233,0,61,0,188,0,216,0,0,0,18,0,86,0,206,0,106,0,187,0,0,0,194,0,87,0,44,0,252,0,118,0,145,0,118,0,234,0,125,0,130,0,240,0,13,0,0,0,77,0,67,0,79,0,81,0,216,0,13,0,200,0,35,0,225,0,0,0,6,0,156,0,0,0,130,0,6,0,106,0,3,0,229,0,118,0,0,0,205,0,89,0,132,0,0,0,251,0,176,0,200,0,0,0,165,0,55,0,107,0,0,0,99,0,24,0,0,0,198,0,0,0,51,0,0,0,251,0,87,0,35,0,3,0,167,0,230,0,81,0,10,0,116,0,92,0,66,0,12,0,0,0,141,0,42,0,163,0,61,0,0,0,98,0,168,0,13,0,157,0,83,0,120,0,0,0,196,0,235,0,206,0,0,0,46,0,163,0,29,0,8,0);
signal scenario_full  : scenario_type := (198,31,198,30,66,31,115,31,163,31,118,31,118,30,118,29,43,31,165,31,11,31,47,31,121,31,121,30,148,31,153,31,147,31,89,31,7,31,142,31,249,31,255,31,255,30,255,29,158,31,158,30,76,31,219,31,219,30,144,31,144,30,193,31,163,31,219,31,249,31,34,31,64,31,18,31,255,31,32,31,222,31,133,31,226,31,17,31,17,30,175,31,175,30,175,29,244,31,244,30,68,31,130,31,58,31,58,30,245,31,150,31,36,31,8,31,203,31,247,31,178,31,178,30,80,31,130,31,130,30,147,31,223,31,5,31,201,31,56,31,56,30,187,31,230,31,198,31,222,31,212,31,201,31,213,31,174,31,33,31,23,31,108,31,17,31,210,31,210,30,210,29,210,28,76,31,128,31,149,31,120,31,172,31,43,31,104,31,104,30,104,29,152,31,152,30,152,29,163,31,163,30,5,31,25,31,99,31,42,31,39,31,39,30,128,31,128,30,35,31,224,31,224,30,147,31,148,31,45,31,179,31,141,31,176,31,82,31,204,31,79,31,79,30,121,31,231,31,235,31,6,31,161,31,11,31,28,31,95,31,95,30,245,31,126,31,126,30,126,29,126,28,1,31,207,31,207,30,249,31,5,31,126,31,130,31,130,30,159,31,78,31,78,30,113,31,155,31,158,31,49,31,138,31,128,31,118,31,118,30,4,31,4,30,101,31,184,31,184,30,130,31,230,31,230,30,204,31,201,31,201,30,150,31,128,31,128,31,79,31,15,31,243,31,171,31,189,31,200,31,200,30,24,31,118,31,102,31,157,31,157,30,157,29,3,31,47,31,47,30,164,31,64,31,64,30,190,31,190,30,1,31,1,30,130,31,130,30,130,29,224,31,224,30,209,31,140,31,29,31,55,31,53,31,184,31,244,31,174,31,133,31,184,31,184,30,205,31,46,31,25,31,184,31,148,31,243,31,243,30,128,31,78,31,75,31,138,31,107,31,11,31,174,31,116,31,128,31,128,30,128,29,244,31,244,30,244,29,24,31,69,31,116,31,116,30,166,31,186,31,183,31,76,31,200,31,240,31,107,31,5,31,19,31,88,31,133,31,183,31,241,31,199,31,113,31,91,31,87,31,40,31,154,31,40,31,66,31,97,31,175,31,208,31,208,30,190,31,190,30,89,31,127,31,214,31,168,31,199,31,87,31,38,31,169,31,1,31,13,31,13,30,13,29,13,28,208,31,255,31,215,31,86,31,244,31,43,31,2,31,151,31,119,31,50,31,68,31,56,31,90,31,186,31,186,30,186,29,186,28,208,31,208,30,143,31,53,31,94,31,149,31,149,30,182,31,61,31,107,31,255,31,117,31,224,31,224,30,224,29,224,28,224,27,104,31,104,30,249,31,249,30,14,31,50,31,27,31,27,30,27,29,250,31,162,31,6,31,204,31,250,31,134,31,232,31,105,31,142,31,39,31,93,31,180,31,131,31,106,31,226,31,167,31,36,31,177,31,81,31,115,31,63,31,40,31,69,31,131,31,145,31,146,31,170,31,210,31,210,30,173,31,246,31,174,31,203,31,203,30,152,31,207,31,153,31,41,31,107,31,243,31,230,31,189,31,189,31,166,31,212,31,135,31,33,31,182,31,129,31,141,31,89,31,126,31,61,31,70,31,70,30,194,31,173,31,10,31,10,30,10,29,10,28,198,31,39,31,143,31,9,31,163,31,163,30,17,31,119,31,190,31,190,30,180,31,180,30,2,31,228,31,228,30,228,29,12,31,236,31,240,31,240,30,240,29,68,31,48,31,48,30,19,31,19,30,41,31,41,30,99,31,239,31,78,31,4,31,68,31,251,31,255,31,255,30,198,31,198,30,13,31,149,31,199,31,213,31,17,31,248,31,248,30,248,29,183,31,203,31,203,30,178,31,138,31,114,31,114,30,23,31,23,30,27,31,46,31,129,31,226,31,85,31,85,30,85,29,161,31,192,31,89,31,89,30,151,31,126,31,37,31,158,31,175,31,43,31,38,31,38,30,60,31,216,31,216,30,116,31,228,31,205,31,14,31,127,31,158,31,250,31,169,31,122,31,122,30,253,31,84,31,129,31,62,31,183,31,82,31,134,31,35,31,212,31,188,31,142,31,34,31,138,31,138,30,79,31,206,31,162,31,42,31,1,31,143,31,39,31,234,31,123,31,69,31,12,31,12,30,37,31,250,31,250,30,149,31,10,31,142,31,159,31,159,30,69,31,37,31,104,31,104,30,104,29,240,31,78,31,13,31,76,31,60,31,78,31,247,31,16,31,16,30,68,31,16,31,249,31,240,31,45,31,103,31,168,31,182,31,177,31,177,30,207,31,93,31,166,31,160,31,255,31,255,30,241,31,241,30,255,31,63,31,63,30,203,31,163,31,163,30,144,31,144,30,144,29,229,31,9,31,130,31,49,31,165,31,62,31,21,31,85,31,61,31,210,31,95,31,32,31,117,31,117,30,176,31,116,31,40,31,146,31,226,31,72,31,225,31,82,31,9,31,27,31,27,30,27,29,188,31,188,30,104,31,104,30,194,31,215,31,215,30,234,31,66,31,98,31,115,31,115,30,253,31,146,31,14,31,212,31,49,31,151,31,18,31,129,31,100,31,105,31,233,31,169,31,137,31,219,31,80,31,74,31,195,31,71,31,71,30,71,29,140,31,209,31,233,31,61,31,188,31,216,31,216,30,18,31,86,31,206,31,106,31,187,31,187,30,194,31,87,31,44,31,252,31,118,31,145,31,118,31,234,31,125,31,130,31,240,31,13,31,13,30,77,31,67,31,79,31,81,31,216,31,13,31,200,31,35,31,225,31,225,30,6,31,156,31,156,30,130,31,6,31,106,31,3,31,229,31,118,31,118,30,205,31,89,31,132,31,132,30,251,31,176,31,200,31,200,30,165,31,55,31,107,31,107,30,99,31,24,31,24,30,198,31,198,30,51,31,51,30,251,31,87,31,35,31,3,31,167,31,230,31,81,31,10,31,116,31,92,31,66,31,12,31,12,30,141,31,42,31,163,31,61,31,61,30,98,31,168,31,13,31,157,31,83,31,120,31,120,30,196,31,235,31,206,31,206,30,46,31,163,31,29,31,8,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
