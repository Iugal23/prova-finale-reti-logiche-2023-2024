-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 739;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,116,0,44,0,188,0,79,0,0,0,85,0,215,0,45,0,245,0,96,0,74,0,0,0,23,0,203,0,134,0,22,0,114,0,7,0,43,0,30,0,74,0,0,0,0,0,6,0,115,0,0,0,133,0,52,0,45,0,0,0,0,0,203,0,6,0,0,0,0,0,0,0,218,0,0,0,0,0,78,0,0,0,123,0,230,0,0,0,196,0,0,0,203,0,0,0,0,0,117,0,133,0,241,0,8,0,203,0,209,0,119,0,2,0,0,0,52,0,204,0,154,0,100,0,62,0,12,0,222,0,209,0,105,0,24,0,232,0,0,0,148,0,60,0,85,0,161,0,0,0,76,0,64,0,5,0,129,0,161,0,241,0,35,0,228,0,9,0,234,0,0,0,159,0,0,0,205,0,230,0,158,0,105,0,216,0,35,0,169,0,182,0,108,0,121,0,53,0,197,0,38,0,237,0,189,0,115,0,139,0,11,0,0,0,197,0,41,0,0,0,16,0,124,0,43,0,221,0,243,0,0,0,176,0,231,0,164,0,50,0,190,0,61,0,166,0,22,0,132,0,233,0,0,0,0,0,0,0,95,0,0,0,0,0,78,0,97,0,0,0,169,0,107,0,109,0,225,0,126,0,0,0,207,0,0,0,177,0,54,0,206,0,0,0,0,0,138,0,250,0,255,0,0,0,195,0,193,0,0,0,11,0,86,0,0,0,87,0,0,0,194,0,77,0,203,0,44,0,0,0,227,0,170,0,0,0,207,0,203,0,255,0,0,0,195,0,0,0,0,0,0,0,100,0,228,0,246,0,104,0,0,0,36,0,124,0,16,0,0,0,155,0,230,0,0,0,10,0,201,0,0,0,0,0,214,0,0,0,17,0,139,0,0,0,178,0,2,0,198,0,40,0,81,0,28,0,226,0,99,0,67,0,71,0,102,0,225,0,241,0,165,0,60,0,65,0,4,0,138,0,135,0,244,0,235,0,132,0,136,0,141,0,0,0,34,0,41,0,140,0,0,0,0,0,17,0,146,0,59,0,67,0,126,0,153,0,83,0,174,0,161,0,155,0,21,0,235,0,2,0,237,0,0,0,109,0,173,0,161,0,203,0,127,0,99,0,213,0,19,0,183,0,100,0,66,0,4,0,184,0,135,0,22,0,0,0,93,0,123,0,96,0,0,0,170,0,201,0,0,0,0,0,97,0,54,0,0,0,53,0,0,0,0,0,247,0,19,0,182,0,129,0,162,0,138,0,152,0,0,0,0,0,0,0,0,0,0,0,145,0,183,0,67,0,239,0,86,0,129,0,0,0,0,0,162,0,68,0,250,0,132,0,153,0,5,0,0,0,184,0,19,0,0,0,0,0,219,0,221,0,158,0,0,0,42,0,39,0,251,0,245,0,248,0,173,0,0,0,250,0,114,0,0,0,0,0,134,0,95,0,162,0,4,0,0,0,75,0,247,0,197,0,183,0,0,0,0,0,111,0,122,0,246,0,208,0,217,0,145,0,231,0,24,0,181,0,7,0,0,0,0,0,247,0,55,0,0,0,66,0,64,0,0,0,126,0,63,0,49,0,95,0,248,0,0,0,219,0,0,0,130,0,189,0,170,0,244,0,127,0,24,0,251,0,245,0,195,0,65,0,54,0,181,0,0,0,60,0,147,0,0,0,78,0,205,0,230,0,203,0,137,0,46,0,91,0,166,0,0,0,77,0,177,0,5,0,157,0,84,0,163,0,125,0,152,0,87,0,6,0,63,0,105,0,15,0,144,0,105,0,211,0,0,0,44,0,201,0,0,0,35,0,43,0,2,0,254,0,5,0,169,0,180,0,0,0,102,0,119,0,247,0,43,0,0,0,135,0,170,0,99,0,26,0,62,0,207,0,205,0,0,0,140,0,240,0,0,0,0,0,0,0,0,0,109,0,0,0,226,0,0,0,66,0,74,0,192,0,0,0,118,0,58,0,0,0,137,0,0,0,166,0,58,0,228,0,29,0,232,0,29,0,0,0,68,0,154,0,52,0,116,0,195,0,135,0,0,0,68,0,0,0,0,0,84,0,209,0,114,0,176,0,117,0,182,0,102,0,82,0,35,0,221,0,186,0,0,0,82,0,225,0,65,0,220,0,141,0,208,0,141,0,0,0,169,0,0,0,210,0,142,0,84,0,112,0,161,0,1,0,233,0,118,0,0,0,18,0,195,0,213,0,63,0,96,0,38,0,127,0,50,0,228,0,61,0,2,0,0,0,0,0,0,0,0,0,246,0,0,0,193,0,0,0,0,0,74,0,24,0,0,0,13,0,41,0,25,0,0,0,49,0,206,0,223,0,162,0,0,0,0,0,169,0,78,0,6,0,0,0,142,0,0,0,74,0,24,0,15,0,233,0,93,0,8,0,28,0,229,0,145,0,122,0,111,0,140,0,61,0,131,0,231,0,0,0,0,0,186,0,46,0,167,0,4,0,29,0,207,0,39,0,96,0,94,0,221,0,185,0,192,0,52,0,0,0,241,0,33,0,229,0,103,0,60,0,120,0,0,0,56,0,133,0,0,0,135,0,0,0,82,0,226,0,29,0,26,0,228,0,104,0,160,0,103,0,195,0,0,0,82,0,45,0,195,0,0,0,195,0,71,0,249,0,252,0,72,0,59,0,113,0,0,0,19,0,89,0,88,0,143,0,236,0,208,0,115,0,186,0,0,0,184,0,147,0,159,0,76,0,161,0,147,0,0,0,219,0,0,0,0,0,58,0,128,0,122,0,20,0,4,0,119,0,18,0,184,0,0,0,30,0,0,0,0,0,17,0,245,0,0,0,173,0,231,0,245,0,227,0,85,0,194,0,215,0,202,0,164,0,91,0,19,0,101,0,52,0,26,0,30,0,11,0,0,0,190,0,0,0,195,0,87,0,244,0,31,0,69,0,228,0,117,0,122,0,124,0,0,0,101,0,202,0,22,0,74,0,99,0,208,0,249,0,192,0,78,0,252,0,177,0,48,0,158,0,213,0,23,0,34,0,214,0,244,0,36,0,174,0,100,0,75,0,237,0,162,0,106,0,76,0,0,0,143,0,183,0,0,0,59,0,77,0,97,0,203,0,230,0,174,0,42,0,221,0,79,0,0,0,152,0,0,0,245,0,44,0,11,0,0,0,83,0,218,0,105,0,188,0,107,0,164,0,0,0,206,0,152,0,105,0,35,0,42,0,29,0,189,0,190,0,167,0,153,0,201,0,115,0,103,0,27,0,118,0,0,0,176,0,184,0,0,0,27,0,233,0,115,0,20,0,6,0,0,0,0,0,23,0,119,0,146,0,223,0);
signal scenario_full  : scenario_type := (0,0,116,31,44,31,188,31,79,31,79,30,85,31,215,31,45,31,245,31,96,31,74,31,74,30,23,31,203,31,134,31,22,31,114,31,7,31,43,31,30,31,74,31,74,30,74,29,6,31,115,31,115,30,133,31,52,31,45,31,45,30,45,29,203,31,6,31,6,30,6,29,6,28,218,31,218,30,218,29,78,31,78,30,123,31,230,31,230,30,196,31,196,30,203,31,203,30,203,29,117,31,133,31,241,31,8,31,203,31,209,31,119,31,2,31,2,30,52,31,204,31,154,31,100,31,62,31,12,31,222,31,209,31,105,31,24,31,232,31,232,30,148,31,60,31,85,31,161,31,161,30,76,31,64,31,5,31,129,31,161,31,241,31,35,31,228,31,9,31,234,31,234,30,159,31,159,30,205,31,230,31,158,31,105,31,216,31,35,31,169,31,182,31,108,31,121,31,53,31,197,31,38,31,237,31,189,31,115,31,139,31,11,31,11,30,197,31,41,31,41,30,16,31,124,31,43,31,221,31,243,31,243,30,176,31,231,31,164,31,50,31,190,31,61,31,166,31,22,31,132,31,233,31,233,30,233,29,233,28,95,31,95,30,95,29,78,31,97,31,97,30,169,31,107,31,109,31,225,31,126,31,126,30,207,31,207,30,177,31,54,31,206,31,206,30,206,29,138,31,250,31,255,31,255,30,195,31,193,31,193,30,11,31,86,31,86,30,87,31,87,30,194,31,77,31,203,31,44,31,44,30,227,31,170,31,170,30,207,31,203,31,255,31,255,30,195,31,195,30,195,29,195,28,100,31,228,31,246,31,104,31,104,30,36,31,124,31,16,31,16,30,155,31,230,31,230,30,10,31,201,31,201,30,201,29,214,31,214,30,17,31,139,31,139,30,178,31,2,31,198,31,40,31,81,31,28,31,226,31,99,31,67,31,71,31,102,31,225,31,241,31,165,31,60,31,65,31,4,31,138,31,135,31,244,31,235,31,132,31,136,31,141,31,141,30,34,31,41,31,140,31,140,30,140,29,17,31,146,31,59,31,67,31,126,31,153,31,83,31,174,31,161,31,155,31,21,31,235,31,2,31,237,31,237,30,109,31,173,31,161,31,203,31,127,31,99,31,213,31,19,31,183,31,100,31,66,31,4,31,184,31,135,31,22,31,22,30,93,31,123,31,96,31,96,30,170,31,201,31,201,30,201,29,97,31,54,31,54,30,53,31,53,30,53,29,247,31,19,31,182,31,129,31,162,31,138,31,152,31,152,30,152,29,152,28,152,27,152,26,145,31,183,31,67,31,239,31,86,31,129,31,129,30,129,29,162,31,68,31,250,31,132,31,153,31,5,31,5,30,184,31,19,31,19,30,19,29,219,31,221,31,158,31,158,30,42,31,39,31,251,31,245,31,248,31,173,31,173,30,250,31,114,31,114,30,114,29,134,31,95,31,162,31,4,31,4,30,75,31,247,31,197,31,183,31,183,30,183,29,111,31,122,31,246,31,208,31,217,31,145,31,231,31,24,31,181,31,7,31,7,30,7,29,247,31,55,31,55,30,66,31,64,31,64,30,126,31,63,31,49,31,95,31,248,31,248,30,219,31,219,30,130,31,189,31,170,31,244,31,127,31,24,31,251,31,245,31,195,31,65,31,54,31,181,31,181,30,60,31,147,31,147,30,78,31,205,31,230,31,203,31,137,31,46,31,91,31,166,31,166,30,77,31,177,31,5,31,157,31,84,31,163,31,125,31,152,31,87,31,6,31,63,31,105,31,15,31,144,31,105,31,211,31,211,30,44,31,201,31,201,30,35,31,43,31,2,31,254,31,5,31,169,31,180,31,180,30,102,31,119,31,247,31,43,31,43,30,135,31,170,31,99,31,26,31,62,31,207,31,205,31,205,30,140,31,240,31,240,30,240,29,240,28,240,27,109,31,109,30,226,31,226,30,66,31,74,31,192,31,192,30,118,31,58,31,58,30,137,31,137,30,166,31,58,31,228,31,29,31,232,31,29,31,29,30,68,31,154,31,52,31,116,31,195,31,135,31,135,30,68,31,68,30,68,29,84,31,209,31,114,31,176,31,117,31,182,31,102,31,82,31,35,31,221,31,186,31,186,30,82,31,225,31,65,31,220,31,141,31,208,31,141,31,141,30,169,31,169,30,210,31,142,31,84,31,112,31,161,31,1,31,233,31,118,31,118,30,18,31,195,31,213,31,63,31,96,31,38,31,127,31,50,31,228,31,61,31,2,31,2,30,2,29,2,28,2,27,246,31,246,30,193,31,193,30,193,29,74,31,24,31,24,30,13,31,41,31,25,31,25,30,49,31,206,31,223,31,162,31,162,30,162,29,169,31,78,31,6,31,6,30,142,31,142,30,74,31,24,31,15,31,233,31,93,31,8,31,28,31,229,31,145,31,122,31,111,31,140,31,61,31,131,31,231,31,231,30,231,29,186,31,46,31,167,31,4,31,29,31,207,31,39,31,96,31,94,31,221,31,185,31,192,31,52,31,52,30,241,31,33,31,229,31,103,31,60,31,120,31,120,30,56,31,133,31,133,30,135,31,135,30,82,31,226,31,29,31,26,31,228,31,104,31,160,31,103,31,195,31,195,30,82,31,45,31,195,31,195,30,195,31,71,31,249,31,252,31,72,31,59,31,113,31,113,30,19,31,89,31,88,31,143,31,236,31,208,31,115,31,186,31,186,30,184,31,147,31,159,31,76,31,161,31,147,31,147,30,219,31,219,30,219,29,58,31,128,31,122,31,20,31,4,31,119,31,18,31,184,31,184,30,30,31,30,30,30,29,17,31,245,31,245,30,173,31,231,31,245,31,227,31,85,31,194,31,215,31,202,31,164,31,91,31,19,31,101,31,52,31,26,31,30,31,11,31,11,30,190,31,190,30,195,31,87,31,244,31,31,31,69,31,228,31,117,31,122,31,124,31,124,30,101,31,202,31,22,31,74,31,99,31,208,31,249,31,192,31,78,31,252,31,177,31,48,31,158,31,213,31,23,31,34,31,214,31,244,31,36,31,174,31,100,31,75,31,237,31,162,31,106,31,76,31,76,30,143,31,183,31,183,30,59,31,77,31,97,31,203,31,230,31,174,31,42,31,221,31,79,31,79,30,152,31,152,30,245,31,44,31,11,31,11,30,83,31,218,31,105,31,188,31,107,31,164,31,164,30,206,31,152,31,105,31,35,31,42,31,29,31,189,31,190,31,167,31,153,31,201,31,115,31,103,31,27,31,118,31,118,30,176,31,184,31,184,30,27,31,233,31,115,31,20,31,6,31,6,30,6,29,23,31,119,31,146,31,223,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
