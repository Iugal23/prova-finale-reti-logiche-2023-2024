-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 703;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (51,0,59,0,230,0,209,0,218,0,43,0,164,0,60,0,114,0,90,0,135,0,0,0,164,0,0,0,252,0,121,0,111,0,151,0,0,0,158,0,157,0,125,0,0,0,116,0,58,0,0,0,128,0,120,0,81,0,199,0,174,0,14,0,0,0,225,0,0,0,71,0,228,0,60,0,0,0,44,0,0,0,0,0,193,0,192,0,184,0,147,0,21,0,42,0,208,0,27,0,125,0,14,0,0,0,0,0,0,0,247,0,8,0,141,0,88,0,248,0,22,0,54,0,55,0,75,0,20,0,160,0,80,0,103,0,19,0,14,0,0,0,19,0,25,0,9,0,87,0,175,0,16,0,0,0,254,0,98,0,113,0,0,0,255,0,188,0,15,0,79,0,49,0,98,0,84,0,210,0,63,0,175,0,230,0,77,0,229,0,60,0,71,0,132,0,125,0,25,0,0,0,0,0,90,0,0,0,0,0,13,0,122,0,20,0,229,0,119,0,162,0,231,0,178,0,10,0,0,0,77,0,67,0,0,0,201,0,16,0,83,0,136,0,0,0,141,0,241,0,187,0,3,0,226,0,1,0,243,0,74,0,1,0,244,0,217,0,204,0,76,0,203,0,52,0,104,0,130,0,196,0,114,0,133,0,106,0,167,0,95,0,119,0,0,0,165,0,175,0,55,0,216,0,173,0,97,0,240,0,0,0,217,0,152,0,37,0,80,0,99,0,14,0,36,0,235,0,84,0,0,0,119,0,36,0,139,0,0,0,0,0,202,0,18,0,119,0,128,0,198,0,73,0,33,0,134,0,0,0,197,0,50,0,137,0,9,0,0,0,244,0,0,0,59,0,37,0,67,0,0,0,180,0,0,0,127,0,241,0,183,0,135,0,178,0,206,0,18,0,23,0,54,0,0,0,102,0,130,0,0,0,194,0,147,0,0,0,54,0,80,0,57,0,170,0,0,0,235,0,186,0,75,0,200,0,201,0,59,0,208,0,22,0,214,0,139,0,116,0,108,0,41,0,176,0,0,0,85,0,101,0,77,0,177,0,0,0,175,0,8,0,247,0,0,0,114,0,35,0,142,0,0,0,210,0,194,0,176,0,158,0,0,0,141,0,14,0,129,0,205,0,45,0,110,0,0,0,69,0,55,0,54,0,25,0,138,0,118,0,94,0,105,0,232,0,0,0,0,0,0,0,89,0,134,0,154,0,0,0,202,0,252,0,123,0,176,0,5,0,0,0,224,0,194,0,174,0,203,0,168,0,151,0,247,0,83,0,181,0,211,0,105,0,0,0,85,0,126,0,200,0,94,0,28,0,238,0,9,0,131,0,219,0,28,0,0,0,32,0,107,0,0,0,3,0,115,0,144,0,20,0,65,0,6,0,168,0,224,0,47,0,39,0,0,0,61,0,14,0,195,0,102,0,0,0,124,0,238,0,0,0,7,0,89,0,0,0,176,0,63,0,184,0,0,0,223,0,250,0,235,0,0,0,46,0,81,0,11,0,173,0,254,0,204,0,0,0,53,0,124,0,156,0,0,0,4,0,0,0,0,0,0,0,211,0,35,0,18,0,156,0,129,0,114,0,112,0,195,0,3,0,35,0,204,0,0,0,222,0,139,0,137,0,102,0,144,0,211,0,246,0,183,0,7,0,216,0,0,0,0,0,93,0,242,0,173,0,172,0,0,0,53,0,156,0,85,0,62,0,0,0,46,0,186,0,158,0,0,0,201,0,48,0,165,0,114,0,0,0,112,0,105,0,15,0,164,0,207,0,105,0,100,0,0,0,85,0,208,0,0,0,92,0,52,0,51,0,0,0,115,0,57,0,183,0,223,0,172,0,167,0,163,0,12,0,126,0,40,0,229,0,203,0,185,0,66,0,213,0,214,0,88,0,25,0,255,0,8,0,0,0,132,0,172,0,0,0,115,0,0,0,219,0,0,0,234,0,73,0,188,0,6,0,8,0,242,0,53,0,253,0,181,0,108,0,71,0,80,0,211,0,6,0,187,0,165,0,176,0,0,0,0,0,58,0,0,0,103,0,243,0,171,0,99,0,167,0,251,0,100,0,13,0,140,0,38,0,115,0,61,0,104,0,247,0,120,0,205,0,134,0,48,0,10,0,104,0,0,0,60,0,238,0,119,0,131,0,0,0,134,0,223,0,0,0,0,0,67,0,137,0,96,0,231,0,0,0,139,0,0,0,212,0,2,0,166,0,110,0,43,0,123,0,13,0,0,0,28,0,129,0,67,0,0,0,183,0,30,0,120,0,17,0,0,0,89,0,139,0,231,0,50,0,88,0,204,0,0,0,100,0,11,0,93,0,176,0,180,0,253,0,176,0,223,0,232,0,233,0,228,0,83,0,36,0,0,0,45,0,0,0,204,0,0,0,69,0,73,0,169,0,210,0,0,0,37,0,193,0,215,0,179,0,0,0,0,0,161,0,156,0,0,0,16,0,136,0,169,0,224,0,18,0,0,0,255,0,130,0,0,0,225,0,0,0,0,0,112,0,151,0,0,0,53,0,75,0,80,0,108,0,48,0,0,0,44,0,118,0,0,0,200,0,79,0,251,0,145,0,0,0,231,0,139,0,250,0,51,0,0,0,137,0,187,0,0,0,0,0,183,0,127,0,230,0,0,0,107,0,18,0,22,0,0,0,143,0,37,0,0,0,178,0,62,0,228,0,9,0,112,0,26,0,234,0,187,0,109,0,57,0,0,0,124,0,226,0,248,0,153,0,13,0,0,0,37,0,249,0,0,0,0,0,0,0,0,0,0,0,0,0,165,0,192,0,143,0,40,0,0,0,223,0,93,0,0,0,255,0,176,0,0,0,21,0,136,0,97,0,13,0,94,0,0,0,165,0,0,0,100,0,212,0,254,0,18,0,0,0,157,0,25,0,58,0,116,0,0,0,48,0,28,0,0,0,119,0,0,0,6,0,226,0,0,0,103,0,100,0,211,0,145,0,90,0,0,0,0,0,0,0,64,0,1,0,235,0,1,0,243,0,69,0,0,0,0,0,167,0,0,0,67,0,11,0,168,0,0,0,173,0,231,0,86,0,132,0,0,0,0,0,192,0,0,0,0,0,227,0,44,0,0,0,169,0,254,0,32,0,61,0,166,0,37,0,0,0,0,0,0,0,220,0,0,0);
signal scenario_full  : scenario_type := (51,31,59,31,230,31,209,31,218,31,43,31,164,31,60,31,114,31,90,31,135,31,135,30,164,31,164,30,252,31,121,31,111,31,151,31,151,30,158,31,157,31,125,31,125,30,116,31,58,31,58,30,128,31,120,31,81,31,199,31,174,31,14,31,14,30,225,31,225,30,71,31,228,31,60,31,60,30,44,31,44,30,44,29,193,31,192,31,184,31,147,31,21,31,42,31,208,31,27,31,125,31,14,31,14,30,14,29,14,28,247,31,8,31,141,31,88,31,248,31,22,31,54,31,55,31,75,31,20,31,160,31,80,31,103,31,19,31,14,31,14,30,19,31,25,31,9,31,87,31,175,31,16,31,16,30,254,31,98,31,113,31,113,30,255,31,188,31,15,31,79,31,49,31,98,31,84,31,210,31,63,31,175,31,230,31,77,31,229,31,60,31,71,31,132,31,125,31,25,31,25,30,25,29,90,31,90,30,90,29,13,31,122,31,20,31,229,31,119,31,162,31,231,31,178,31,10,31,10,30,77,31,67,31,67,30,201,31,16,31,83,31,136,31,136,30,141,31,241,31,187,31,3,31,226,31,1,31,243,31,74,31,1,31,244,31,217,31,204,31,76,31,203,31,52,31,104,31,130,31,196,31,114,31,133,31,106,31,167,31,95,31,119,31,119,30,165,31,175,31,55,31,216,31,173,31,97,31,240,31,240,30,217,31,152,31,37,31,80,31,99,31,14,31,36,31,235,31,84,31,84,30,119,31,36,31,139,31,139,30,139,29,202,31,18,31,119,31,128,31,198,31,73,31,33,31,134,31,134,30,197,31,50,31,137,31,9,31,9,30,244,31,244,30,59,31,37,31,67,31,67,30,180,31,180,30,127,31,241,31,183,31,135,31,178,31,206,31,18,31,23,31,54,31,54,30,102,31,130,31,130,30,194,31,147,31,147,30,54,31,80,31,57,31,170,31,170,30,235,31,186,31,75,31,200,31,201,31,59,31,208,31,22,31,214,31,139,31,116,31,108,31,41,31,176,31,176,30,85,31,101,31,77,31,177,31,177,30,175,31,8,31,247,31,247,30,114,31,35,31,142,31,142,30,210,31,194,31,176,31,158,31,158,30,141,31,14,31,129,31,205,31,45,31,110,31,110,30,69,31,55,31,54,31,25,31,138,31,118,31,94,31,105,31,232,31,232,30,232,29,232,28,89,31,134,31,154,31,154,30,202,31,252,31,123,31,176,31,5,31,5,30,224,31,194,31,174,31,203,31,168,31,151,31,247,31,83,31,181,31,211,31,105,31,105,30,85,31,126,31,200,31,94,31,28,31,238,31,9,31,131,31,219,31,28,31,28,30,32,31,107,31,107,30,3,31,115,31,144,31,20,31,65,31,6,31,168,31,224,31,47,31,39,31,39,30,61,31,14,31,195,31,102,31,102,30,124,31,238,31,238,30,7,31,89,31,89,30,176,31,63,31,184,31,184,30,223,31,250,31,235,31,235,30,46,31,81,31,11,31,173,31,254,31,204,31,204,30,53,31,124,31,156,31,156,30,4,31,4,30,4,29,4,28,211,31,35,31,18,31,156,31,129,31,114,31,112,31,195,31,3,31,35,31,204,31,204,30,222,31,139,31,137,31,102,31,144,31,211,31,246,31,183,31,7,31,216,31,216,30,216,29,93,31,242,31,173,31,172,31,172,30,53,31,156,31,85,31,62,31,62,30,46,31,186,31,158,31,158,30,201,31,48,31,165,31,114,31,114,30,112,31,105,31,15,31,164,31,207,31,105,31,100,31,100,30,85,31,208,31,208,30,92,31,52,31,51,31,51,30,115,31,57,31,183,31,223,31,172,31,167,31,163,31,12,31,126,31,40,31,229,31,203,31,185,31,66,31,213,31,214,31,88,31,25,31,255,31,8,31,8,30,132,31,172,31,172,30,115,31,115,30,219,31,219,30,234,31,73,31,188,31,6,31,8,31,242,31,53,31,253,31,181,31,108,31,71,31,80,31,211,31,6,31,187,31,165,31,176,31,176,30,176,29,58,31,58,30,103,31,243,31,171,31,99,31,167,31,251,31,100,31,13,31,140,31,38,31,115,31,61,31,104,31,247,31,120,31,205,31,134,31,48,31,10,31,104,31,104,30,60,31,238,31,119,31,131,31,131,30,134,31,223,31,223,30,223,29,67,31,137,31,96,31,231,31,231,30,139,31,139,30,212,31,2,31,166,31,110,31,43,31,123,31,13,31,13,30,28,31,129,31,67,31,67,30,183,31,30,31,120,31,17,31,17,30,89,31,139,31,231,31,50,31,88,31,204,31,204,30,100,31,11,31,93,31,176,31,180,31,253,31,176,31,223,31,232,31,233,31,228,31,83,31,36,31,36,30,45,31,45,30,204,31,204,30,69,31,73,31,169,31,210,31,210,30,37,31,193,31,215,31,179,31,179,30,179,29,161,31,156,31,156,30,16,31,136,31,169,31,224,31,18,31,18,30,255,31,130,31,130,30,225,31,225,30,225,29,112,31,151,31,151,30,53,31,75,31,80,31,108,31,48,31,48,30,44,31,118,31,118,30,200,31,79,31,251,31,145,31,145,30,231,31,139,31,250,31,51,31,51,30,137,31,187,31,187,30,187,29,183,31,127,31,230,31,230,30,107,31,18,31,22,31,22,30,143,31,37,31,37,30,178,31,62,31,228,31,9,31,112,31,26,31,234,31,187,31,109,31,57,31,57,30,124,31,226,31,248,31,153,31,13,31,13,30,37,31,249,31,249,30,249,29,249,28,249,27,249,26,249,25,165,31,192,31,143,31,40,31,40,30,223,31,93,31,93,30,255,31,176,31,176,30,21,31,136,31,97,31,13,31,94,31,94,30,165,31,165,30,100,31,212,31,254,31,18,31,18,30,157,31,25,31,58,31,116,31,116,30,48,31,28,31,28,30,119,31,119,30,6,31,226,31,226,30,103,31,100,31,211,31,145,31,90,31,90,30,90,29,90,28,64,31,1,31,235,31,1,31,243,31,69,31,69,30,69,29,167,31,167,30,67,31,11,31,168,31,168,30,173,31,231,31,86,31,132,31,132,30,132,29,192,31,192,30,192,29,227,31,44,31,44,30,169,31,254,31,32,31,61,31,166,31,37,31,37,30,37,29,37,28,220,31,220,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
