-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_700 is
end project_tb_700;

architecture project_tb_arch_700 of project_tb_700 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 829;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (168,0,181,0,82,0,151,0,177,0,114,0,0,0,97,0,50,0,18,0,110,0,14,0,84,0,0,0,55,0,189,0,0,0,185,0,66,0,95,0,80,0,222,0,203,0,33,0,118,0,0,0,0,0,62,0,159,0,102,0,28,0,93,0,195,0,43,0,224,0,61,0,220,0,8,0,90,0,19,0,42,0,135,0,208,0,0,0,210,0,34,0,205,0,101,0,196,0,86,0,68,0,161,0,223,0,18,0,0,0,148,0,0,0,167,0,255,0,72,0,213,0,0,0,26,0,0,0,0,0,182,0,173,0,127,0,146,0,84,0,118,0,104,0,82,0,78,0,156,0,181,0,59,0,250,0,154,0,242,0,242,0,88,0,203,0,70,0,15,0,154,0,206,0,72,0,24,0,68,0,131,0,15,0,0,0,192,0,111,0,147,0,232,0,12,0,27,0,121,0,127,0,39,0,0,0,58,0,154,0,166,0,26,0,215,0,0,0,33,0,73,0,159,0,88,0,51,0,0,0,92,0,123,0,185,0,200,0,107,0,183,0,33,0,53,0,194,0,3,0,0,0,9,0,0,0,219,0,203,0,17,0,227,0,69,0,197,0,0,0,196,0,105,0,59,0,0,0,64,0,150,0,0,0,0,0,54,0,178,0,106,0,219,0,0,0,0,0,0,0,22,0,29,0,8,0,0,0,254,0,210,0,214,0,67,0,32,0,96,0,0,0,65,0,73,0,0,0,233,0,0,0,28,0,152,0,137,0,246,0,0,0,0,0,193,0,245,0,241,0,234,0,0,0,19,0,0,0,198,0,24,0,0,0,0,0,157,0,0,0,77,0,200,0,119,0,0,0,76,0,55,0,181,0,41,0,131,0,22,0,125,0,0,0,63,0,172,0,165,0,132,0,0,0,149,0,149,0,79,0,93,0,72,0,183,0,0,0,231,0,33,0,0,0,0,0,31,0,207,0,25,0,142,0,28,0,118,0,168,0,175,0,61,0,55,0,230,0,209,0,98,0,0,0,222,0,66,0,213,0,43,0,196,0,132,0,255,0,135,0,0,0,11,0,0,0,194,0,130,0,197,0,29,0,0,0,0,0,248,0,167,0,104,0,15,0,132,0,246,0,0,0,167,0,91,0,113,0,127,0,184,0,228,0,216,0,21,0,34,0,245,0,0,0,33,0,118,0,192,0,89,0,0,0,236,0,0,0,81,0,0,0,6,0,242,0,55,0,109,0,246,0,0,0,137,0,68,0,25,0,151,0,178,0,131,0,0,0,174,0,155,0,0,0,206,0,28,0,85,0,0,0,43,0,0,0,0,0,132,0,0,0,48,0,248,0,241,0,113,0,146,0,0,0,143,0,93,0,0,0,0,0,0,0,194,0,87,0,86,0,51,0,33,0,95,0,136,0,157,0,0,0,181,0,89,0,212,0,50,0,156,0,117,0,111,0,45,0,0,0,88,0,202,0,40,0,191,0,148,0,79,0,44,0,0,0,0,0,132,0,62,0,144,0,41,0,0,0,124,0,236,0,0,0,174,0,94,0,191,0,255,0,0,0,0,0,81,0,111,0,99,0,136,0,0,0,0,0,235,0,35,0,72,0,140,0,32,0,0,0,183,0,223,0,0,0,118,0,153,0,0,0,0,0,142,0,20,0,0,0,119,0,48,0,101,0,0,0,149,0,27,0,52,0,250,0,201,0,253,0,123,0,211,0,17,0,68,0,180,0,2,0,0,0,20,0,76,0,80,0,117,0,130,0,174,0,90,0,0,0,0,0,137,0,89,0,99,0,52,0,27,0,0,0,19,0,56,0,196,0,207,0,86,0,81,0,181,0,236,0,79,0,0,0,0,0,0,0,0,0,67,0,177,0,4,0,0,0,148,0,89,0,20,0,156,0,22,0,22,0,0,0,0,0,108,0,20,0,0,0,251,0,228,0,207,0,2,0,0,0,0,0,164,0,191,0,239,0,189,0,31,0,21,0,40,0,35,0,101,0,0,0,4,0,0,0,41,0,96,0,120,0,141,0,230,0,11,0,0,0,0,0,0,0,249,0,156,0,72,0,216,0,213,0,0,0,103,0,70,0,130,0,124,0,0,0,195,0,161,0,153,0,0,0,93,0,74,0,182,0,206,0,110,0,27,0,183,0,103,0,127,0,65,0,171,0,96,0,152,0,157,0,27,0,187,0,152,0,225,0,248,0,0,0,97,0,0,0,9,0,0,0,109,0,233,0,74,0,174,0,0,0,66,0,0,0,217,0,59,0,5,0,249,0,184,0,239,0,0,0,234,0,122,0,66,0,13,0,28,0,15,0,251,0,0,0,12,0,13,0,0,0,5,0,39,0,39,0,195,0,78,0,255,0,153,0,37,0,0,0,37,0,144,0,157,0,98,0,122,0,149,0,0,0,161,0,49,0,84,0,0,0,210,0,80,0,183,0,112,0,0,0,147,0,99,0,16,0,109,0,0,0,241,0,60,0,246,0,36,0,239,0,0,0,186,0,53,0,0,0,0,0,181,0,181,0,9,0,42,0,238,0,0,0,0,0,45,0,67,0,0,0,125,0,42,0,33,0,25,0,123,0,62,0,248,0,64,0,246,0,33,0,0,0,200,0,0,0,67,0,106,0,70,0,195,0,176,0,214,0,191,0,0,0,0,0,112,0,229,0,2,0,106,0,169,0,149,0,231,0,80,0,43,0,46,0,143,0,240,0,144,0,216,0,104,0,160,0,0,0,91,0,0,0,115,0,0,0,0,0,245,0,0,0,208,0,177,0,38,0,69,0,0,0,150,0,252,0,175,0,99,0,0,0,74,0,203,0,185,0,0,0,10,0,148,0,185,0,183,0,0,0,135,0,137,0,180,0,184,0,149,0,195,0,218,0,68,0,173,0,29,0,57,0,68,0,211,0,175,0,0,0,198,0,125,0,203,0,17,0,217,0,219,0,225,0,0,0,171,0,249,0,0,0,175,0,8,0,237,0,200,0,64,0,137,0,82,0,0,0,60,0,0,0,255,0,119,0,71,0,184,0,0,0,167,0,144,0,53,0,0,0,0,0,111,0,0,0,145,0,184,0,251,0,60,0,239,0,0,0,180,0,228,0,82,0,49,0,148,0,98,0,0,0,156,0,246,0,73,0,6,0,238,0,248,0,113,0,120,0,0,0,75,0,181,0,108,0,155,0,0,0,115,0,52,0,161,0,18,0,0,0,134,0,134,0,120,0,8,0,127,0,46,0,72,0,12,0,0,0,124,0,224,0,69,0,186,0,0,0,94,0,0,0,254,0,0,0,41,0,32,0,157,0,16,0,116,0,164,0,70,0,17,0,8,0,196,0,38,0,224,0,76,0,33,0,78,0,198,0,242,0,20,0,56,0,31,0,98,0,166,0,139,0,0,0,202,0,0,0,7,0,223,0,115,0,245,0,54,0,114,0,254,0,27,0,162,0,37,0,47,0,0,0,119,0,137,0,221,0,1,0,68,0,199,0,97,0,176,0,215,0,0,0,0,0,0,0,0,0,105,0,36,0,150,0,113,0,0,0,0,0,37,0,39,0,90,0,120,0,226,0,35,0,137,0,211,0,104,0,53,0,0,0,189,0,69,0,223,0,157,0,19,0,239,0,221,0,245,0,248,0,161,0,0,0,253,0,132,0,74,0,77,0,119,0,29,0,48,0,198,0,178,0,11,0,224,0,199,0,124,0,56,0,225,0,0,0);
signal scenario_full  : scenario_type := (168,31,181,31,82,31,151,31,177,31,114,31,114,30,97,31,50,31,18,31,110,31,14,31,84,31,84,30,55,31,189,31,189,30,185,31,66,31,95,31,80,31,222,31,203,31,33,31,118,31,118,30,118,29,62,31,159,31,102,31,28,31,93,31,195,31,43,31,224,31,61,31,220,31,8,31,90,31,19,31,42,31,135,31,208,31,208,30,210,31,34,31,205,31,101,31,196,31,86,31,68,31,161,31,223,31,18,31,18,30,148,31,148,30,167,31,255,31,72,31,213,31,213,30,26,31,26,30,26,29,182,31,173,31,127,31,146,31,84,31,118,31,104,31,82,31,78,31,156,31,181,31,59,31,250,31,154,31,242,31,242,31,88,31,203,31,70,31,15,31,154,31,206,31,72,31,24,31,68,31,131,31,15,31,15,30,192,31,111,31,147,31,232,31,12,31,27,31,121,31,127,31,39,31,39,30,58,31,154,31,166,31,26,31,215,31,215,30,33,31,73,31,159,31,88,31,51,31,51,30,92,31,123,31,185,31,200,31,107,31,183,31,33,31,53,31,194,31,3,31,3,30,9,31,9,30,219,31,203,31,17,31,227,31,69,31,197,31,197,30,196,31,105,31,59,31,59,30,64,31,150,31,150,30,150,29,54,31,178,31,106,31,219,31,219,30,219,29,219,28,22,31,29,31,8,31,8,30,254,31,210,31,214,31,67,31,32,31,96,31,96,30,65,31,73,31,73,30,233,31,233,30,28,31,152,31,137,31,246,31,246,30,246,29,193,31,245,31,241,31,234,31,234,30,19,31,19,30,198,31,24,31,24,30,24,29,157,31,157,30,77,31,200,31,119,31,119,30,76,31,55,31,181,31,41,31,131,31,22,31,125,31,125,30,63,31,172,31,165,31,132,31,132,30,149,31,149,31,79,31,93,31,72,31,183,31,183,30,231,31,33,31,33,30,33,29,31,31,207,31,25,31,142,31,28,31,118,31,168,31,175,31,61,31,55,31,230,31,209,31,98,31,98,30,222,31,66,31,213,31,43,31,196,31,132,31,255,31,135,31,135,30,11,31,11,30,194,31,130,31,197,31,29,31,29,30,29,29,248,31,167,31,104,31,15,31,132,31,246,31,246,30,167,31,91,31,113,31,127,31,184,31,228,31,216,31,21,31,34,31,245,31,245,30,33,31,118,31,192,31,89,31,89,30,236,31,236,30,81,31,81,30,6,31,242,31,55,31,109,31,246,31,246,30,137,31,68,31,25,31,151,31,178,31,131,31,131,30,174,31,155,31,155,30,206,31,28,31,85,31,85,30,43,31,43,30,43,29,132,31,132,30,48,31,248,31,241,31,113,31,146,31,146,30,143,31,93,31,93,30,93,29,93,28,194,31,87,31,86,31,51,31,33,31,95,31,136,31,157,31,157,30,181,31,89,31,212,31,50,31,156,31,117,31,111,31,45,31,45,30,88,31,202,31,40,31,191,31,148,31,79,31,44,31,44,30,44,29,132,31,62,31,144,31,41,31,41,30,124,31,236,31,236,30,174,31,94,31,191,31,255,31,255,30,255,29,81,31,111,31,99,31,136,31,136,30,136,29,235,31,35,31,72,31,140,31,32,31,32,30,183,31,223,31,223,30,118,31,153,31,153,30,153,29,142,31,20,31,20,30,119,31,48,31,101,31,101,30,149,31,27,31,52,31,250,31,201,31,253,31,123,31,211,31,17,31,68,31,180,31,2,31,2,30,20,31,76,31,80,31,117,31,130,31,174,31,90,31,90,30,90,29,137,31,89,31,99,31,52,31,27,31,27,30,19,31,56,31,196,31,207,31,86,31,81,31,181,31,236,31,79,31,79,30,79,29,79,28,79,27,67,31,177,31,4,31,4,30,148,31,89,31,20,31,156,31,22,31,22,31,22,30,22,29,108,31,20,31,20,30,251,31,228,31,207,31,2,31,2,30,2,29,164,31,191,31,239,31,189,31,31,31,21,31,40,31,35,31,101,31,101,30,4,31,4,30,41,31,96,31,120,31,141,31,230,31,11,31,11,30,11,29,11,28,249,31,156,31,72,31,216,31,213,31,213,30,103,31,70,31,130,31,124,31,124,30,195,31,161,31,153,31,153,30,93,31,74,31,182,31,206,31,110,31,27,31,183,31,103,31,127,31,65,31,171,31,96,31,152,31,157,31,27,31,187,31,152,31,225,31,248,31,248,30,97,31,97,30,9,31,9,30,109,31,233,31,74,31,174,31,174,30,66,31,66,30,217,31,59,31,5,31,249,31,184,31,239,31,239,30,234,31,122,31,66,31,13,31,28,31,15,31,251,31,251,30,12,31,13,31,13,30,5,31,39,31,39,31,195,31,78,31,255,31,153,31,37,31,37,30,37,31,144,31,157,31,98,31,122,31,149,31,149,30,161,31,49,31,84,31,84,30,210,31,80,31,183,31,112,31,112,30,147,31,99,31,16,31,109,31,109,30,241,31,60,31,246,31,36,31,239,31,239,30,186,31,53,31,53,30,53,29,181,31,181,31,9,31,42,31,238,31,238,30,238,29,45,31,67,31,67,30,125,31,42,31,33,31,25,31,123,31,62,31,248,31,64,31,246,31,33,31,33,30,200,31,200,30,67,31,106,31,70,31,195,31,176,31,214,31,191,31,191,30,191,29,112,31,229,31,2,31,106,31,169,31,149,31,231,31,80,31,43,31,46,31,143,31,240,31,144,31,216,31,104,31,160,31,160,30,91,31,91,30,115,31,115,30,115,29,245,31,245,30,208,31,177,31,38,31,69,31,69,30,150,31,252,31,175,31,99,31,99,30,74,31,203,31,185,31,185,30,10,31,148,31,185,31,183,31,183,30,135,31,137,31,180,31,184,31,149,31,195,31,218,31,68,31,173,31,29,31,57,31,68,31,211,31,175,31,175,30,198,31,125,31,203,31,17,31,217,31,219,31,225,31,225,30,171,31,249,31,249,30,175,31,8,31,237,31,200,31,64,31,137,31,82,31,82,30,60,31,60,30,255,31,119,31,71,31,184,31,184,30,167,31,144,31,53,31,53,30,53,29,111,31,111,30,145,31,184,31,251,31,60,31,239,31,239,30,180,31,228,31,82,31,49,31,148,31,98,31,98,30,156,31,246,31,73,31,6,31,238,31,248,31,113,31,120,31,120,30,75,31,181,31,108,31,155,31,155,30,115,31,52,31,161,31,18,31,18,30,134,31,134,31,120,31,8,31,127,31,46,31,72,31,12,31,12,30,124,31,224,31,69,31,186,31,186,30,94,31,94,30,254,31,254,30,41,31,32,31,157,31,16,31,116,31,164,31,70,31,17,31,8,31,196,31,38,31,224,31,76,31,33,31,78,31,198,31,242,31,20,31,56,31,31,31,98,31,166,31,139,31,139,30,202,31,202,30,7,31,223,31,115,31,245,31,54,31,114,31,254,31,27,31,162,31,37,31,47,31,47,30,119,31,137,31,221,31,1,31,68,31,199,31,97,31,176,31,215,31,215,30,215,29,215,28,215,27,105,31,36,31,150,31,113,31,113,30,113,29,37,31,39,31,90,31,120,31,226,31,35,31,137,31,211,31,104,31,53,31,53,30,189,31,69,31,223,31,157,31,19,31,239,31,221,31,245,31,248,31,161,31,161,30,253,31,132,31,74,31,77,31,119,31,29,31,48,31,198,31,178,31,11,31,224,31,199,31,124,31,56,31,225,31,225,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
