-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_396 is
end project_tb_396;

architecture project_tb_arch_396 of project_tb_396 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 707;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (208,0,117,0,226,0,166,0,123,0,0,0,131,0,79,0,83,0,235,0,221,0,69,0,131,0,0,0,0,0,0,0,190,0,106,0,0,0,9,0,33,0,102,0,225,0,124,0,0,0,172,0,217,0,212,0,155,0,43,0,22,0,138,0,67,0,94,0,18,0,76,0,247,0,0,0,0,0,228,0,129,0,0,0,78,0,0,0,0,0,55,0,217,0,38,0,88,0,0,0,69,0,25,0,153,0,144,0,103,0,254,0,191,0,0,0,251,0,219,0,0,0,0,0,109,0,0,0,6,0,63,0,8,0,6,0,61,0,186,0,147,0,5,0,190,0,95,0,245,0,200,0,118,0,170,0,9,0,182,0,98,0,177,0,156,0,191,0,239,0,56,0,110,0,0,0,26,0,162,0,46,0,113,0,126,0,71,0,57,0,142,0,8,0,229,0,111,0,215,0,0,0,154,0,66,0,220,0,0,0,238,0,219,0,120,0,171,0,64,0,122,0,212,0,26,0,107,0,0,0,222,0,141,0,242,0,85,0,75,0,223,0,5,0,190,0,127,0,0,0,52,0,85,0,14,0,104,0,214,0,0,0,140,0,86,0,73,0,164,0,92,0,233,0,201,0,174,0,0,0,90,0,0,0,0,0,2,0,88,0,248,0,92,0,128,0,0,0,178,0,65,0,43,0,0,0,254,0,162,0,95,0,44,0,0,0,236,0,127,0,246,0,0,0,79,0,42,0,82,0,236,0,230,0,217,0,79,0,0,0,220,0,0,0,75,0,138,0,0,0,206,0,0,0,0,0,0,0,157,0,0,0,176,0,133,0,0,0,0,0,78,0,76,0,0,0,125,0,41,0,157,0,109,0,130,0,231,0,146,0,0,0,195,0,0,0,54,0,88,0,0,0,87,0,170,0,159,0,0,0,242,0,9,0,0,0,212,0,8,0,0,0,40,0,105,0,54,0,169,0,152,0,0,0,11,0,0,0,98,0,134,0,51,0,238,0,105,0,0,0,148,0,131,0,124,0,0,0,243,0,157,0,177,0,126,0,0,0,76,0,17,0,36,0,168,0,144,0,86,0,19,0,0,0,178,0,170,0,35,0,0,0,100,0,83,0,237,0,106,0,229,0,44,0,0,0,0,0,125,0,166,0,212,0,58,0,140,0,116,0,43,0,0,0,177,0,181,0,0,0,0,0,222,0,218,0,220,0,139,0,0,0,107,0,253,0,224,0,99,0,41,0,41,0,90,0,224,0,64,0,22,0,125,0,0,0,57,0,179,0,108,0,74,0,51,0,0,0,0,0,220,0,0,0,0,0,142,0,169,0,3,0,64,0,124,0,131,0,0,0,9,0,208,0,193,0,0,0,0,0,185,0,0,0,114,0,9,0,3,0,233,0,76,0,185,0,195,0,0,0,6,0,234,0,136,0,72,0,13,0,120,0,237,0,17,0,1,0,123,0,0,0,0,0,16,0,0,0,47,0,117,0,231,0,114,0,55,0,198,0,237,0,0,0,64,0,239,0,0,0,0,0,9,0,123,0,30,0,112,0,0,0,0,0,240,0,106,0,107,0,219,0,78,0,131,0,0,0,247,0,113,0,111,0,236,0,70,0,24,0,0,0,0,0,40,0,18,0,213,0,204,0,178,0,213,0,4,0,46,0,199,0,160,0,0,0,35,0,137,0,204,0,89,0,7,0,0,0,46,0,4,0,0,0,126,0,83,0,0,0,0,0,98,0,0,0,0,0,45,0,126,0,183,0,0,0,96,0,47,0,136,0,35,0,35,0,103,0,106,0,204,0,0,0,171,0,206,0,7,0,0,0,140,0,228,0,182,0,0,0,111,0,0,0,117,0,164,0,93,0,92,0,0,0,0,0,0,0,40,0,122,0,129,0,0,0,49,0,124,0,22,0,165,0,138,0,188,0,233,0,100,0,133,0,20,0,91,0,217,0,15,0,39,0,217,0,194,0,147,0,92,0,203,0,169,0,227,0,98,0,24,0,31,0,80,0,92,0,93,0,76,0,48,0,128,0,106,0,91,0,0,0,146,0,192,0,69,0,141,0,0,0,0,0,180,0,0,0,50,0,236,0,107,0,4,0,188,0,22,0,0,0,126,0,0,0,100,0,144,0,49,0,192,0,43,0,130,0,178,0,237,0,140,0,233,0,76,0,0,0,205,0,182,0,0,0,164,0,0,0,221,0,136,0,70,0,232,0,255,0,105,0,238,0,0,0,0,0,122,0,2,0,25,0,144,0,134,0,17,0,205,0,146,0,0,0,190,0,234,0,0,0,146,0,0,0,39,0,0,0,14,0,232,0,64,0,132,0,0,0,144,0,173,0,0,0,181,0,223,0,23,0,93,0,105,0,145,0,11,0,0,0,176,0,228,0,0,0,125,0,48,0,0,0,214,0,38,0,236,0,232,0,113,0,63,0,108,0,208,0,0,0,117,0,80,0,128,0,0,0,139,0,200,0,78,0,49,0,173,0,194,0,199,0,0,0,51,0,230,0,238,0,227,0,169,0,207,0,0,0,181,0,117,0,214,0,81,0,40,0,234,0,208,0,101,0,244,0,192,0,17,0,183,0,253,0,221,0,121,0,244,0,156,0,61,0,68,0,58,0,91,0,0,0,6,0,115,0,0,0,203,0,0,0,43,0,216,0,37,0,179,0,6,0,0,0,95,0,0,0,0,0,57,0,119,0,0,0,0,0,112,0,0,0,34,0,179,0,42,0,81,0,81,0,0,0,0,0,0,0,0,0,0,0,0,0,82,0,91,0,136,0,90,0,10,0,236,0,37,0,16,0,150,0,78,0,88,0,121,0,238,0,225,0,93,0,0,0,222,0,90,0,23,0,101,0,0,0,25,0,8,0,147,0,0,0,101,0,167,0,96,0,206,0,179,0,183,0,52,0,110,0,0,0,73,0,179,0,86,0,0,0,198,0,207,0,42,0,0,0,0,0,227,0,13,0,229,0,64,0,0,0,0,0,220,0,5,0,2,0,12,0,0,0,151,0,0,0,102,0,0,0,87,0,195,0,238,0,0,0,238,0,13,0,0,0,153,0,130,0,218,0,5,0,0,0,145,0,149,0,0,0,0,0,155,0,148,0,35,0,240,0,0,0,35,0,143,0,19,0,191,0,105,0,91,0,79,0,104,0,0,0,187,0);
signal scenario_full  : scenario_type := (208,31,117,31,226,31,166,31,123,31,123,30,131,31,79,31,83,31,235,31,221,31,69,31,131,31,131,30,131,29,131,28,190,31,106,31,106,30,9,31,33,31,102,31,225,31,124,31,124,30,172,31,217,31,212,31,155,31,43,31,22,31,138,31,67,31,94,31,18,31,76,31,247,31,247,30,247,29,228,31,129,31,129,30,78,31,78,30,78,29,55,31,217,31,38,31,88,31,88,30,69,31,25,31,153,31,144,31,103,31,254,31,191,31,191,30,251,31,219,31,219,30,219,29,109,31,109,30,6,31,63,31,8,31,6,31,61,31,186,31,147,31,5,31,190,31,95,31,245,31,200,31,118,31,170,31,9,31,182,31,98,31,177,31,156,31,191,31,239,31,56,31,110,31,110,30,26,31,162,31,46,31,113,31,126,31,71,31,57,31,142,31,8,31,229,31,111,31,215,31,215,30,154,31,66,31,220,31,220,30,238,31,219,31,120,31,171,31,64,31,122,31,212,31,26,31,107,31,107,30,222,31,141,31,242,31,85,31,75,31,223,31,5,31,190,31,127,31,127,30,52,31,85,31,14,31,104,31,214,31,214,30,140,31,86,31,73,31,164,31,92,31,233,31,201,31,174,31,174,30,90,31,90,30,90,29,2,31,88,31,248,31,92,31,128,31,128,30,178,31,65,31,43,31,43,30,254,31,162,31,95,31,44,31,44,30,236,31,127,31,246,31,246,30,79,31,42,31,82,31,236,31,230,31,217,31,79,31,79,30,220,31,220,30,75,31,138,31,138,30,206,31,206,30,206,29,206,28,157,31,157,30,176,31,133,31,133,30,133,29,78,31,76,31,76,30,125,31,41,31,157,31,109,31,130,31,231,31,146,31,146,30,195,31,195,30,54,31,88,31,88,30,87,31,170,31,159,31,159,30,242,31,9,31,9,30,212,31,8,31,8,30,40,31,105,31,54,31,169,31,152,31,152,30,11,31,11,30,98,31,134,31,51,31,238,31,105,31,105,30,148,31,131,31,124,31,124,30,243,31,157,31,177,31,126,31,126,30,76,31,17,31,36,31,168,31,144,31,86,31,19,31,19,30,178,31,170,31,35,31,35,30,100,31,83,31,237,31,106,31,229,31,44,31,44,30,44,29,125,31,166,31,212,31,58,31,140,31,116,31,43,31,43,30,177,31,181,31,181,30,181,29,222,31,218,31,220,31,139,31,139,30,107,31,253,31,224,31,99,31,41,31,41,31,90,31,224,31,64,31,22,31,125,31,125,30,57,31,179,31,108,31,74,31,51,31,51,30,51,29,220,31,220,30,220,29,142,31,169,31,3,31,64,31,124,31,131,31,131,30,9,31,208,31,193,31,193,30,193,29,185,31,185,30,114,31,9,31,3,31,233,31,76,31,185,31,195,31,195,30,6,31,234,31,136,31,72,31,13,31,120,31,237,31,17,31,1,31,123,31,123,30,123,29,16,31,16,30,47,31,117,31,231,31,114,31,55,31,198,31,237,31,237,30,64,31,239,31,239,30,239,29,9,31,123,31,30,31,112,31,112,30,112,29,240,31,106,31,107,31,219,31,78,31,131,31,131,30,247,31,113,31,111,31,236,31,70,31,24,31,24,30,24,29,40,31,18,31,213,31,204,31,178,31,213,31,4,31,46,31,199,31,160,31,160,30,35,31,137,31,204,31,89,31,7,31,7,30,46,31,4,31,4,30,126,31,83,31,83,30,83,29,98,31,98,30,98,29,45,31,126,31,183,31,183,30,96,31,47,31,136,31,35,31,35,31,103,31,106,31,204,31,204,30,171,31,206,31,7,31,7,30,140,31,228,31,182,31,182,30,111,31,111,30,117,31,164,31,93,31,92,31,92,30,92,29,92,28,40,31,122,31,129,31,129,30,49,31,124,31,22,31,165,31,138,31,188,31,233,31,100,31,133,31,20,31,91,31,217,31,15,31,39,31,217,31,194,31,147,31,92,31,203,31,169,31,227,31,98,31,24,31,31,31,80,31,92,31,93,31,76,31,48,31,128,31,106,31,91,31,91,30,146,31,192,31,69,31,141,31,141,30,141,29,180,31,180,30,50,31,236,31,107,31,4,31,188,31,22,31,22,30,126,31,126,30,100,31,144,31,49,31,192,31,43,31,130,31,178,31,237,31,140,31,233,31,76,31,76,30,205,31,182,31,182,30,164,31,164,30,221,31,136,31,70,31,232,31,255,31,105,31,238,31,238,30,238,29,122,31,2,31,25,31,144,31,134,31,17,31,205,31,146,31,146,30,190,31,234,31,234,30,146,31,146,30,39,31,39,30,14,31,232,31,64,31,132,31,132,30,144,31,173,31,173,30,181,31,223,31,23,31,93,31,105,31,145,31,11,31,11,30,176,31,228,31,228,30,125,31,48,31,48,30,214,31,38,31,236,31,232,31,113,31,63,31,108,31,208,31,208,30,117,31,80,31,128,31,128,30,139,31,200,31,78,31,49,31,173,31,194,31,199,31,199,30,51,31,230,31,238,31,227,31,169,31,207,31,207,30,181,31,117,31,214,31,81,31,40,31,234,31,208,31,101,31,244,31,192,31,17,31,183,31,253,31,221,31,121,31,244,31,156,31,61,31,68,31,58,31,91,31,91,30,6,31,115,31,115,30,203,31,203,30,43,31,216,31,37,31,179,31,6,31,6,30,95,31,95,30,95,29,57,31,119,31,119,30,119,29,112,31,112,30,34,31,179,31,42,31,81,31,81,31,81,30,81,29,81,28,81,27,81,26,81,25,82,31,91,31,136,31,90,31,10,31,236,31,37,31,16,31,150,31,78,31,88,31,121,31,238,31,225,31,93,31,93,30,222,31,90,31,23,31,101,31,101,30,25,31,8,31,147,31,147,30,101,31,167,31,96,31,206,31,179,31,183,31,52,31,110,31,110,30,73,31,179,31,86,31,86,30,198,31,207,31,42,31,42,30,42,29,227,31,13,31,229,31,64,31,64,30,64,29,220,31,5,31,2,31,12,31,12,30,151,31,151,30,102,31,102,30,87,31,195,31,238,31,238,30,238,31,13,31,13,30,153,31,130,31,218,31,5,31,5,30,145,31,149,31,149,30,149,29,155,31,148,31,35,31,240,31,240,30,35,31,143,31,19,31,191,31,105,31,91,31,79,31,104,31,104,30,187,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
