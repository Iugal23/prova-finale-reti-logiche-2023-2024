-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 406;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,98,0,194,0,44,0,112,0,96,0,170,0,164,0,64,0,195,0,0,0,26,0,138,0,95,0,85,0,72,0,249,0,223,0,38,0,1,0,154,0,216,0,0,0,213,0,16,0,223,0,191,0,8,0,162,0,0,0,195,0,153,0,209,0,60,0,0,0,115,0,104,0,206,0,82,0,8,0,14,0,214,0,215,0,0,0,75,0,88,0,0,0,170,0,233,0,104,0,84,0,0,0,170,0,139,0,0,0,45,0,75,0,110,0,135,0,231,0,247,0,0,0,51,0,0,0,42,0,218,0,0,0,0,0,172,0,206,0,104,0,143,0,67,0,0,0,7,0,24,0,175,0,127,0,243,0,38,0,0,0,0,0,160,0,14,0,70,0,0,0,41,0,185,0,172,0,0,0,117,0,0,0,51,0,0,0,207,0,91,0,0,0,139,0,6,0,0,0,0,0,82,0,254,0,0,0,143,0,182,0,206,0,21,0,5,0,72,0,92,0,211,0,182,0,178,0,116,0,221,0,83,0,174,0,219,0,0,0,247,0,120,0,49,0,224,0,145,0,0,0,202,0,243,0,238,0,215,0,0,0,0,0,0,0,0,0,0,0,192,0,22,0,0,0,94,0,0,0,144,0,209,0,51,0,101,0,0,0,254,0,125,0,138,0,164,0,141,0,253,0,180,0,210,0,48,0,62,0,0,0,221,0,0,0,91,0,225,0,0,0,75,0,12,0,221,0,120,0,84,0,94,0,163,0,18,0,120,0,67,0,0,0,167,0,164,0,71,0,171,0,0,0,0,0,108,0,18,0,74,0,109,0,61,0,28,0,170,0,119,0,10,0,254,0,224,0,196,0,47,0,0,0,247,0,61,0,0,0,68,0,8,0,108,0,0,0,192,0,141,0,0,0,173,0,97,0,3,0,99,0,0,0,0,0,179,0,143,0,3,0,62,0,46,0,0,0,103,0,192,0,217,0,38,0,36,0,37,0,152,0,9,0,0,0,44,0,11,0,100,0,180,0,30,0,139,0,36,0,62,0,0,0,0,0,198,0,50,0,0,0,0,0,37,0,210,0,0,0,44,0,107,0,205,0,0,0,3,0,102,0,2,0,21,0,142,0,186,0,109,0,116,0,224,0,125,0,252,0,31,0,98,0,233,0,14,0,0,0,24,0,7,0,157,0,46,0,0,0,42,0,102,0,0,0,213,0,197,0,0,0,100,0,192,0,210,0,184,0,80,0,179,0,0,0,1,0,59,0,196,0,231,0,244,0,50,0,11,0,0,0,176,0,8,0,0,0,33,0,170,0,0,0,0,0,163,0,60,0,0,0,156,0,225,0,120,0,163,0,188,0,50,0,148,0,0,0,252,0,178,0,0,0,97,0,0,0,0,0,83,0,198,0,91,0,193,0,180,0,122,0,139,0,220,0,123,0,9,0,15,0,35,0,213,0,216,0,247,0,102,0,225,0,92,0,246,0,0,0,226,0,0,0,220,0,50,0,140,0,86,0,82,0,115,0,98,0,124,0,13,0,186,0,165,0,73,0,45,0,153,0,0,0,235,0,150,0,117,0,140,0,133,0,0,0,0,0,92,0,0,0,241,0,71,0,123,0,0,0,230,0,249,0,82,0,147,0,97,0,132,0,60,0,94,0,4,0,213,0,32,0,5,0,0,0,104,0,124,0,230,0,77,0,162,0,0,0,44,0,213,0,0,0,198,0,47,0,124,0,184,0,152,0,58,0,0,0,0,0,169,0,219,0,126,0,32,0,0,0,119,0,0,0,0,0,40,0,200,0,31,0,226,0,0,0,189,0,26,0,213,0);
signal scenario_full  : scenario_type := (0,0,98,31,194,31,44,31,112,31,96,31,170,31,164,31,64,31,195,31,195,30,26,31,138,31,95,31,85,31,72,31,249,31,223,31,38,31,1,31,154,31,216,31,216,30,213,31,16,31,223,31,191,31,8,31,162,31,162,30,195,31,153,31,209,31,60,31,60,30,115,31,104,31,206,31,82,31,8,31,14,31,214,31,215,31,215,30,75,31,88,31,88,30,170,31,233,31,104,31,84,31,84,30,170,31,139,31,139,30,45,31,75,31,110,31,135,31,231,31,247,31,247,30,51,31,51,30,42,31,218,31,218,30,218,29,172,31,206,31,104,31,143,31,67,31,67,30,7,31,24,31,175,31,127,31,243,31,38,31,38,30,38,29,160,31,14,31,70,31,70,30,41,31,185,31,172,31,172,30,117,31,117,30,51,31,51,30,207,31,91,31,91,30,139,31,6,31,6,30,6,29,82,31,254,31,254,30,143,31,182,31,206,31,21,31,5,31,72,31,92,31,211,31,182,31,178,31,116,31,221,31,83,31,174,31,219,31,219,30,247,31,120,31,49,31,224,31,145,31,145,30,202,31,243,31,238,31,215,31,215,30,215,29,215,28,215,27,215,26,192,31,22,31,22,30,94,31,94,30,144,31,209,31,51,31,101,31,101,30,254,31,125,31,138,31,164,31,141,31,253,31,180,31,210,31,48,31,62,31,62,30,221,31,221,30,91,31,225,31,225,30,75,31,12,31,221,31,120,31,84,31,94,31,163,31,18,31,120,31,67,31,67,30,167,31,164,31,71,31,171,31,171,30,171,29,108,31,18,31,74,31,109,31,61,31,28,31,170,31,119,31,10,31,254,31,224,31,196,31,47,31,47,30,247,31,61,31,61,30,68,31,8,31,108,31,108,30,192,31,141,31,141,30,173,31,97,31,3,31,99,31,99,30,99,29,179,31,143,31,3,31,62,31,46,31,46,30,103,31,192,31,217,31,38,31,36,31,37,31,152,31,9,31,9,30,44,31,11,31,100,31,180,31,30,31,139,31,36,31,62,31,62,30,62,29,198,31,50,31,50,30,50,29,37,31,210,31,210,30,44,31,107,31,205,31,205,30,3,31,102,31,2,31,21,31,142,31,186,31,109,31,116,31,224,31,125,31,252,31,31,31,98,31,233,31,14,31,14,30,24,31,7,31,157,31,46,31,46,30,42,31,102,31,102,30,213,31,197,31,197,30,100,31,192,31,210,31,184,31,80,31,179,31,179,30,1,31,59,31,196,31,231,31,244,31,50,31,11,31,11,30,176,31,8,31,8,30,33,31,170,31,170,30,170,29,163,31,60,31,60,30,156,31,225,31,120,31,163,31,188,31,50,31,148,31,148,30,252,31,178,31,178,30,97,31,97,30,97,29,83,31,198,31,91,31,193,31,180,31,122,31,139,31,220,31,123,31,9,31,15,31,35,31,213,31,216,31,247,31,102,31,225,31,92,31,246,31,246,30,226,31,226,30,220,31,50,31,140,31,86,31,82,31,115,31,98,31,124,31,13,31,186,31,165,31,73,31,45,31,153,31,153,30,235,31,150,31,117,31,140,31,133,31,133,30,133,29,92,31,92,30,241,31,71,31,123,31,123,30,230,31,249,31,82,31,147,31,97,31,132,31,60,31,94,31,4,31,213,31,32,31,5,31,5,30,104,31,124,31,230,31,77,31,162,31,162,30,44,31,213,31,213,30,198,31,47,31,124,31,184,31,152,31,58,31,58,30,58,29,169,31,219,31,126,31,32,31,32,30,119,31,119,30,119,29,40,31,200,31,31,31,226,31,226,30,189,31,26,31,213,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
