-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_947 is
end project_tb_947;

architecture project_tb_arch_947 of project_tb_947 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 597;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (235,0,15,0,119,0,82,0,70,0,102,0,113,0,117,0,223,0,0,0,0,0,28,0,193,0,164,0,168,0,2,0,50,0,23,0,197,0,0,0,0,0,223,0,32,0,229,0,254,0,173,0,21,0,26,0,0,0,5,0,181,0,145,0,203,0,140,0,195,0,61,0,48,0,6,0,120,0,213,0,121,0,0,0,188,0,0,0,242,0,36,0,250,0,222,0,16,0,0,0,114,0,162,0,47,0,195,0,6,0,0,0,67,0,156,0,0,0,62,0,82,0,6,0,0,0,176,0,127,0,113,0,88,0,223,0,157,0,230,0,30,0,123,0,0,0,187,0,0,0,47,0,153,0,254,0,0,0,236,0,50,0,0,0,156,0,78,0,0,0,167,0,200,0,55,0,206,0,203,0,93,0,62,0,187,0,0,0,32,0,102,0,151,0,206,0,0,0,5,0,240,0,0,0,227,0,70,0,101,0,170,0,229,0,0,0,207,0,250,0,174,0,173,0,0,0,0,0,79,0,9,0,88,0,160,0,34,0,84,0,63,0,147,0,85,0,68,0,109,0,42,0,11,0,255,0,221,0,0,0,87,0,0,0,86,0,210,0,113,0,85,0,41,0,94,0,142,0,42,0,207,0,172,0,113,0,0,0,0,0,53,0,166,0,0,0,128,0,127,0,142,0,27,0,191,0,86,0,219,0,197,0,201,0,0,0,0,0,143,0,148,0,76,0,113,0,0,0,2,0,43,0,156,0,17,0,107,0,147,0,188,0,29,0,0,0,166,0,0,0,231,0,92,0,0,0,153,0,46,0,0,0,241,0,35,0,83,0,0,0,0,0,0,0,78,0,116,0,122,0,69,0,178,0,231,0,29,0,0,0,188,0,146,0,253,0,56,0,173,0,189,0,56,0,151,0,27,0,4,0,0,0,61,0,206,0,112,0,59,0,152,0,149,0,43,0,87,0,49,0,238,0,103,0,21,0,6,0,125,0,138,0,169,0,234,0,54,0,171,0,4,0,245,0,0,0,56,0,110,0,211,0,0,0,249,0,60,0,92,0,250,0,0,0,181,0,91,0,96,0,153,0,58,0,48,0,164,0,4,0,114,0,84,0,67,0,55,0,0,0,229,0,0,0,7,0,0,0,0,0,67,0,0,0,0,0,218,0,129,0,151,0,7,0,5,0,206,0,64,0,17,0,98,0,191,0,0,0,195,0,68,0,197,0,169,0,4,0,0,0,90,0,166,0,0,0,184,0,246,0,67,0,199,0,92,0,147,0,169,0,97,0,251,0,0,0,93,0,232,0,21,0,95,0,0,0,36,0,3,0,0,0,0,0,110,0,169,0,101,0,0,0,0,0,55,0,46,0,97,0,252,0,19,0,184,0,11,0,7,0,21,0,0,0,61,0,35,0,0,0,75,0,217,0,112,0,215,0,206,0,0,0,143,0,0,0,184,0,102,0,90,0,105,0,2,0,190,0,74,0,0,0,0,0,172,0,158,0,184,0,200,0,0,0,160,0,1,0,106,0,0,0,0,0,53,0,0,0,0,0,0,0,155,0,0,0,237,0,149,0,142,0,243,0,11,0,4,0,219,0,55,0,103,0,33,0,201,0,243,0,129,0,219,0,226,0,10,0,150,0,41,0,119,0,0,0,47,0,241,0,236,0,237,0,145,0,255,0,0,0,0,0,88,0,0,0,156,0,166,0,99,0,101,0,253,0,128,0,111,0,208,0,77,0,160,0,83,0,0,0,0,0,209,0,0,0,0,0,197,0,175,0,217,0,186,0,0,0,242,0,0,0,152,0,0,0,116,0,0,0,0,0,194,0,71,0,127,0,148,0,25,0,0,0,79,0,69,0,24,0,0,0,80,0,99,0,246,0,244,0,0,0,0,0,72,0,132,0,146,0,0,0,39,0,214,0,0,0,252,0,0,0,215,0,0,0,49,0,143,0,226,0,18,0,222,0,159,0,113,0,199,0,199,0,228,0,240,0,90,0,0,0,0,0,76,0,0,0,40,0,242,0,78,0,203,0,0,0,84,0,214,0,170,0,0,0,0,0,50,0,0,0,112,0,0,0,0,0,2,0,206,0,0,0,125,0,134,0,112,0,233,0,44,0,0,0,6,0,103,0,39,0,121,0,0,0,115,0,93,0,27,0,0,0,0,0,177,0,197,0,119,0,0,0,0,0,0,0,154,0,165,0,135,0,41,0,214,0,0,0,0,0,0,0,0,0,57,0,85,0,0,0,69,0,13,0,243,0,0,0,23,0,164,0,0,0,43,0,49,0,5,0,0,0,0,0,237,0,0,0,0,0,0,0,225,0,202,0,0,0,228,0,77,0,125,0,126,0,121,0,0,0,253,0,0,0,0,0,178,0,118,0,0,0,54,0,9,0,0,0,205,0,46,0,208,0,176,0,0,0,20,0,45,0,225,0,0,0,0,0,12,0,0,0,246,0,125,0,245,0,134,0,128,0,231,0,6,0,167,0,133,0,134,0,145,0,86,0,84,0,38,0,191,0,0,0,202,0,123,0,218,0,112,0,0,0,51,0,174,0,5,0,16,0,131,0,245,0,0,0,136,0,18,0,0,0,170,0,184,0,92,0,216,0,167,0,187,0,6,0,246,0,3,0,93,0,0,0,63,0,140,0,41,0,202,0,57,0,105,0,235,0,194,0);
signal scenario_full  : scenario_type := (235,31,15,31,119,31,82,31,70,31,102,31,113,31,117,31,223,31,223,30,223,29,28,31,193,31,164,31,168,31,2,31,50,31,23,31,197,31,197,30,197,29,223,31,32,31,229,31,254,31,173,31,21,31,26,31,26,30,5,31,181,31,145,31,203,31,140,31,195,31,61,31,48,31,6,31,120,31,213,31,121,31,121,30,188,31,188,30,242,31,36,31,250,31,222,31,16,31,16,30,114,31,162,31,47,31,195,31,6,31,6,30,67,31,156,31,156,30,62,31,82,31,6,31,6,30,176,31,127,31,113,31,88,31,223,31,157,31,230,31,30,31,123,31,123,30,187,31,187,30,47,31,153,31,254,31,254,30,236,31,50,31,50,30,156,31,78,31,78,30,167,31,200,31,55,31,206,31,203,31,93,31,62,31,187,31,187,30,32,31,102,31,151,31,206,31,206,30,5,31,240,31,240,30,227,31,70,31,101,31,170,31,229,31,229,30,207,31,250,31,174,31,173,31,173,30,173,29,79,31,9,31,88,31,160,31,34,31,84,31,63,31,147,31,85,31,68,31,109,31,42,31,11,31,255,31,221,31,221,30,87,31,87,30,86,31,210,31,113,31,85,31,41,31,94,31,142,31,42,31,207,31,172,31,113,31,113,30,113,29,53,31,166,31,166,30,128,31,127,31,142,31,27,31,191,31,86,31,219,31,197,31,201,31,201,30,201,29,143,31,148,31,76,31,113,31,113,30,2,31,43,31,156,31,17,31,107,31,147,31,188,31,29,31,29,30,166,31,166,30,231,31,92,31,92,30,153,31,46,31,46,30,241,31,35,31,83,31,83,30,83,29,83,28,78,31,116,31,122,31,69,31,178,31,231,31,29,31,29,30,188,31,146,31,253,31,56,31,173,31,189,31,56,31,151,31,27,31,4,31,4,30,61,31,206,31,112,31,59,31,152,31,149,31,43,31,87,31,49,31,238,31,103,31,21,31,6,31,125,31,138,31,169,31,234,31,54,31,171,31,4,31,245,31,245,30,56,31,110,31,211,31,211,30,249,31,60,31,92,31,250,31,250,30,181,31,91,31,96,31,153,31,58,31,48,31,164,31,4,31,114,31,84,31,67,31,55,31,55,30,229,31,229,30,7,31,7,30,7,29,67,31,67,30,67,29,218,31,129,31,151,31,7,31,5,31,206,31,64,31,17,31,98,31,191,31,191,30,195,31,68,31,197,31,169,31,4,31,4,30,90,31,166,31,166,30,184,31,246,31,67,31,199,31,92,31,147,31,169,31,97,31,251,31,251,30,93,31,232,31,21,31,95,31,95,30,36,31,3,31,3,30,3,29,110,31,169,31,101,31,101,30,101,29,55,31,46,31,97,31,252,31,19,31,184,31,11,31,7,31,21,31,21,30,61,31,35,31,35,30,75,31,217,31,112,31,215,31,206,31,206,30,143,31,143,30,184,31,102,31,90,31,105,31,2,31,190,31,74,31,74,30,74,29,172,31,158,31,184,31,200,31,200,30,160,31,1,31,106,31,106,30,106,29,53,31,53,30,53,29,53,28,155,31,155,30,237,31,149,31,142,31,243,31,11,31,4,31,219,31,55,31,103,31,33,31,201,31,243,31,129,31,219,31,226,31,10,31,150,31,41,31,119,31,119,30,47,31,241,31,236,31,237,31,145,31,255,31,255,30,255,29,88,31,88,30,156,31,166,31,99,31,101,31,253,31,128,31,111,31,208,31,77,31,160,31,83,31,83,30,83,29,209,31,209,30,209,29,197,31,175,31,217,31,186,31,186,30,242,31,242,30,152,31,152,30,116,31,116,30,116,29,194,31,71,31,127,31,148,31,25,31,25,30,79,31,69,31,24,31,24,30,80,31,99,31,246,31,244,31,244,30,244,29,72,31,132,31,146,31,146,30,39,31,214,31,214,30,252,31,252,30,215,31,215,30,49,31,143,31,226,31,18,31,222,31,159,31,113,31,199,31,199,31,228,31,240,31,90,31,90,30,90,29,76,31,76,30,40,31,242,31,78,31,203,31,203,30,84,31,214,31,170,31,170,30,170,29,50,31,50,30,112,31,112,30,112,29,2,31,206,31,206,30,125,31,134,31,112,31,233,31,44,31,44,30,6,31,103,31,39,31,121,31,121,30,115,31,93,31,27,31,27,30,27,29,177,31,197,31,119,31,119,30,119,29,119,28,154,31,165,31,135,31,41,31,214,31,214,30,214,29,214,28,214,27,57,31,85,31,85,30,69,31,13,31,243,31,243,30,23,31,164,31,164,30,43,31,49,31,5,31,5,30,5,29,237,31,237,30,237,29,237,28,225,31,202,31,202,30,228,31,77,31,125,31,126,31,121,31,121,30,253,31,253,30,253,29,178,31,118,31,118,30,54,31,9,31,9,30,205,31,46,31,208,31,176,31,176,30,20,31,45,31,225,31,225,30,225,29,12,31,12,30,246,31,125,31,245,31,134,31,128,31,231,31,6,31,167,31,133,31,134,31,145,31,86,31,84,31,38,31,191,31,191,30,202,31,123,31,218,31,112,31,112,30,51,31,174,31,5,31,16,31,131,31,245,31,245,30,136,31,18,31,18,30,170,31,184,31,92,31,216,31,167,31,187,31,6,31,246,31,3,31,93,31,93,30,63,31,140,31,41,31,202,31,57,31,105,31,235,31,194,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
