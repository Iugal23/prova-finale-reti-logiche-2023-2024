-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 235;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,19,0,101,0,209,0,104,0,0,0,222,0,2,0,110,0,119,0,177,0,144,0,98,0,18,0,128,0,172,0,0,0,0,0,196,0,0,0,32,0,122,0,194,0,231,0,2,0,70,0,67,0,170,0,56,0,107,0,0,0,207,0,8,0,38,0,246,0,78,0,156,0,214,0,148,0,57,0,166,0,87,0,0,0,197,0,235,0,72,0,0,0,156,0,0,0,148,0,0,0,0,0,181,0,183,0,0,0,88,0,180,0,150,0,199,0,183,0,0,0,20,0,157,0,252,0,0,0,79,0,0,0,195,0,70,0,91,0,45,0,0,0,67,0,135,0,206,0,153,0,172,0,218,0,181,0,19,0,102,0,190,0,246,0,208,0,156,0,0,0,171,0,231,0,63,0,59,0,145,0,15,0,4,0,0,0,225,0,55,0,52,0,0,0,26,0,89,0,35,0,0,0,134,0,92,0,140,0,0,0,112,0,159,0,235,0,215,0,220,0,0,0,196,0,118,0,215,0,129,0,253,0,7,0,0,0,252,0,0,0,17,0,132,0,185,0,15,0,186,0,0,0,93,0,0,0,43,0,0,0,181,0,0,0,137,0,20,0,42,0,0,0,93,0,0,0,102,0,6,0,155,0,13,0,194,0,167,0,253,0,241,0,0,0,137,0,44,0,94,0,0,0,196,0,166,0,185,0,217,0,181,0,117,0,183,0,5,0,205,0,65,0,136,0,3,0,0,0,0,0,58,0,97,0,88,0,0,0,119,0,170,0,240,0,79,0,233,0,108,0,27,0,0,0,95,0,47,0,252,0,106,0,140,0,251,0,142,0,73,0,223,0,229,0,205,0,248,0,150,0,253,0,0,0,150,0,143,0,236,0,156,0,0,0,191,0,220,0,161,0,159,0,200,0,0,0,158,0,231,0,92,0,151,0,84,0,49,0,105,0,201,0,253,0,217,0,0,0,217,0,5,0,90,0,0,0,61,0,221,0,81,0,186,0,93,0,193,0,10,0,46,0,201,0,112,0,67,0,244,0,153,0,57,0,89,0,91,0);
signal scenario_full  : scenario_type := (0,0,19,31,101,31,209,31,104,31,104,30,222,31,2,31,110,31,119,31,177,31,144,31,98,31,18,31,128,31,172,31,172,30,172,29,196,31,196,30,32,31,122,31,194,31,231,31,2,31,70,31,67,31,170,31,56,31,107,31,107,30,207,31,8,31,38,31,246,31,78,31,156,31,214,31,148,31,57,31,166,31,87,31,87,30,197,31,235,31,72,31,72,30,156,31,156,30,148,31,148,30,148,29,181,31,183,31,183,30,88,31,180,31,150,31,199,31,183,31,183,30,20,31,157,31,252,31,252,30,79,31,79,30,195,31,70,31,91,31,45,31,45,30,67,31,135,31,206,31,153,31,172,31,218,31,181,31,19,31,102,31,190,31,246,31,208,31,156,31,156,30,171,31,231,31,63,31,59,31,145,31,15,31,4,31,4,30,225,31,55,31,52,31,52,30,26,31,89,31,35,31,35,30,134,31,92,31,140,31,140,30,112,31,159,31,235,31,215,31,220,31,220,30,196,31,118,31,215,31,129,31,253,31,7,31,7,30,252,31,252,30,17,31,132,31,185,31,15,31,186,31,186,30,93,31,93,30,43,31,43,30,181,31,181,30,137,31,20,31,42,31,42,30,93,31,93,30,102,31,6,31,155,31,13,31,194,31,167,31,253,31,241,31,241,30,137,31,44,31,94,31,94,30,196,31,166,31,185,31,217,31,181,31,117,31,183,31,5,31,205,31,65,31,136,31,3,31,3,30,3,29,58,31,97,31,88,31,88,30,119,31,170,31,240,31,79,31,233,31,108,31,27,31,27,30,95,31,47,31,252,31,106,31,140,31,251,31,142,31,73,31,223,31,229,31,205,31,248,31,150,31,253,31,253,30,150,31,143,31,236,31,156,31,156,30,191,31,220,31,161,31,159,31,200,31,200,30,158,31,231,31,92,31,151,31,84,31,49,31,105,31,201,31,253,31,217,31,217,30,217,31,5,31,90,31,90,30,61,31,221,31,81,31,186,31,93,31,193,31,10,31,46,31,201,31,112,31,67,31,244,31,153,31,57,31,89,31,91,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
