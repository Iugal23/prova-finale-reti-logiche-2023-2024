-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_965 is
end project_tb_965;

architecture project_tb_arch_965 of project_tb_965 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 649;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (7,0,10,0,237,0,137,0,0,0,118,0,146,0,133,0,59,0,228,0,203,0,104,0,246,0,0,0,224,0,0,0,160,0,42,0,245,0,16,0,0,0,224,0,36,0,125,0,58,0,157,0,149,0,35,0,222,0,209,0,192,0,71,0,228,0,0,0,0,0,233,0,50,0,193,0,0,0,19,0,236,0,15,0,201,0,96,0,0,0,121,0,0,0,97,0,189,0,180,0,57,0,111,0,65,0,216,0,133,0,222,0,59,0,0,0,250,0,222,0,92,0,0,0,85,0,75,0,0,0,75,0,40,0,63,0,180,0,240,0,0,0,20,0,159,0,0,0,0,0,48,0,179,0,234,0,93,0,33,0,24,0,0,0,100,0,194,0,70,0,123,0,187,0,0,0,143,0,0,0,168,0,54,0,0,0,215,0,13,0,155,0,115,0,110,0,239,0,157,0,51,0,208,0,222,0,237,0,127,0,188,0,131,0,140,0,38,0,81,0,109,0,2,0,126,0,75,0,34,0,98,0,33,0,0,0,0,0,108,0,235,0,190,0,0,0,149,0,92,0,52,0,236,0,99,0,0,0,75,0,129,0,55,0,33,0,110,0,189,0,0,0,54,0,253,0,97,0,0,0,113,0,191,0,0,0,157,0,200,0,119,0,126,0,105,0,39,0,116,0,228,0,0,0,22,0,190,0,97,0,129,0,0,0,0,0,170,0,0,0,59,0,135,0,228,0,0,0,122,0,208,0,94,0,0,0,221,0,0,0,81,0,74,0,105,0,31,0,167,0,140,0,0,0,38,0,167,0,197,0,82,0,210,0,252,0,13,0,215,0,231,0,135,0,121,0,158,0,177,0,12,0,128,0,0,0,183,0,224,0,0,0,134,0,178,0,58,0,191,0,66,0,0,0,248,0,35,0,178,0,219,0,0,0,138,0,90,0,253,0,160,0,106,0,232,0,170,0,154,0,124,0,152,0,23,0,142,0,0,0,106,0,238,0,213,0,0,0,65,0,88,0,115,0,167,0,155,0,15,0,0,0,217,0,5,0,38,0,34,0,148,0,86,0,169,0,111,0,102,0,130,0,245,0,133,0,0,0,96,0,82,0,121,0,0,0,138,0,0,0,177,0,2,0,56,0,49,0,166,0,3,0,98,0,198,0,48,0,3,0,176,0,173,0,92,0,253,0,0,0,188,0,0,0,0,0,67,0,120,0,172,0,22,0,13,0,47,0,162,0,219,0,106,0,34,0,15,0,98,0,115,0,189,0,15,0,123,0,18,0,241,0,0,0,0,0,203,0,54,0,173,0,212,0,0,0,44,0,232,0,0,0,219,0,0,0,185,0,187,0,191,0,172,0,243,0,235,0,226,0,106,0,112,0,31,0,250,0,0,0,91,0,72,0,106,0,8,0,131,0,127,0,184,0,75,0,169,0,247,0,65,0,222,0,33,0,0,0,157,0,161,0,176,0,57,0,216,0,204,0,46,0,0,0,162,0,220,0,3,0,0,0,206,0,0,0,217,0,26,0,80,0,107,0,165,0,49,0,231,0,87,0,28,0,6,0,0,0,225,0,60,0,60,0,0,0,50,0,105,0,0,0,216,0,49,0,0,0,82,0,163,0,116,0,26,0,190,0,137,0,61,0,0,0,154,0,0,0,164,0,90,0,0,0,49,0,216,0,102,0,39,0,204,0,145,0,99,0,34,0,94,0,152,0,150,0,248,0,0,0,249,0,162,0,67,0,18,0,0,0,111,0,117,0,0,0,54,0,73,0,178,0,25,0,19,0,0,0,0,0,125,0,64,0,71,0,51,0,144,0,248,0,0,0,55,0,218,0,57,0,84,0,80,0,18,0,130,0,152,0,161,0,0,0,46,0,149,0,244,0,12,0,57,0,52,0,67,0,224,0,79,0,118,0,163,0,0,0,236,0,193,0,159,0,164,0,185,0,226,0,195,0,181,0,205,0,0,0,193,0,0,0,19,0,98,0,0,0,136,0,200,0,0,0,0,0,16,0,47,0,0,0,121,0,2,0,139,0,0,0,234,0,0,0,112,0,150,0,223,0,0,0,0,0,0,0,86,0,203,0,200,0,27,0,162,0,183,0,122,0,15,0,89,0,0,0,119,0,0,0,199,0,0,0,72,0,190,0,0,0,93,0,78,0,0,0,0,0,168,0,0,0,155,0,251,0,239,0,182,0,45,0,241,0,183,0,198,0,121,0,0,0,21,0,63,0,156,0,176,0,159,0,0,0,150,0,48,0,223,0,0,0,45,0,248,0,17,0,85,0,162,0,15,0,30,0,122,0,65,0,243,0,0,0,0,0,161,0,214,0,201,0,0,0,215,0,80,0,0,0,0,0,0,0,0,0,221,0,66,0,237,0,199,0,153,0,150,0,0,0,111,0,14,0,1,0,36,0,110,0,88,0,156,0,22,0,158,0,0,0,181,0,0,0,60,0,0,0,58,0,73,0,0,0,0,0,159,0,1,0,0,0,255,0,90,0,33,0,92,0,107,0,8,0,99,0,117,0,0,0,16,0,227,0,129,0,117,0,204,0,124,0,36,0,29,0,0,0,123,0,51,0,227,0,0,0,0,0,65,0,225,0,76,0,226,0,33,0,192,0,0,0,16,0,166,0,234,0,29,0,20,0,0,0,33,0,87,0,45,0,147,0,0,0,0,0,0,0,76,0,70,0,0,0,209,0,141,0,238,0,124,0,0,0,147,0,160,0,225,0,8,0,78,0,108,0,157,0,121,0,58,0,221,0,83,0,71,0,154,0,2,0,24,0,157,0,184,0,110,0,30,0,0,0,207,0,129,0,135,0,123,0,200,0,41,0,0,0,0,0,100,0,220,0,143,0,244,0,230,0,131,0,0,0,250,0,236,0,25,0,131,0,24,0,24,0,170,0);
signal scenario_full  : scenario_type := (7,31,10,31,237,31,137,31,137,30,118,31,146,31,133,31,59,31,228,31,203,31,104,31,246,31,246,30,224,31,224,30,160,31,42,31,245,31,16,31,16,30,224,31,36,31,125,31,58,31,157,31,149,31,35,31,222,31,209,31,192,31,71,31,228,31,228,30,228,29,233,31,50,31,193,31,193,30,19,31,236,31,15,31,201,31,96,31,96,30,121,31,121,30,97,31,189,31,180,31,57,31,111,31,65,31,216,31,133,31,222,31,59,31,59,30,250,31,222,31,92,31,92,30,85,31,75,31,75,30,75,31,40,31,63,31,180,31,240,31,240,30,20,31,159,31,159,30,159,29,48,31,179,31,234,31,93,31,33,31,24,31,24,30,100,31,194,31,70,31,123,31,187,31,187,30,143,31,143,30,168,31,54,31,54,30,215,31,13,31,155,31,115,31,110,31,239,31,157,31,51,31,208,31,222,31,237,31,127,31,188,31,131,31,140,31,38,31,81,31,109,31,2,31,126,31,75,31,34,31,98,31,33,31,33,30,33,29,108,31,235,31,190,31,190,30,149,31,92,31,52,31,236,31,99,31,99,30,75,31,129,31,55,31,33,31,110,31,189,31,189,30,54,31,253,31,97,31,97,30,113,31,191,31,191,30,157,31,200,31,119,31,126,31,105,31,39,31,116,31,228,31,228,30,22,31,190,31,97,31,129,31,129,30,129,29,170,31,170,30,59,31,135,31,228,31,228,30,122,31,208,31,94,31,94,30,221,31,221,30,81,31,74,31,105,31,31,31,167,31,140,31,140,30,38,31,167,31,197,31,82,31,210,31,252,31,13,31,215,31,231,31,135,31,121,31,158,31,177,31,12,31,128,31,128,30,183,31,224,31,224,30,134,31,178,31,58,31,191,31,66,31,66,30,248,31,35,31,178,31,219,31,219,30,138,31,90,31,253,31,160,31,106,31,232,31,170,31,154,31,124,31,152,31,23,31,142,31,142,30,106,31,238,31,213,31,213,30,65,31,88,31,115,31,167,31,155,31,15,31,15,30,217,31,5,31,38,31,34,31,148,31,86,31,169,31,111,31,102,31,130,31,245,31,133,31,133,30,96,31,82,31,121,31,121,30,138,31,138,30,177,31,2,31,56,31,49,31,166,31,3,31,98,31,198,31,48,31,3,31,176,31,173,31,92,31,253,31,253,30,188,31,188,30,188,29,67,31,120,31,172,31,22,31,13,31,47,31,162,31,219,31,106,31,34,31,15,31,98,31,115,31,189,31,15,31,123,31,18,31,241,31,241,30,241,29,203,31,54,31,173,31,212,31,212,30,44,31,232,31,232,30,219,31,219,30,185,31,187,31,191,31,172,31,243,31,235,31,226,31,106,31,112,31,31,31,250,31,250,30,91,31,72,31,106,31,8,31,131,31,127,31,184,31,75,31,169,31,247,31,65,31,222,31,33,31,33,30,157,31,161,31,176,31,57,31,216,31,204,31,46,31,46,30,162,31,220,31,3,31,3,30,206,31,206,30,217,31,26,31,80,31,107,31,165,31,49,31,231,31,87,31,28,31,6,31,6,30,225,31,60,31,60,31,60,30,50,31,105,31,105,30,216,31,49,31,49,30,82,31,163,31,116,31,26,31,190,31,137,31,61,31,61,30,154,31,154,30,164,31,90,31,90,30,49,31,216,31,102,31,39,31,204,31,145,31,99,31,34,31,94,31,152,31,150,31,248,31,248,30,249,31,162,31,67,31,18,31,18,30,111,31,117,31,117,30,54,31,73,31,178,31,25,31,19,31,19,30,19,29,125,31,64,31,71,31,51,31,144,31,248,31,248,30,55,31,218,31,57,31,84,31,80,31,18,31,130,31,152,31,161,31,161,30,46,31,149,31,244,31,12,31,57,31,52,31,67,31,224,31,79,31,118,31,163,31,163,30,236,31,193,31,159,31,164,31,185,31,226,31,195,31,181,31,205,31,205,30,193,31,193,30,19,31,98,31,98,30,136,31,200,31,200,30,200,29,16,31,47,31,47,30,121,31,2,31,139,31,139,30,234,31,234,30,112,31,150,31,223,31,223,30,223,29,223,28,86,31,203,31,200,31,27,31,162,31,183,31,122,31,15,31,89,31,89,30,119,31,119,30,199,31,199,30,72,31,190,31,190,30,93,31,78,31,78,30,78,29,168,31,168,30,155,31,251,31,239,31,182,31,45,31,241,31,183,31,198,31,121,31,121,30,21,31,63,31,156,31,176,31,159,31,159,30,150,31,48,31,223,31,223,30,45,31,248,31,17,31,85,31,162,31,15,31,30,31,122,31,65,31,243,31,243,30,243,29,161,31,214,31,201,31,201,30,215,31,80,31,80,30,80,29,80,28,80,27,221,31,66,31,237,31,199,31,153,31,150,31,150,30,111,31,14,31,1,31,36,31,110,31,88,31,156,31,22,31,158,31,158,30,181,31,181,30,60,31,60,30,58,31,73,31,73,30,73,29,159,31,1,31,1,30,255,31,90,31,33,31,92,31,107,31,8,31,99,31,117,31,117,30,16,31,227,31,129,31,117,31,204,31,124,31,36,31,29,31,29,30,123,31,51,31,227,31,227,30,227,29,65,31,225,31,76,31,226,31,33,31,192,31,192,30,16,31,166,31,234,31,29,31,20,31,20,30,33,31,87,31,45,31,147,31,147,30,147,29,147,28,76,31,70,31,70,30,209,31,141,31,238,31,124,31,124,30,147,31,160,31,225,31,8,31,78,31,108,31,157,31,121,31,58,31,221,31,83,31,71,31,154,31,2,31,24,31,157,31,184,31,110,31,30,31,30,30,207,31,129,31,135,31,123,31,200,31,41,31,41,30,41,29,100,31,220,31,143,31,244,31,230,31,131,31,131,30,250,31,236,31,25,31,131,31,24,31,24,31,170,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
