-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_80 is
end project_tb_80;

architecture project_tb_arch_80 of project_tb_80 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 417;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (4,0,111,0,57,0,0,0,155,0,161,0,67,0,119,0,22,0,0,0,178,0,128,0,8,0,138,0,5,0,134,0,221,0,211,0,1,0,140,0,70,0,231,0,0,0,101,0,0,0,148,0,58,0,0,0,198,0,0,0,0,0,109,0,0,0,0,0,63,0,44,0,129,0,235,0,0,0,190,0,139,0,0,0,171,0,126,0,173,0,0,0,0,0,0,0,0,0,86,0,50,0,222,0,84,0,223,0,210,0,163,0,115,0,81,0,163,0,209,0,0,0,206,0,247,0,132,0,68,0,99,0,162,0,33,0,0,0,186,0,28,0,200,0,246,0,67,0,33,0,238,0,220,0,189,0,207,0,135,0,136,0,179,0,162,0,148,0,30,0,0,0,229,0,0,0,200,0,200,0,162,0,157,0,47,0,34,0,0,0,85,0,30,0,77,0,30,0,242,0,138,0,1,0,88,0,237,0,65,0,238,0,50,0,192,0,246,0,58,0,32,0,0,0,170,0,66,0,156,0,83,0,212,0,0,0,48,0,6,0,0,0,100,0,250,0,49,0,45,0,185,0,69,0,152,0,114,0,122,0,109,0,203,0,182,0,223,0,116,0,46,0,129,0,0,0,175,0,87,0,143,0,202,0,101,0,52,0,179,0,40,0,0,0,170,0,235,0,94,0,69,0,74,0,162,0,43,0,10,0,199,0,155,0,99,0,0,0,243,0,88,0,60,0,160,0,159,0,207,0,0,0,0,0,117,0,186,0,201,0,172,0,0,0,103,0,127,0,0,0,11,0,9,0,58,0,148,0,25,0,127,0,64,0,234,0,197,0,0,0,0,0,250,0,53,0,236,0,39,0,0,0,202,0,0,0,241,0,156,0,139,0,0,0,237,0,211,0,32,0,145,0,35,0,0,0,242,0,130,0,97,0,0,0,248,0,17,0,204,0,11,0,76,0,29,0,233,0,19,0,52,0,26,0,190,0,70,0,0,0,187,0,146,0,69,0,240,0,173,0,0,0,21,0,97,0,0,0,221,0,41,0,23,0,156,0,0,0,165,0,0,0,221,0,26,0,74,0,131,0,48,0,225,0,84,0,117,0,40,0,97,0,145,0,87,0,0,0,127,0,180,0,1,0,78,0,27,0,78,0,84,0,119,0,158,0,249,0,35,0,62,0,82,0,166,0,117,0,4,0,228,0,142,0,3,0,191,0,0,0,159,0,29,0,179,0,218,0,26,0,180,0,252,0,241,0,0,0,203,0,172,0,62,0,159,0,171,0,0,0,0,0,129,0,11,0,0,0,237,0,0,0,182,0,194,0,74,0,0,0,94,0,150,0,171,0,14,0,93,0,195,0,147,0,236,0,99,0,218,0,110,0,194,0,0,0,85,0,0,0,47,0,154,0,196,0,234,0,53,0,237,0,252,0,114,0,20,0,202,0,45,0,132,0,222,0,93,0,0,0,0,0,89,0,207,0,0,0,148,0,0,0,118,0,81,0,11,0,0,0,0,0,76,0,113,0,160,0,52,0,0,0,195,0,0,0,193,0,129,0,0,0,49,0,0,0,87,0,30,0,149,0,0,0,63,0,180,0,208,0,52,0,241,0,33,0,118,0,52,0,162,0,185,0,28,0,82,0,150,0,26,0,0,0,20,0,14,0,235,0,84,0,0,0,223,0,176,0,0,0,232,0,77,0,86,0,30,0,223,0,32,0,246,0,225,0,0,0,80,0,115,0,163,0,29,0,45,0,225,0,143,0,101,0,189,0,217,0,54,0,28,0,41,0,0,0,3,0,32,0,177,0,0,0,0,0,51,0,0,0,17,0,176,0,0,0,188,0,170,0,23,0,192,0,45,0,0,0,215,0,0,0,112,0);
signal scenario_full  : scenario_type := (4,31,111,31,57,31,57,30,155,31,161,31,67,31,119,31,22,31,22,30,178,31,128,31,8,31,138,31,5,31,134,31,221,31,211,31,1,31,140,31,70,31,231,31,231,30,101,31,101,30,148,31,58,31,58,30,198,31,198,30,198,29,109,31,109,30,109,29,63,31,44,31,129,31,235,31,235,30,190,31,139,31,139,30,171,31,126,31,173,31,173,30,173,29,173,28,173,27,86,31,50,31,222,31,84,31,223,31,210,31,163,31,115,31,81,31,163,31,209,31,209,30,206,31,247,31,132,31,68,31,99,31,162,31,33,31,33,30,186,31,28,31,200,31,246,31,67,31,33,31,238,31,220,31,189,31,207,31,135,31,136,31,179,31,162,31,148,31,30,31,30,30,229,31,229,30,200,31,200,31,162,31,157,31,47,31,34,31,34,30,85,31,30,31,77,31,30,31,242,31,138,31,1,31,88,31,237,31,65,31,238,31,50,31,192,31,246,31,58,31,32,31,32,30,170,31,66,31,156,31,83,31,212,31,212,30,48,31,6,31,6,30,100,31,250,31,49,31,45,31,185,31,69,31,152,31,114,31,122,31,109,31,203,31,182,31,223,31,116,31,46,31,129,31,129,30,175,31,87,31,143,31,202,31,101,31,52,31,179,31,40,31,40,30,170,31,235,31,94,31,69,31,74,31,162,31,43,31,10,31,199,31,155,31,99,31,99,30,243,31,88,31,60,31,160,31,159,31,207,31,207,30,207,29,117,31,186,31,201,31,172,31,172,30,103,31,127,31,127,30,11,31,9,31,58,31,148,31,25,31,127,31,64,31,234,31,197,31,197,30,197,29,250,31,53,31,236,31,39,31,39,30,202,31,202,30,241,31,156,31,139,31,139,30,237,31,211,31,32,31,145,31,35,31,35,30,242,31,130,31,97,31,97,30,248,31,17,31,204,31,11,31,76,31,29,31,233,31,19,31,52,31,26,31,190,31,70,31,70,30,187,31,146,31,69,31,240,31,173,31,173,30,21,31,97,31,97,30,221,31,41,31,23,31,156,31,156,30,165,31,165,30,221,31,26,31,74,31,131,31,48,31,225,31,84,31,117,31,40,31,97,31,145,31,87,31,87,30,127,31,180,31,1,31,78,31,27,31,78,31,84,31,119,31,158,31,249,31,35,31,62,31,82,31,166,31,117,31,4,31,228,31,142,31,3,31,191,31,191,30,159,31,29,31,179,31,218,31,26,31,180,31,252,31,241,31,241,30,203,31,172,31,62,31,159,31,171,31,171,30,171,29,129,31,11,31,11,30,237,31,237,30,182,31,194,31,74,31,74,30,94,31,150,31,171,31,14,31,93,31,195,31,147,31,236,31,99,31,218,31,110,31,194,31,194,30,85,31,85,30,47,31,154,31,196,31,234,31,53,31,237,31,252,31,114,31,20,31,202,31,45,31,132,31,222,31,93,31,93,30,93,29,89,31,207,31,207,30,148,31,148,30,118,31,81,31,11,31,11,30,11,29,76,31,113,31,160,31,52,31,52,30,195,31,195,30,193,31,129,31,129,30,49,31,49,30,87,31,30,31,149,31,149,30,63,31,180,31,208,31,52,31,241,31,33,31,118,31,52,31,162,31,185,31,28,31,82,31,150,31,26,31,26,30,20,31,14,31,235,31,84,31,84,30,223,31,176,31,176,30,232,31,77,31,86,31,30,31,223,31,32,31,246,31,225,31,225,30,80,31,115,31,163,31,29,31,45,31,225,31,143,31,101,31,189,31,217,31,54,31,28,31,41,31,41,30,3,31,32,31,177,31,177,30,177,29,51,31,51,30,17,31,176,31,176,30,188,31,170,31,23,31,192,31,45,31,45,30,215,31,215,30,112,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
