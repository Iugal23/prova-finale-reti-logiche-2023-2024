-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_303 is
end project_tb_303;

architecture project_tb_arch_303 of project_tb_303 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 669;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (102,0,215,0,101,0,237,0,0,0,167,0,61,0,0,0,0,0,37,0,66,0,235,0,117,0,197,0,0,0,0,0,9,0,180,0,151,0,57,0,49,0,0,0,84,0,51,0,0,0,93,0,44,0,9,0,0,0,61,0,151,0,181,0,148,0,146,0,17,0,0,0,0,0,99,0,1,0,142,0,97,0,84,0,123,0,99,0,0,0,93,0,29,0,155,0,91,0,98,0,116,0,2,0,145,0,134,0,31,0,158,0,0,0,218,0,0,0,252,0,177,0,127,0,0,0,116,0,153,0,86,0,69,0,53,0,61,0,0,0,249,0,161,0,12,0,180,0,18,0,53,0,39,0,156,0,202,0,137,0,95,0,0,0,237,0,47,0,129,0,144,0,50,0,243,0,129,0,122,0,230,0,226,0,0,0,122,0,207,0,98,0,0,0,0,0,9,0,103,0,0,0,233,0,0,0,204,0,48,0,121,0,0,0,112,0,81,0,161,0,231,0,132,0,186,0,250,0,72,0,58,0,242,0,70,0,0,0,123,0,48,0,242,0,239,0,204,0,147,0,188,0,167,0,146,0,198,0,0,0,209,0,245,0,153,0,0,0,0,0,224,0,236,0,211,0,3,0,152,0,0,0,150,0,117,0,0,0,0,0,143,0,166,0,49,0,197,0,191,0,2,0,4,0,201,0,211,0,210,0,199,0,18,0,124,0,194,0,35,0,0,0,188,0,0,0,132,0,228,0,141,0,92,0,148,0,186,0,1,0,18,0,0,0,86,0,24,0,173,0,74,0,138,0,0,0,239,0,0,0,58,0,91,0,86,0,59,0,173,0,85,0,210,0,27,0,235,0,0,0,77,0,0,0,16,0,204,0,226,0,227,0,184,0,240,0,0,0,85,0,0,0,0,0,0,0,137,0,0,0,0,0,0,0,62,0,22,0,93,0,192,0,61,0,54,0,185,0,133,0,0,0,1,0,180,0,124,0,159,0,107,0,52,0,244,0,235,0,54,0,29,0,75,0,0,0,0,0,251,0,248,0,27,0,245,0,0,0,86,0,150,0,241,0,225,0,43,0,85,0,147,0,148,0,0,0,6,0,0,0,53,0,86,0,0,0,242,0,255,0,210,0,4,0,10,0,255,0,147,0,78,0,248,0,24,0,131,0,74,0,125,0,0,0,213,0,114,0,116,0,25,0,142,0,221,0,213,0,205,0,66,0,253,0,9,0,0,0,211,0,250,0,231,0,0,0,251,0,121,0,151,0,33,0,106,0,130,0,0,0,245,0,60,0,0,0,136,0,57,0,103,0,246,0,111,0,104,0,39,0,143,0,161,0,7,0,76,0,199,0,124,0,74,0,45,0,180,0,88,0,215,0,207,0,84,0,0,0,0,0,0,0,80,0,0,0,206,0,255,0,0,0,170,0,231,0,207,0,93,0,160,0,30,0,0,0,242,0,180,0,217,0,228,0,37,0,170,0,238,0,0,0,127,0,58,0,96,0,134,0,62,0,200,0,225,0,76,0,134,0,91,0,189,0,17,0,0,0,207,0,98,0,78,0,136,0,150,0,42,0,60,0,96,0,213,0,31,0,223,0,232,0,37,0,112,0,0,0,0,0,237,0,248,0,187,0,83,0,34,0,159,0,0,0,243,0,197,0,93,0,141,0,0,0,9,0,121,0,82,0,247,0,15,0,35,0,66,0,128,0,0,0,198,0,71,0,182,0,115,0,227,0,164,0,166,0,1,0,154,0,230,0,63,0,53,0,149,0,123,0,184,0,93,0,0,0,215,0,14,0,132,0,206,0,154,0,205,0,239,0,15,0,142,0,212,0,33,0,210,0,229,0,0,0,126,0,0,0,42,0,42,0,186,0,224,0,176,0,0,0,185,0,233,0,127,0,54,0,0,0,206,0,167,0,104,0,94,0,27,0,5,0,243,0,150,0,115,0,206,0,0,0,206,0,174,0,0,0,0,0,203,0,117,0,57,0,85,0,57,0,104,0,222,0,88,0,43,0,0,0,234,0,94,0,125,0,198,0,147,0,0,0,0,0,76,0,0,0,12,0,0,0,0,0,0,0,44,0,156,0,100,0,35,0,180,0,233,0,248,0,114,0,0,0,0,0,0,0,157,0,165,0,202,0,0,0,122,0,64,0,242,0,0,0,0,0,26,0,13,0,221,0,28,0,0,0,0,0,159,0,0,0,213,0,152,0,175,0,199,0,151,0,136,0,28,0,49,0,0,0,234,0,214,0,0,0,42,0,200,0,18,0,0,0,8,0,21,0,6,0,151,0,17,0,253,0,48,0,128,0,0,0,222,0,180,0,84,0,0,0,193,0,0,0,19,0,226,0,101,0,0,0,44,0,48,0,164,0,122,0,223,0,0,0,0,0,71,0,0,0,135,0,56,0,89,0,167,0,0,0,0,0,210,0,158,0,137,0,87,0,38,0,19,0,0,0,214,0,0,0,210,0,184,0,160,0,197,0,185,0,109,0,0,0,238,0,0,0,0,0,208,0,15,0,65,0,139,0,0,0,166,0,122,0,208,0,138,0,103,0,175,0,0,0,96,0,39,0,163,0,195,0,26,0,0,0,180,0,240,0,147,0,0,0,213,0,76,0,51,0,95,0,171,0,0,0,248,0,238,0,117,0,118,0,51,0,18,0,169,0,52,0,164,0,138,0,27,0,190,0,203,0,34,0,0,0,64,0,141,0,81,0,34,0,27,0,134,0,156,0,243,0,109,0,233,0,164,0,67,0,233,0,226,0,6,0,233,0,93,0,183,0,238,0,61,0,153,0,146,0,122,0,223,0,0,0,0,0,121,0,190,0,117,0,123,0,174,0,233,0,176,0,239,0,107,0,3,0,178,0,1,0,0,0,0,0,250,0,213,0,19,0,2,0,189,0,50,0,247,0,104,0,108,0,123,0,153,0,0,0,193,0,171,0,249,0,165,0,108,0,0,0,76,0,239,0,146,0,136,0,113,0,0,0,49,0,0,0);
signal scenario_full  : scenario_type := (102,31,215,31,101,31,237,31,237,30,167,31,61,31,61,30,61,29,37,31,66,31,235,31,117,31,197,31,197,30,197,29,9,31,180,31,151,31,57,31,49,31,49,30,84,31,51,31,51,30,93,31,44,31,9,31,9,30,61,31,151,31,181,31,148,31,146,31,17,31,17,30,17,29,99,31,1,31,142,31,97,31,84,31,123,31,99,31,99,30,93,31,29,31,155,31,91,31,98,31,116,31,2,31,145,31,134,31,31,31,158,31,158,30,218,31,218,30,252,31,177,31,127,31,127,30,116,31,153,31,86,31,69,31,53,31,61,31,61,30,249,31,161,31,12,31,180,31,18,31,53,31,39,31,156,31,202,31,137,31,95,31,95,30,237,31,47,31,129,31,144,31,50,31,243,31,129,31,122,31,230,31,226,31,226,30,122,31,207,31,98,31,98,30,98,29,9,31,103,31,103,30,233,31,233,30,204,31,48,31,121,31,121,30,112,31,81,31,161,31,231,31,132,31,186,31,250,31,72,31,58,31,242,31,70,31,70,30,123,31,48,31,242,31,239,31,204,31,147,31,188,31,167,31,146,31,198,31,198,30,209,31,245,31,153,31,153,30,153,29,224,31,236,31,211,31,3,31,152,31,152,30,150,31,117,31,117,30,117,29,143,31,166,31,49,31,197,31,191,31,2,31,4,31,201,31,211,31,210,31,199,31,18,31,124,31,194,31,35,31,35,30,188,31,188,30,132,31,228,31,141,31,92,31,148,31,186,31,1,31,18,31,18,30,86,31,24,31,173,31,74,31,138,31,138,30,239,31,239,30,58,31,91,31,86,31,59,31,173,31,85,31,210,31,27,31,235,31,235,30,77,31,77,30,16,31,204,31,226,31,227,31,184,31,240,31,240,30,85,31,85,30,85,29,85,28,137,31,137,30,137,29,137,28,62,31,22,31,93,31,192,31,61,31,54,31,185,31,133,31,133,30,1,31,180,31,124,31,159,31,107,31,52,31,244,31,235,31,54,31,29,31,75,31,75,30,75,29,251,31,248,31,27,31,245,31,245,30,86,31,150,31,241,31,225,31,43,31,85,31,147,31,148,31,148,30,6,31,6,30,53,31,86,31,86,30,242,31,255,31,210,31,4,31,10,31,255,31,147,31,78,31,248,31,24,31,131,31,74,31,125,31,125,30,213,31,114,31,116,31,25,31,142,31,221,31,213,31,205,31,66,31,253,31,9,31,9,30,211,31,250,31,231,31,231,30,251,31,121,31,151,31,33,31,106,31,130,31,130,30,245,31,60,31,60,30,136,31,57,31,103,31,246,31,111,31,104,31,39,31,143,31,161,31,7,31,76,31,199,31,124,31,74,31,45,31,180,31,88,31,215,31,207,31,84,31,84,30,84,29,84,28,80,31,80,30,206,31,255,31,255,30,170,31,231,31,207,31,93,31,160,31,30,31,30,30,242,31,180,31,217,31,228,31,37,31,170,31,238,31,238,30,127,31,58,31,96,31,134,31,62,31,200,31,225,31,76,31,134,31,91,31,189,31,17,31,17,30,207,31,98,31,78,31,136,31,150,31,42,31,60,31,96,31,213,31,31,31,223,31,232,31,37,31,112,31,112,30,112,29,237,31,248,31,187,31,83,31,34,31,159,31,159,30,243,31,197,31,93,31,141,31,141,30,9,31,121,31,82,31,247,31,15,31,35,31,66,31,128,31,128,30,198,31,71,31,182,31,115,31,227,31,164,31,166,31,1,31,154,31,230,31,63,31,53,31,149,31,123,31,184,31,93,31,93,30,215,31,14,31,132,31,206,31,154,31,205,31,239,31,15,31,142,31,212,31,33,31,210,31,229,31,229,30,126,31,126,30,42,31,42,31,186,31,224,31,176,31,176,30,185,31,233,31,127,31,54,31,54,30,206,31,167,31,104,31,94,31,27,31,5,31,243,31,150,31,115,31,206,31,206,30,206,31,174,31,174,30,174,29,203,31,117,31,57,31,85,31,57,31,104,31,222,31,88,31,43,31,43,30,234,31,94,31,125,31,198,31,147,31,147,30,147,29,76,31,76,30,12,31,12,30,12,29,12,28,44,31,156,31,100,31,35,31,180,31,233,31,248,31,114,31,114,30,114,29,114,28,157,31,165,31,202,31,202,30,122,31,64,31,242,31,242,30,242,29,26,31,13,31,221,31,28,31,28,30,28,29,159,31,159,30,213,31,152,31,175,31,199,31,151,31,136,31,28,31,49,31,49,30,234,31,214,31,214,30,42,31,200,31,18,31,18,30,8,31,21,31,6,31,151,31,17,31,253,31,48,31,128,31,128,30,222,31,180,31,84,31,84,30,193,31,193,30,19,31,226,31,101,31,101,30,44,31,48,31,164,31,122,31,223,31,223,30,223,29,71,31,71,30,135,31,56,31,89,31,167,31,167,30,167,29,210,31,158,31,137,31,87,31,38,31,19,31,19,30,214,31,214,30,210,31,184,31,160,31,197,31,185,31,109,31,109,30,238,31,238,30,238,29,208,31,15,31,65,31,139,31,139,30,166,31,122,31,208,31,138,31,103,31,175,31,175,30,96,31,39,31,163,31,195,31,26,31,26,30,180,31,240,31,147,31,147,30,213,31,76,31,51,31,95,31,171,31,171,30,248,31,238,31,117,31,118,31,51,31,18,31,169,31,52,31,164,31,138,31,27,31,190,31,203,31,34,31,34,30,64,31,141,31,81,31,34,31,27,31,134,31,156,31,243,31,109,31,233,31,164,31,67,31,233,31,226,31,6,31,233,31,93,31,183,31,238,31,61,31,153,31,146,31,122,31,223,31,223,30,223,29,121,31,190,31,117,31,123,31,174,31,233,31,176,31,239,31,107,31,3,31,178,31,1,31,1,30,1,29,250,31,213,31,19,31,2,31,189,31,50,31,247,31,104,31,108,31,123,31,153,31,153,30,193,31,171,31,249,31,165,31,108,31,108,30,76,31,239,31,146,31,136,31,113,31,113,30,49,31,49,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
