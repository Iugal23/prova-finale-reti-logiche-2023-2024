-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_382 is
end project_tb_382;

architecture project_tb_arch_382 of project_tb_382 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 930;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,182,0,0,0,118,0,205,0,219,0,224,0,0,0,0,0,101,0,122,0,140,0,212,0,222,0,154,0,15,0,242,0,207,0,29,0,201,0,0,0,98,0,15,0,238,0,124,0,0,0,56,0,223,0,121,0,26,0,2,0,0,0,144,0,131,0,210,0,222,0,172,0,93,0,246,0,114,0,0,0,111,0,0,0,0,0,0,0,136,0,53,0,41,0,120,0,144,0,193,0,244,0,0,0,63,0,154,0,0,0,171,0,122,0,61,0,251,0,168,0,170,0,89,0,130,0,215,0,34,0,247,0,228,0,45,0,0,0,0,0,180,0,105,0,62,0,127,0,149,0,16,0,229,0,15,0,189,0,242,0,68,0,0,0,0,0,250,0,125,0,206,0,0,0,141,0,120,0,62,0,0,0,164,0,14,0,88,0,54,0,154,0,60,0,0,0,125,0,79,0,75,0,113,0,94,0,0,0,44,0,28,0,31,0,238,0,31,0,0,0,70,0,58,0,42,0,21,0,219,0,0,0,39,0,22,0,61,0,209,0,138,0,136,0,248,0,68,0,98,0,8,0,77,0,125,0,94,0,0,0,0,0,83,0,100,0,0,0,0,0,0,0,47,0,102,0,0,0,220,0,0,0,183,0,0,0,46,0,0,0,0,0,252,0,0,0,94,0,0,0,247,0,0,0,0,0,90,0,221,0,100,0,0,0,121,0,174,0,64,0,124,0,31,0,81,0,6,0,194,0,44,0,164,0,0,0,129,0,138,0,170,0,12,0,61,0,241,0,103,0,0,0,27,0,196,0,240,0,138,0,220,0,41,0,45,0,136,0,135,0,136,0,172,0,5,0,204,0,62,0,123,0,243,0,24,0,0,0,0,0,49,0,82,0,208,0,88,0,171,0,69,0,128,0,23,0,0,0,11,0,250,0,0,0,172,0,127,0,0,0,104,0,74,0,107,0,46,0,183,0,83,0,230,0,0,0,169,0,238,0,199,0,0,0,85,0,126,0,0,0,237,0,147,0,160,0,7,0,129,0,197,0,72,0,29,0,192,0,53,0,148,0,53,0,23,0,122,0,0,0,0,0,208,0,52,0,0,0,225,0,183,0,206,0,180,0,82,0,0,0,45,0,0,0,7,0,67,0,163,0,174,0,226,0,0,0,34,0,201,0,95,0,0,0,209,0,0,0,100,0,150,0,0,0,102,0,199,0,0,0,149,0,33,0,72,0,9,0,0,0,242,0,17,0,56,0,120,0,190,0,0,0,74,0,65,0,0,0,138,0,206,0,112,0,232,0,22,0,60,0,179,0,196,0,10,0,95,0,207,0,93,0,197,0,79,0,107,0,177,0,0,0,55,0,0,0,134,0,59,0,0,0,186,0,187,0,0,0,0,0,231,0,208,0,140,0,234,0,102,0,106,0,0,0,0,0,85,0,0,0,206,0,228,0,0,0,0,0,0,0,203,0,119,0,132,0,0,0,0,0,0,0,93,0,95,0,0,0,157,0,241,0,19,0,68,0,8,0,150,0,34,0,0,0,67,0,153,0,2,0,206,0,98,0,215,0,172,0,28,0,6,0,109,0,0,0,236,0,12,0,8,0,219,0,49,0,0,0,74,0,82,0,26,0,71,0,0,0,48,0,15,0,0,0,54,0,231,0,0,0,121,0,174,0,0,0,21,0,76,0,25,0,140,0,207,0,87,0,0,0,120,0,193,0,170,0,22,0,200,0,0,0,0,0,58,0,166,0,137,0,196,0,78,0,248,0,243,0,85,0,66,0,0,0,158,0,99,0,3,0,154,0,70,0,23,0,0,0,183,0,61,0,76,0,0,0,18,0,7,0,64,0,150,0,0,0,53,0,0,0,0,0,95,0,212,0,203,0,203,0,225,0,115,0,0,0,68,0,190,0,254,0,118,0,130,0,160,0,108,0,155,0,1,0,41,0,248,0,48,0,109,0,200,0,209,0,179,0,13,0,183,0,149,0,121,0,240,0,0,0,234,0,19,0,0,0,97,0,66,0,116,0,248,0,146,0,61,0,164,0,180,0,90,0,37,0,48,0,50,0,0,0,0,0,102,0,219,0,123,0,177,0,158,0,0,0,177,0,186,0,0,0,0,0,106,0,85,0,0,0,254,0,42,0,132,0,0,0,165,0,3,0,135,0,114,0,121,0,68,0,136,0,0,0,0,0,205,0,213,0,198,0,242,0,173,0,0,0,236,0,0,0,25,0,170,0,55,0,246,0,1,0,102,0,230,0,130,0,225,0,66,0,211,0,128,0,29,0,146,0,0,0,218,0,208,0,251,0,0,0,247,0,114,0,0,0,224,0,204,0,76,0,33,0,73,0,105,0,180,0,246,0,242,0,223,0,156,0,229,0,55,0,0,0,60,0,0,0,199,0,0,0,0,0,0,0,67,0,83,0,0,0,97,0,154,0,0,0,0,0,8,0,149,0,255,0,212,0,115,0,229,0,0,0,153,0,0,0,112,0,227,0,17,0,67,0,158,0,216,0,33,0,79,0,59,0,250,0,191,0,255,0,202,0,109,0,0,0,192,0,68,0,146,0,0,0,0,0,55,0,184,0,0,0,251,0,190,0,32,0,7,0,110,0,0,0,227,0,0,0,0,0,0,0,89,0,86,0,25,0,178,0,70,0,67,0,0,0,50,0,255,0,0,0,162,0,85,0,74,0,222,0,168,0,247,0,151,0,247,0,33,0,23,0,245,0,77,0,225,0,55,0,227,0,207,0,238,0,0,0,0,0,76,0,86,0,150,0,79,0,11,0,0,0,182,0,23,0,75,0,37,0,71,0,248,0,14,0,224,0,149,0,143,0,101,0,0,0,0,0,59,0,234,0,75,0,239,0,13,0,0,0,140,0,10,0,144,0,93,0,0,0,128,0,244,0,214,0,0,0,68,0,0,0,24,0,232,0,50,0,223,0,0,0,0,0,154,0,213,0,113,0,0,0,234,0,209,0,202,0,0,0,0,0,185,0,196,0,248,0,149,0,107,0,253,0,0,0,0,0,111,0,0,0,0,0,113,0,206,0,44,0,157,0,69,0,12,0,49,0,107,0,100,0,16,0,0,0,4,0,114,0,149,0,204,0,78,0,41,0,67,0,0,0,96,0,4,0,215,0,121,0,18,0,0,0,44,0,82,0,17,0,0,0,56,0,128,0,126,0,147,0,0,0,9,0,132,0,164,0,227,0,0,0,84,0,151,0,31,0,177,0,6,0,196,0,222,0,237,0,173,0,0,0,228,0,78,0,32,0,130,0,131,0,215,0,0,0,130,0,6,0,88,0,0,0,0,0,156,0,0,0,115,0,127,0,200,0,118,0,37,0,0,0,0,0,202,0,200,0,118,0,0,0,78,0,61,0,0,0,211,0,96,0,0,0,0,0,109,0,56,0,238,0,30,0,143,0,38,0,222,0,11,0,0,0,234,0,123,0,116,0,243,0,121,0,84,0,0,0,0,0,15,0,3,0,71,0,149,0,107,0,155,0,199,0,235,0,0,0,24,0,56,0,104,0,2,0,0,0,233,0,98,0,68,0,90,0,0,0,27,0,34,0,103,0,226,0,55,0,0,0,0,0,166,0,38,0,117,0,186,0,26,0,33,0,109,0,87,0,0,0,215,0,56,0,209,0,168,0,40,0,0,0,109,0,0,0,37,0,45,0,0,0,114,0,220,0,192,0,141,0,230,0,236,0,35,0,156,0,157,0,83,0,158,0,89,0,195,0,26,0,115,0,129,0,180,0,73,0,207,0,41,0,45,0,171,0,244,0,237,0,153,0,246,0,128,0,122,0,147,0,195,0,61,0,111,0,206,0,207,0,193,0,0,0,0,0,216,0,0,0,229,0,181,0,207,0,145,0,61,0,146,0,207,0,187,0,0,0,0,0,129,0,75,0,0,0,128,0,40,0,0,0,148,0,220,0,162,0,0,0,218,0,0,0,36,0,180,0,205,0,231,0,166,0,161,0,55,0,81,0,165,0,97,0,248,0,177,0,157,0,129,0,0,0,0,0,251,0,0,0,98,0,242,0,0,0,254,0,34,0,225,0,50,0,0,0,0,0,0,0,219,0,194,0,218,0,139,0,213,0,55,0,219,0,233,0,43,0,209,0,17,0,240,0,90,0,10,0,0,0,164,0,90,0);
signal scenario_full  : scenario_type := (0,0,0,0,182,31,182,30,118,31,205,31,219,31,224,31,224,30,224,29,101,31,122,31,140,31,212,31,222,31,154,31,15,31,242,31,207,31,29,31,201,31,201,30,98,31,15,31,238,31,124,31,124,30,56,31,223,31,121,31,26,31,2,31,2,30,144,31,131,31,210,31,222,31,172,31,93,31,246,31,114,31,114,30,111,31,111,30,111,29,111,28,136,31,53,31,41,31,120,31,144,31,193,31,244,31,244,30,63,31,154,31,154,30,171,31,122,31,61,31,251,31,168,31,170,31,89,31,130,31,215,31,34,31,247,31,228,31,45,31,45,30,45,29,180,31,105,31,62,31,127,31,149,31,16,31,229,31,15,31,189,31,242,31,68,31,68,30,68,29,250,31,125,31,206,31,206,30,141,31,120,31,62,31,62,30,164,31,14,31,88,31,54,31,154,31,60,31,60,30,125,31,79,31,75,31,113,31,94,31,94,30,44,31,28,31,31,31,238,31,31,31,31,30,70,31,58,31,42,31,21,31,219,31,219,30,39,31,22,31,61,31,209,31,138,31,136,31,248,31,68,31,98,31,8,31,77,31,125,31,94,31,94,30,94,29,83,31,100,31,100,30,100,29,100,28,47,31,102,31,102,30,220,31,220,30,183,31,183,30,46,31,46,30,46,29,252,31,252,30,94,31,94,30,247,31,247,30,247,29,90,31,221,31,100,31,100,30,121,31,174,31,64,31,124,31,31,31,81,31,6,31,194,31,44,31,164,31,164,30,129,31,138,31,170,31,12,31,61,31,241,31,103,31,103,30,27,31,196,31,240,31,138,31,220,31,41,31,45,31,136,31,135,31,136,31,172,31,5,31,204,31,62,31,123,31,243,31,24,31,24,30,24,29,49,31,82,31,208,31,88,31,171,31,69,31,128,31,23,31,23,30,11,31,250,31,250,30,172,31,127,31,127,30,104,31,74,31,107,31,46,31,183,31,83,31,230,31,230,30,169,31,238,31,199,31,199,30,85,31,126,31,126,30,237,31,147,31,160,31,7,31,129,31,197,31,72,31,29,31,192,31,53,31,148,31,53,31,23,31,122,31,122,30,122,29,208,31,52,31,52,30,225,31,183,31,206,31,180,31,82,31,82,30,45,31,45,30,7,31,67,31,163,31,174,31,226,31,226,30,34,31,201,31,95,31,95,30,209,31,209,30,100,31,150,31,150,30,102,31,199,31,199,30,149,31,33,31,72,31,9,31,9,30,242,31,17,31,56,31,120,31,190,31,190,30,74,31,65,31,65,30,138,31,206,31,112,31,232,31,22,31,60,31,179,31,196,31,10,31,95,31,207,31,93,31,197,31,79,31,107,31,177,31,177,30,55,31,55,30,134,31,59,31,59,30,186,31,187,31,187,30,187,29,231,31,208,31,140,31,234,31,102,31,106,31,106,30,106,29,85,31,85,30,206,31,228,31,228,30,228,29,228,28,203,31,119,31,132,31,132,30,132,29,132,28,93,31,95,31,95,30,157,31,241,31,19,31,68,31,8,31,150,31,34,31,34,30,67,31,153,31,2,31,206,31,98,31,215,31,172,31,28,31,6,31,109,31,109,30,236,31,12,31,8,31,219,31,49,31,49,30,74,31,82,31,26,31,71,31,71,30,48,31,15,31,15,30,54,31,231,31,231,30,121,31,174,31,174,30,21,31,76,31,25,31,140,31,207,31,87,31,87,30,120,31,193,31,170,31,22,31,200,31,200,30,200,29,58,31,166,31,137,31,196,31,78,31,248,31,243,31,85,31,66,31,66,30,158,31,99,31,3,31,154,31,70,31,23,31,23,30,183,31,61,31,76,31,76,30,18,31,7,31,64,31,150,31,150,30,53,31,53,30,53,29,95,31,212,31,203,31,203,31,225,31,115,31,115,30,68,31,190,31,254,31,118,31,130,31,160,31,108,31,155,31,1,31,41,31,248,31,48,31,109,31,200,31,209,31,179,31,13,31,183,31,149,31,121,31,240,31,240,30,234,31,19,31,19,30,97,31,66,31,116,31,248,31,146,31,61,31,164,31,180,31,90,31,37,31,48,31,50,31,50,30,50,29,102,31,219,31,123,31,177,31,158,31,158,30,177,31,186,31,186,30,186,29,106,31,85,31,85,30,254,31,42,31,132,31,132,30,165,31,3,31,135,31,114,31,121,31,68,31,136,31,136,30,136,29,205,31,213,31,198,31,242,31,173,31,173,30,236,31,236,30,25,31,170,31,55,31,246,31,1,31,102,31,230,31,130,31,225,31,66,31,211,31,128,31,29,31,146,31,146,30,218,31,208,31,251,31,251,30,247,31,114,31,114,30,224,31,204,31,76,31,33,31,73,31,105,31,180,31,246,31,242,31,223,31,156,31,229,31,55,31,55,30,60,31,60,30,199,31,199,30,199,29,199,28,67,31,83,31,83,30,97,31,154,31,154,30,154,29,8,31,149,31,255,31,212,31,115,31,229,31,229,30,153,31,153,30,112,31,227,31,17,31,67,31,158,31,216,31,33,31,79,31,59,31,250,31,191,31,255,31,202,31,109,31,109,30,192,31,68,31,146,31,146,30,146,29,55,31,184,31,184,30,251,31,190,31,32,31,7,31,110,31,110,30,227,31,227,30,227,29,227,28,89,31,86,31,25,31,178,31,70,31,67,31,67,30,50,31,255,31,255,30,162,31,85,31,74,31,222,31,168,31,247,31,151,31,247,31,33,31,23,31,245,31,77,31,225,31,55,31,227,31,207,31,238,31,238,30,238,29,76,31,86,31,150,31,79,31,11,31,11,30,182,31,23,31,75,31,37,31,71,31,248,31,14,31,224,31,149,31,143,31,101,31,101,30,101,29,59,31,234,31,75,31,239,31,13,31,13,30,140,31,10,31,144,31,93,31,93,30,128,31,244,31,214,31,214,30,68,31,68,30,24,31,232,31,50,31,223,31,223,30,223,29,154,31,213,31,113,31,113,30,234,31,209,31,202,31,202,30,202,29,185,31,196,31,248,31,149,31,107,31,253,31,253,30,253,29,111,31,111,30,111,29,113,31,206,31,44,31,157,31,69,31,12,31,49,31,107,31,100,31,16,31,16,30,4,31,114,31,149,31,204,31,78,31,41,31,67,31,67,30,96,31,4,31,215,31,121,31,18,31,18,30,44,31,82,31,17,31,17,30,56,31,128,31,126,31,147,31,147,30,9,31,132,31,164,31,227,31,227,30,84,31,151,31,31,31,177,31,6,31,196,31,222,31,237,31,173,31,173,30,228,31,78,31,32,31,130,31,131,31,215,31,215,30,130,31,6,31,88,31,88,30,88,29,156,31,156,30,115,31,127,31,200,31,118,31,37,31,37,30,37,29,202,31,200,31,118,31,118,30,78,31,61,31,61,30,211,31,96,31,96,30,96,29,109,31,56,31,238,31,30,31,143,31,38,31,222,31,11,31,11,30,234,31,123,31,116,31,243,31,121,31,84,31,84,30,84,29,15,31,3,31,71,31,149,31,107,31,155,31,199,31,235,31,235,30,24,31,56,31,104,31,2,31,2,30,233,31,98,31,68,31,90,31,90,30,27,31,34,31,103,31,226,31,55,31,55,30,55,29,166,31,38,31,117,31,186,31,26,31,33,31,109,31,87,31,87,30,215,31,56,31,209,31,168,31,40,31,40,30,109,31,109,30,37,31,45,31,45,30,114,31,220,31,192,31,141,31,230,31,236,31,35,31,156,31,157,31,83,31,158,31,89,31,195,31,26,31,115,31,129,31,180,31,73,31,207,31,41,31,45,31,171,31,244,31,237,31,153,31,246,31,128,31,122,31,147,31,195,31,61,31,111,31,206,31,207,31,193,31,193,30,193,29,216,31,216,30,229,31,181,31,207,31,145,31,61,31,146,31,207,31,187,31,187,30,187,29,129,31,75,31,75,30,128,31,40,31,40,30,148,31,220,31,162,31,162,30,218,31,218,30,36,31,180,31,205,31,231,31,166,31,161,31,55,31,81,31,165,31,97,31,248,31,177,31,157,31,129,31,129,30,129,29,251,31,251,30,98,31,242,31,242,30,254,31,34,31,225,31,50,31,50,30,50,29,50,28,219,31,194,31,218,31,139,31,213,31,55,31,219,31,233,31,43,31,209,31,17,31,240,31,90,31,10,31,10,30,164,31,90,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
