-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_37 is
end project_tb_37;

architecture project_tb_arch_37 of project_tb_37 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 257;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (154,0,147,0,90,0,209,0,140,0,17,0,188,0,152,0,40,0,138,0,9,0,4,0,0,0,206,0,217,0,83,0,211,0,237,0,170,0,218,0,122,0,80,0,129,0,22,0,0,0,2,0,219,0,98,0,195,0,0,0,0,0,227,0,151,0,253,0,26,0,95,0,85,0,0,0,0,0,156,0,42,0,207,0,0,0,0,0,121,0,133,0,122,0,155,0,194,0,126,0,26,0,0,0,0,0,46,0,129,0,118,0,86,0,0,0,0,0,0,0,243,0,89,0,0,0,225,0,7,0,59,0,249,0,16,0,0,0,169,0,0,0,41,0,252,0,0,0,173,0,113,0,123,0,69,0,115,0,200,0,64,0,17,0,0,0,97,0,175,0,30,0,171,0,0,0,0,0,193,0,142,0,0,0,45,0,68,0,29,0,77,0,90,0,0,0,144,0,0,0,129,0,162,0,0,0,220,0,191,0,99,0,0,0,77,0,254,0,116,0,7,0,91,0,107,0,60,0,107,0,245,0,102,0,141,0,27,0,213,0,198,0,149,0,29,0,59,0,220,0,188,0,64,0,0,0,0,0,125,0,0,0,156,0,195,0,0,0,37,0,0,0,79,0,39,0,109,0,141,0,0,0,0,0,104,0,0,0,167,0,43,0,210,0,57,0,16,0,90,0,9,0,0,0,111,0,93,0,95,0,32,0,97,0,199,0,33,0,0,0,18,0,0,0,255,0,0,0,0,0,0,0,237,0,97,0,139,0,228,0,249,0,207,0,13,0,0,0,0,0,40,0,141,0,188,0,118,0,230,0,107,0,194,0,101,0,81,0,31,0,61,0,249,0,168,0,73,0,97,0,138,0,188,0,238,0,154,0,0,0,252,0,72,0,143,0,143,0,73,0,161,0,201,0,76,0,166,0,85,0,81,0,142,0,232,0,147,0,40,0,249,0,114,0,237,0,162,0,0,0,243,0,150,0,120,0,68,0,83,0,0,0,191,0,118,0,186,0,26,0,187,0,233,0,194,0,83,0,138,0,56,0,0,0,93,0,0,0,246,0,166,0,0,0,0,0,81,0,192,0,0,0,2,0,81,0,152,0,0,0,237,0,184,0,229,0,81,0,121,0,133,0,143,0,227,0,0,0,12,0,143,0,12,0);
signal scenario_full  : scenario_type := (154,31,147,31,90,31,209,31,140,31,17,31,188,31,152,31,40,31,138,31,9,31,4,31,4,30,206,31,217,31,83,31,211,31,237,31,170,31,218,31,122,31,80,31,129,31,22,31,22,30,2,31,219,31,98,31,195,31,195,30,195,29,227,31,151,31,253,31,26,31,95,31,85,31,85,30,85,29,156,31,42,31,207,31,207,30,207,29,121,31,133,31,122,31,155,31,194,31,126,31,26,31,26,30,26,29,46,31,129,31,118,31,86,31,86,30,86,29,86,28,243,31,89,31,89,30,225,31,7,31,59,31,249,31,16,31,16,30,169,31,169,30,41,31,252,31,252,30,173,31,113,31,123,31,69,31,115,31,200,31,64,31,17,31,17,30,97,31,175,31,30,31,171,31,171,30,171,29,193,31,142,31,142,30,45,31,68,31,29,31,77,31,90,31,90,30,144,31,144,30,129,31,162,31,162,30,220,31,191,31,99,31,99,30,77,31,254,31,116,31,7,31,91,31,107,31,60,31,107,31,245,31,102,31,141,31,27,31,213,31,198,31,149,31,29,31,59,31,220,31,188,31,64,31,64,30,64,29,125,31,125,30,156,31,195,31,195,30,37,31,37,30,79,31,39,31,109,31,141,31,141,30,141,29,104,31,104,30,167,31,43,31,210,31,57,31,16,31,90,31,9,31,9,30,111,31,93,31,95,31,32,31,97,31,199,31,33,31,33,30,18,31,18,30,255,31,255,30,255,29,255,28,237,31,97,31,139,31,228,31,249,31,207,31,13,31,13,30,13,29,40,31,141,31,188,31,118,31,230,31,107,31,194,31,101,31,81,31,31,31,61,31,249,31,168,31,73,31,97,31,138,31,188,31,238,31,154,31,154,30,252,31,72,31,143,31,143,31,73,31,161,31,201,31,76,31,166,31,85,31,81,31,142,31,232,31,147,31,40,31,249,31,114,31,237,31,162,31,162,30,243,31,150,31,120,31,68,31,83,31,83,30,191,31,118,31,186,31,26,31,187,31,233,31,194,31,83,31,138,31,56,31,56,30,93,31,93,30,246,31,166,31,166,30,166,29,81,31,192,31,192,30,2,31,81,31,152,31,152,30,237,31,184,31,229,31,81,31,121,31,133,31,143,31,227,31,227,30,12,31,143,31,12,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
