-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 855;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (10,0,237,0,220,0,97,0,234,0,224,0,53,0,0,0,140,0,242,0,251,0,0,0,17,0,0,0,219,0,153,0,13,0,122,0,242,0,0,0,220,0,116,0,23,0,193,0,0,0,45,0,137,0,35,0,242,0,0,0,35,0,209,0,235,0,185,0,242,0,70,0,134,0,142,0,68,0,74,0,4,0,224,0,56,0,58,0,76,0,13,0,56,0,5,0,195,0,0,0,0,0,0,0,0,0,14,0,36,0,217,0,162,0,122,0,137,0,217,0,158,0,222,0,94,0,33,0,0,0,87,0,8,0,236,0,0,0,31,0,68,0,45,0,233,0,178,0,47,0,0,0,186,0,0,0,195,0,225,0,0,0,66,0,66,0,45,0,104,0,80,0,54,0,114,0,252,0,109,0,165,0,0,0,165,0,43,0,205,0,84,0,6,0,168,0,0,0,215,0,27,0,46,0,57,0,133,0,216,0,204,0,176,0,47,0,67,0,50,0,118,0,10,0,196,0,16,0,250,0,16,0,0,0,232,0,0,0,0,0,253,0,0,0,191,0,87,0,0,0,202,0,90,0,18,0,241,0,70,0,115,0,153,0,7,0,0,0,0,0,214,0,48,0,180,0,191,0,45,0,196,0,83,0,224,0,72,0,11,0,0,0,91,0,0,0,152,0,33,0,245,0,173,0,151,0,243,0,177,0,152,0,55,0,59,0,77,0,113,0,87,0,31,0,147,0,153,0,82,0,37,0,11,0,83,0,112,0,0,0,0,0,42,0,159,0,112,0,201,0,0,0,81,0,157,0,223,0,179,0,43,0,0,0,76,0,87,0,172,0,0,0,178,0,0,0,159,0,238,0,79,0,193,0,0,0,120,0,0,0,7,0,0,0,26,0,174,0,115,0,247,0,187,0,188,0,35,0,241,0,171,0,103,0,60,0,206,0,54,0,187,0,0,0,168,0,255,0,39,0,0,0,246,0,0,0,0,0,0,0,162,0,222,0,49,0,68,0,0,0,139,0,0,0,40,0,184,0,0,0,62,0,66,0,215,0,0,0,0,0,206,0,0,0,0,0,229,0,254,0,242,0,132,0,217,0,0,0,242,0,115,0,182,0,96,0,163,0,23,0,155,0,0,0,236,0,0,0,106,0,250,0,174,0,183,0,57,0,192,0,85,0,141,0,69,0,44,0,30,0,23,0,174,0,2,0,0,0,0,0,220,0,237,0,195,0,87,0,163,0,23,0,243,0,0,0,184,0,223,0,155,0,95,0,153,0,82,0,40,0,0,0,106,0,210,0,114,0,97,0,164,0,240,0,0,0,218,0,240,0,83,0,204,0,243,0,91,0,95,0,132,0,45,0,178,0,103,0,37,0,0,0,45,0,87,0,136,0,222,0,155,0,184,0,212,0,0,0,3,0,157,0,225,0,0,0,105,0,0,0,0,0,170,0,198,0,136,0,185,0,211,0,195,0,81,0,90,0,0,0,252,0,27,0,0,0,181,0,189,0,0,0,242,0,206,0,0,0,159,0,0,0,155,0,74,0,135,0,168,0,135,0,208,0,167,0,246,0,115,0,0,0,156,0,196,0,73,0,100,0,236,0,138,0,74,0,92,0,193,0,75,0,87,0,0,0,62,0,248,0,0,0,85,0,7,0,0,0,25,0,174,0,244,0,163,0,229,0,203,0,122,0,214,0,2,0,36,0,19,0,0,0,0,0,17,0,236,0,217,0,188,0,0,0,152,0,255,0,0,0,176,0,0,0,0,0,24,0,91,0,114,0,73,0,222,0,119,0,178,0,121,0,152,0,82,0,166,0,105,0,237,0,63,0,122,0,41,0,0,0,0,0,232,0,79,0,152,0,0,0,205,0,0,0,210,0,223,0,89,0,0,0,233,0,147,0,0,0,147,0,118,0,0,0,190,0,93,0,39,0,201,0,0,0,181,0,23,0,13,0,162,0,95,0,0,0,140,0,197,0,0,0,50,0,76,0,4,0,168,0,154,0,0,0,16,0,178,0,102,0,208,0,0,0,246,0,36,0,169,0,0,0,169,0,117,0,162,0,48,0,171,0,122,0,13,0,177,0,88,0,0,0,201,0,222,0,221,0,148,0,108,0,193,0,17,0,249,0,5,0,18,0,198,0,84,0,119,0,79,0,245,0,177,0,10,0,0,0,157,0,118,0,234,0,55,0,0,0,5,0,0,0,0,0,123,0,15,0,0,0,119,0,28,0,139,0,231,0,31,0,241,0,246,0,214,0,250,0,0,0,106,0,45,0,8,0,0,0,33,0,219,0,209,0,209,0,155,0,0,0,151,0,39,0,48,0,102,0,85,0,164,0,252,0,16,0,0,0,213,0,125,0,174,0,109,0,173,0,94,0,0,0,193,0,177,0,114,0,0,0,0,0,197,0,209,0,0,0,23,0,249,0,0,0,111,0,150,0,139,0,91,0,247,0,0,0,18,0,232,0,158,0,203,0,152,0,179,0,0,0,1,0,0,0,145,0,159,0,0,0,189,0,89,0,201,0,0,0,123,0,118,0,76,0,146,0,120,0,0,0,0,0,52,0,162,0,206,0,40,0,0,0,21,0,77,0,0,0,209,0,78,0,0,0,141,0,196,0,65,0,0,0,0,0,250,0,215,0,89,0,238,0,223,0,235,0,201,0,211,0,207,0,215,0,0,0,0,0,197,0,0,0,160,0,0,0,195,0,229,0,176,0,30,0,244,0,23,0,154,0,221,0,238,0,26,0,110,0,62,0,66,0,0,0,129,0,117,0,234,0,252,0,0,0,58,0,86,0,39,0,45,0,207,0,0,0,41,0,1,0,0,0,188,0,0,0,38,0,113,0,218,0,89,0,168,0,127,0,180,0,58,0,19,0,0,0,38,0,131,0,35,0,2,0,0,0,29,0,167,0,0,0,197,0,7,0,165,0,6,0,53,0,0,0,179,0,115,0,3,0,105,0,202,0,0,0,93,0,0,0,5,0,0,0,75,0,130,0,25,0,74,0,245,0,213,0,0,0,201,0,168,0,0,0,0,0,214,0,189,0,208,0,147,0,108,0,74,0,77,0,167,0,95,0,165,0,110,0,176,0,104,0,78,0,161,0,101,0,24,0,189,0,222,0,0,0,125,0,0,0,0,0,13,0,0,0,201,0,164,0,0,0,0,0,72,0,77,0,41,0,0,0,170,0,200,0,222,0,155,0,236,0,0,0,199,0,211,0,84,0,58,0,245,0,0,0,4,0,192,0,138,0,93,0,247,0,251,0,165,0,16,0,127,0,77,0,246,0,151,0,107,0,148,0,130,0,0,0,167,0,47,0,78,0,99,0,13,0,0,0,53,0,46,0,37,0,0,0,0,0,183,0,176,0,102,0,78,0,250,0,21,0,0,0,201,0,157,0,125,0,0,0,62,0,0,0,13,0,152,0,0,0,86,0,184,0,79,0,253,0,0,0,187,0,46,0,20,0,0,0,228,0,166,0,186,0,98,0,111,0,173,0,210,0,0,0,0,0,169,0,0,0,36,0,12,0,17,0,107,0,210,0,52,0,187,0,246,0,195,0,81,0,192,0,24,0,87,0,122,0,0,0,66,0,141,0,0,0,255,0,0,0,234,0,0,0,84,0,118,0,209,0,168,0,77,0,148,0,142,0,214,0,127,0,0,0,0,0,0,0,0,0,128,0,1,0,73,0,0,0,218,0,162,0,177,0,34,0,0,0,227,0,60,0,10,0,117,0,72,0,227,0,115,0,187,0,230,0,196,0,0,0,0,0,240,0,217,0,44,0,171,0,0,0,150,0,28,0,0,0,180,0,226,0,213,0,213,0,126,0);
signal scenario_full  : scenario_type := (10,31,237,31,220,31,97,31,234,31,224,31,53,31,53,30,140,31,242,31,251,31,251,30,17,31,17,30,219,31,153,31,13,31,122,31,242,31,242,30,220,31,116,31,23,31,193,31,193,30,45,31,137,31,35,31,242,31,242,30,35,31,209,31,235,31,185,31,242,31,70,31,134,31,142,31,68,31,74,31,4,31,224,31,56,31,58,31,76,31,13,31,56,31,5,31,195,31,195,30,195,29,195,28,195,27,14,31,36,31,217,31,162,31,122,31,137,31,217,31,158,31,222,31,94,31,33,31,33,30,87,31,8,31,236,31,236,30,31,31,68,31,45,31,233,31,178,31,47,31,47,30,186,31,186,30,195,31,225,31,225,30,66,31,66,31,45,31,104,31,80,31,54,31,114,31,252,31,109,31,165,31,165,30,165,31,43,31,205,31,84,31,6,31,168,31,168,30,215,31,27,31,46,31,57,31,133,31,216,31,204,31,176,31,47,31,67,31,50,31,118,31,10,31,196,31,16,31,250,31,16,31,16,30,232,31,232,30,232,29,253,31,253,30,191,31,87,31,87,30,202,31,90,31,18,31,241,31,70,31,115,31,153,31,7,31,7,30,7,29,214,31,48,31,180,31,191,31,45,31,196,31,83,31,224,31,72,31,11,31,11,30,91,31,91,30,152,31,33,31,245,31,173,31,151,31,243,31,177,31,152,31,55,31,59,31,77,31,113,31,87,31,31,31,147,31,153,31,82,31,37,31,11,31,83,31,112,31,112,30,112,29,42,31,159,31,112,31,201,31,201,30,81,31,157,31,223,31,179,31,43,31,43,30,76,31,87,31,172,31,172,30,178,31,178,30,159,31,238,31,79,31,193,31,193,30,120,31,120,30,7,31,7,30,26,31,174,31,115,31,247,31,187,31,188,31,35,31,241,31,171,31,103,31,60,31,206,31,54,31,187,31,187,30,168,31,255,31,39,31,39,30,246,31,246,30,246,29,246,28,162,31,222,31,49,31,68,31,68,30,139,31,139,30,40,31,184,31,184,30,62,31,66,31,215,31,215,30,215,29,206,31,206,30,206,29,229,31,254,31,242,31,132,31,217,31,217,30,242,31,115,31,182,31,96,31,163,31,23,31,155,31,155,30,236,31,236,30,106,31,250,31,174,31,183,31,57,31,192,31,85,31,141,31,69,31,44,31,30,31,23,31,174,31,2,31,2,30,2,29,220,31,237,31,195,31,87,31,163,31,23,31,243,31,243,30,184,31,223,31,155,31,95,31,153,31,82,31,40,31,40,30,106,31,210,31,114,31,97,31,164,31,240,31,240,30,218,31,240,31,83,31,204,31,243,31,91,31,95,31,132,31,45,31,178,31,103,31,37,31,37,30,45,31,87,31,136,31,222,31,155,31,184,31,212,31,212,30,3,31,157,31,225,31,225,30,105,31,105,30,105,29,170,31,198,31,136,31,185,31,211,31,195,31,81,31,90,31,90,30,252,31,27,31,27,30,181,31,189,31,189,30,242,31,206,31,206,30,159,31,159,30,155,31,74,31,135,31,168,31,135,31,208,31,167,31,246,31,115,31,115,30,156,31,196,31,73,31,100,31,236,31,138,31,74,31,92,31,193,31,75,31,87,31,87,30,62,31,248,31,248,30,85,31,7,31,7,30,25,31,174,31,244,31,163,31,229,31,203,31,122,31,214,31,2,31,36,31,19,31,19,30,19,29,17,31,236,31,217,31,188,31,188,30,152,31,255,31,255,30,176,31,176,30,176,29,24,31,91,31,114,31,73,31,222,31,119,31,178,31,121,31,152,31,82,31,166,31,105,31,237,31,63,31,122,31,41,31,41,30,41,29,232,31,79,31,152,31,152,30,205,31,205,30,210,31,223,31,89,31,89,30,233,31,147,31,147,30,147,31,118,31,118,30,190,31,93,31,39,31,201,31,201,30,181,31,23,31,13,31,162,31,95,31,95,30,140,31,197,31,197,30,50,31,76,31,4,31,168,31,154,31,154,30,16,31,178,31,102,31,208,31,208,30,246,31,36,31,169,31,169,30,169,31,117,31,162,31,48,31,171,31,122,31,13,31,177,31,88,31,88,30,201,31,222,31,221,31,148,31,108,31,193,31,17,31,249,31,5,31,18,31,198,31,84,31,119,31,79,31,245,31,177,31,10,31,10,30,157,31,118,31,234,31,55,31,55,30,5,31,5,30,5,29,123,31,15,31,15,30,119,31,28,31,139,31,231,31,31,31,241,31,246,31,214,31,250,31,250,30,106,31,45,31,8,31,8,30,33,31,219,31,209,31,209,31,155,31,155,30,151,31,39,31,48,31,102,31,85,31,164,31,252,31,16,31,16,30,213,31,125,31,174,31,109,31,173,31,94,31,94,30,193,31,177,31,114,31,114,30,114,29,197,31,209,31,209,30,23,31,249,31,249,30,111,31,150,31,139,31,91,31,247,31,247,30,18,31,232,31,158,31,203,31,152,31,179,31,179,30,1,31,1,30,145,31,159,31,159,30,189,31,89,31,201,31,201,30,123,31,118,31,76,31,146,31,120,31,120,30,120,29,52,31,162,31,206,31,40,31,40,30,21,31,77,31,77,30,209,31,78,31,78,30,141,31,196,31,65,31,65,30,65,29,250,31,215,31,89,31,238,31,223,31,235,31,201,31,211,31,207,31,215,31,215,30,215,29,197,31,197,30,160,31,160,30,195,31,229,31,176,31,30,31,244,31,23,31,154,31,221,31,238,31,26,31,110,31,62,31,66,31,66,30,129,31,117,31,234,31,252,31,252,30,58,31,86,31,39,31,45,31,207,31,207,30,41,31,1,31,1,30,188,31,188,30,38,31,113,31,218,31,89,31,168,31,127,31,180,31,58,31,19,31,19,30,38,31,131,31,35,31,2,31,2,30,29,31,167,31,167,30,197,31,7,31,165,31,6,31,53,31,53,30,179,31,115,31,3,31,105,31,202,31,202,30,93,31,93,30,5,31,5,30,75,31,130,31,25,31,74,31,245,31,213,31,213,30,201,31,168,31,168,30,168,29,214,31,189,31,208,31,147,31,108,31,74,31,77,31,167,31,95,31,165,31,110,31,176,31,104,31,78,31,161,31,101,31,24,31,189,31,222,31,222,30,125,31,125,30,125,29,13,31,13,30,201,31,164,31,164,30,164,29,72,31,77,31,41,31,41,30,170,31,200,31,222,31,155,31,236,31,236,30,199,31,211,31,84,31,58,31,245,31,245,30,4,31,192,31,138,31,93,31,247,31,251,31,165,31,16,31,127,31,77,31,246,31,151,31,107,31,148,31,130,31,130,30,167,31,47,31,78,31,99,31,13,31,13,30,53,31,46,31,37,31,37,30,37,29,183,31,176,31,102,31,78,31,250,31,21,31,21,30,201,31,157,31,125,31,125,30,62,31,62,30,13,31,152,31,152,30,86,31,184,31,79,31,253,31,253,30,187,31,46,31,20,31,20,30,228,31,166,31,186,31,98,31,111,31,173,31,210,31,210,30,210,29,169,31,169,30,36,31,12,31,17,31,107,31,210,31,52,31,187,31,246,31,195,31,81,31,192,31,24,31,87,31,122,31,122,30,66,31,141,31,141,30,255,31,255,30,234,31,234,30,84,31,118,31,209,31,168,31,77,31,148,31,142,31,214,31,127,31,127,30,127,29,127,28,127,27,128,31,1,31,73,31,73,30,218,31,162,31,177,31,34,31,34,30,227,31,60,31,10,31,117,31,72,31,227,31,115,31,187,31,230,31,196,31,196,30,196,29,240,31,217,31,44,31,171,31,171,30,150,31,28,31,28,30,180,31,226,31,213,31,213,31,126,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
