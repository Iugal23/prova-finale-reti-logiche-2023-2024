-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_477 is
end project_tb_477;

architecture project_tb_arch_477 of project_tb_477 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 524;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (218,0,67,0,0,0,243,0,38,0,0,0,0,0,66,0,213,0,148,0,228,0,0,0,158,0,152,0,222,0,0,0,21,0,234,0,0,0,36,0,105,0,140,0,110,0,45,0,0,0,76,0,69,0,194,0,31,0,114,0,252,0,17,0,127,0,0,0,132,0,0,0,0,0,0,0,204,0,126,0,80,0,178,0,0,0,15,0,176,0,240,0,25,0,15,0,47,0,0,0,0,0,76,0,114,0,229,0,0,0,174,0,0,0,0,0,226,0,0,0,217,0,210,0,0,0,210,0,240,0,0,0,22,0,57,0,138,0,219,0,0,0,36,0,67,0,0,0,7,0,107,0,108,0,0,0,204,0,237,0,111,0,0,0,0,0,0,0,143,0,38,0,172,0,213,0,7,0,117,0,56,0,115,0,0,0,128,0,0,0,202,0,0,0,69,0,13,0,0,0,226,0,166,0,166,0,214,0,0,0,165,0,183,0,0,0,207,0,245,0,0,0,194,0,91,0,36,0,0,0,100,0,143,0,0,0,57,0,0,0,35,0,104,0,37,0,7,0,20,0,12,0,89,0,0,0,22,0,231,0,0,0,36,0,42,0,95,0,11,0,0,0,170,0,0,0,189,0,155,0,0,0,0,0,0,0,137,0,223,0,173,0,27,0,224,0,231,0,140,0,221,0,0,0,0,0,0,0,19,0,51,0,210,0,0,0,135,0,0,0,0,0,164,0,21,0,217,0,126,0,120,0,159,0,128,0,0,0,201,0,67,0,0,0,0,0,0,0,37,0,58,0,0,0,234,0,37,0,95,0,178,0,116,0,228,0,0,0,179,0,2,0,184,0,0,0,48,0,145,0,44,0,253,0,86,0,184,0,156,0,135,0,210,0,50,0,0,0,43,0,137,0,0,0,43,0,64,0,69,0,171,0,224,0,0,0,33,0,250,0,16,0,207,0,28,0,244,0,0,0,101,0,13,0,11,0,217,0,196,0,89,0,115,0,0,0,0,0,174,0,0,0,216,0,29,0,177,0,0,0,129,0,0,0,0,0,141,0,233,0,21,0,16,0,47,0,116,0,66,0,49,0,0,0,47,0,6,0,137,0,147,0,109,0,204,0,0,0,157,0,0,0,55,0,94,0,0,0,225,0,14,0,0,0,0,0,201,0,35,0,210,0,149,0,255,0,155,0,45,0,113,0,89,0,73,0,6,0,154,0,0,0,58,0,250,0,226,0,83,0,152,0,211,0,113,0,110,0,213,0,79,0,202,0,0,0,0,0,0,0,50,0,180,0,104,0,171,0,0,0,166,0,157,0,0,0,50,0,209,0,0,0,0,0,11,0,143,0,197,0,0,0,0,0,229,0,175,0,0,0,0,0,232,0,37,0,0,0,0,0,4,0,120,0,66,0,233,0,103,0,43,0,66,0,0,0,13,0,184,0,145,0,0,0,35,0,241,0,0,0,53,0,211,0,148,0,179,0,248,0,0,0,122,0,0,0,219,0,180,0,154,0,103,0,117,0,11,0,0,0,200,0,159,0,166,0,86,0,45,0,219,0,139,0,175,0,220,0,96,0,0,0,35,0,154,0,236,0,146,0,20,0,93,0,6,0,0,0,0,0,178,0,99,0,0,0,116,0,130,0,0,0,222,0,163,0,185,0,0,0,54,0,0,0,0,0,71,0,166,0,126,0,0,0,0,0,144,0,215,0,16,0,190,0,93,0,63,0,0,0,210,0,149,0,0,0,5,0,0,0,142,0,21,0,117,0,107,0,247,0,59,0,112,0,134,0,0,0,111,0,195,0,0,0,16,0,119,0,148,0,240,0,133,0,0,0,0,0,254,0,160,0,53,0,0,0,160,0,0,0,182,0,32,0,93,0,151,0,223,0,44,0,230,0,173,0,26,0,11,0,82,0,130,0,7,0,208,0,217,0,249,0,250,0,0,0,5,0,0,0,229,0,108,0,0,0,178,0,125,0,49,0,143,0,15,0,0,0,57,0,0,0,58,0,166,0,63,0,0,0,140,0,6,0,181,0,215,0,0,0,126,0,8,0,46,0,246,0,183,0,0,0,46,0,63,0,174,0,89,0,241,0,170,0,104,0,70,0,166,0,56,0,25,0,90,0,106,0,168,0,62,0,203,0,62,0,113,0,228,0,204,0,173,0,0,0,166,0,0,0,62,0,0,0,21,0,12,0,99,0,192,0,205,0,243,0,0,0,199,0,0,0,246,0,118,0,118,0,0,0,231,0,30,0,0,0,200,0,0,0,0,0,253,0,27,0,250,0,183,0,119,0,31,0,0,0,235,0,0,0,97,0,0,0,90,0,9,0,91,0,111,0,127,0,0,0,0,0);
signal scenario_full  : scenario_type := (218,31,67,31,67,30,243,31,38,31,38,30,38,29,66,31,213,31,148,31,228,31,228,30,158,31,152,31,222,31,222,30,21,31,234,31,234,30,36,31,105,31,140,31,110,31,45,31,45,30,76,31,69,31,194,31,31,31,114,31,252,31,17,31,127,31,127,30,132,31,132,30,132,29,132,28,204,31,126,31,80,31,178,31,178,30,15,31,176,31,240,31,25,31,15,31,47,31,47,30,47,29,76,31,114,31,229,31,229,30,174,31,174,30,174,29,226,31,226,30,217,31,210,31,210,30,210,31,240,31,240,30,22,31,57,31,138,31,219,31,219,30,36,31,67,31,67,30,7,31,107,31,108,31,108,30,204,31,237,31,111,31,111,30,111,29,111,28,143,31,38,31,172,31,213,31,7,31,117,31,56,31,115,31,115,30,128,31,128,30,202,31,202,30,69,31,13,31,13,30,226,31,166,31,166,31,214,31,214,30,165,31,183,31,183,30,207,31,245,31,245,30,194,31,91,31,36,31,36,30,100,31,143,31,143,30,57,31,57,30,35,31,104,31,37,31,7,31,20,31,12,31,89,31,89,30,22,31,231,31,231,30,36,31,42,31,95,31,11,31,11,30,170,31,170,30,189,31,155,31,155,30,155,29,155,28,137,31,223,31,173,31,27,31,224,31,231,31,140,31,221,31,221,30,221,29,221,28,19,31,51,31,210,31,210,30,135,31,135,30,135,29,164,31,21,31,217,31,126,31,120,31,159,31,128,31,128,30,201,31,67,31,67,30,67,29,67,28,37,31,58,31,58,30,234,31,37,31,95,31,178,31,116,31,228,31,228,30,179,31,2,31,184,31,184,30,48,31,145,31,44,31,253,31,86,31,184,31,156,31,135,31,210,31,50,31,50,30,43,31,137,31,137,30,43,31,64,31,69,31,171,31,224,31,224,30,33,31,250,31,16,31,207,31,28,31,244,31,244,30,101,31,13,31,11,31,217,31,196,31,89,31,115,31,115,30,115,29,174,31,174,30,216,31,29,31,177,31,177,30,129,31,129,30,129,29,141,31,233,31,21,31,16,31,47,31,116,31,66,31,49,31,49,30,47,31,6,31,137,31,147,31,109,31,204,31,204,30,157,31,157,30,55,31,94,31,94,30,225,31,14,31,14,30,14,29,201,31,35,31,210,31,149,31,255,31,155,31,45,31,113,31,89,31,73,31,6,31,154,31,154,30,58,31,250,31,226,31,83,31,152,31,211,31,113,31,110,31,213,31,79,31,202,31,202,30,202,29,202,28,50,31,180,31,104,31,171,31,171,30,166,31,157,31,157,30,50,31,209,31,209,30,209,29,11,31,143,31,197,31,197,30,197,29,229,31,175,31,175,30,175,29,232,31,37,31,37,30,37,29,4,31,120,31,66,31,233,31,103,31,43,31,66,31,66,30,13,31,184,31,145,31,145,30,35,31,241,31,241,30,53,31,211,31,148,31,179,31,248,31,248,30,122,31,122,30,219,31,180,31,154,31,103,31,117,31,11,31,11,30,200,31,159,31,166,31,86,31,45,31,219,31,139,31,175,31,220,31,96,31,96,30,35,31,154,31,236,31,146,31,20,31,93,31,6,31,6,30,6,29,178,31,99,31,99,30,116,31,130,31,130,30,222,31,163,31,185,31,185,30,54,31,54,30,54,29,71,31,166,31,126,31,126,30,126,29,144,31,215,31,16,31,190,31,93,31,63,31,63,30,210,31,149,31,149,30,5,31,5,30,142,31,21,31,117,31,107,31,247,31,59,31,112,31,134,31,134,30,111,31,195,31,195,30,16,31,119,31,148,31,240,31,133,31,133,30,133,29,254,31,160,31,53,31,53,30,160,31,160,30,182,31,32,31,93,31,151,31,223,31,44,31,230,31,173,31,26,31,11,31,82,31,130,31,7,31,208,31,217,31,249,31,250,31,250,30,5,31,5,30,229,31,108,31,108,30,178,31,125,31,49,31,143,31,15,31,15,30,57,31,57,30,58,31,166,31,63,31,63,30,140,31,6,31,181,31,215,31,215,30,126,31,8,31,46,31,246,31,183,31,183,30,46,31,63,31,174,31,89,31,241,31,170,31,104,31,70,31,166,31,56,31,25,31,90,31,106,31,168,31,62,31,203,31,62,31,113,31,228,31,204,31,173,31,173,30,166,31,166,30,62,31,62,30,21,31,12,31,99,31,192,31,205,31,243,31,243,30,199,31,199,30,246,31,118,31,118,31,118,30,231,31,30,31,30,30,200,31,200,30,200,29,253,31,27,31,250,31,183,31,119,31,31,31,31,30,235,31,235,30,97,31,97,30,90,31,9,31,91,31,111,31,127,31,127,30,127,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
