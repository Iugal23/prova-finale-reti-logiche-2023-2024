-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_5 is
end project_tb_5;

architecture project_tb_arch_5 of project_tb_5 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 905;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (35,0,148,0,65,0,246,0,151,0,89,0,51,0,0,0,3,0,18,0,76,0,172,0,0,0,103,0,206,0,77,0,148,0,6,0,145,0,196,0,117,0,49,0,0,0,233,0,0,0,96,0,55,0,0,0,130,0,189,0,0,0,0,0,219,0,194,0,0,0,170,0,0,0,0,0,0,0,200,0,222,0,0,0,64,0,0,0,160,0,12,0,109,0,42,0,0,0,212,0,197,0,8,0,0,0,17,0,35,0,89,0,98,0,132,0,194,0,0,0,27,0,11,0,0,0,0,0,2,0,108,0,240,0,82,0,93,0,0,0,214,0,105,0,229,0,156,0,127,0,200,0,59,0,109,0,173,0,0,0,64,0,92,0,226,0,0,0,0,0,71,0,154,0,67,0,96,0,47,0,13,0,0,0,0,0,8,0,47,0,236,0,3,0,0,0,129,0,0,0,107,0,195,0,75,0,187,0,203,0,238,0,190,0,0,0,0,0,0,0,0,0,0,0,66,0,8,0,0,0,185,0,0,0,166,0,114,0,42,0,224,0,1,0,0,0,119,0,249,0,120,0,250,0,201,0,3,0,0,0,30,0,0,0,32,0,75,0,24,0,98,0,37,0,203,0,11,0,25,0,136,0,0,0,251,0,242,0,224,0,11,0,44,0,164,0,46,0,0,0,170,0,0,0,117,0,168,0,207,0,31,0,0,0,212,0,99,0,195,0,0,0,79,0,43,0,231,0,0,0,210,0,132,0,177,0,68,0,205,0,198,0,114,0,94,0,0,0,38,0,0,0,251,0,216,0,80,0,188,0,22,0,241,0,0,0,45,0,184,0,0,0,98,0,191,0,0,0,166,0,119,0,0,0,0,0,32,0,134,0,224,0,193,0,0,0,124,0,6,0,164,0,146,0,251,0,117,0,115,0,87,0,162,0,171,0,152,0,224,0,185,0,0,0,81,0,23,0,111,0,25,0,0,0,11,0,8,0,81,0,187,0,24,0,27,0,132,0,73,0,0,0,120,0,250,0,0,0,81,0,42,0,0,0,220,0,253,0,198,0,202,0,42,0,42,0,47,0,113,0,93,0,0,0,0,0,0,0,179,0,0,0,0,0,62,0,156,0,0,0,129,0,95,0,250,0,0,0,87,0,148,0,12,0,0,0,160,0,8,0,217,0,100,0,130,0,39,0,91,0,117,0,4,0,81,0,0,0,153,0,13,0,78,0,162,0,32,0,61,0,172,0,197,0,57,0,183,0,44,0,35,0,222,0,243,0,28,0,113,0,238,0,192,0,64,0,42,0,61,0,143,0,0,0,144,0,51,0,233,0,16,0,246,0,77,0,0,0,46,0,238,0,21,0,132,0,0,0,34,0,82,0,48,0,252,0,0,0,0,0,0,0,153,0,156,0,6,0,61,0,83,0,157,0,0,0,126,0,184,0,100,0,34,0,27,0,0,0,0,0,179,0,0,0,171,0,112,0,152,0,0,0,46,0,151,0,132,0,0,0,195,0,2,0,161,0,12,0,212,0,251,0,146,0,255,0,0,0,25,0,0,0,28,0,0,0,107,0,0,0,0,0,0,0,189,0,235,0,0,0,40,0,65,0,0,0,117,0,25,0,65,0,252,0,52,0,7,0,0,0,0,0,109,0,175,0,220,0,120,0,239,0,171,0,248,0,124,0,0,0,132,0,242,0,112,0,118,0,95,0,181,0,24,0,169,0,184,0,165,0,24,0,93,0,225,0,116,0,145,0,155,0,39,0,86,0,49,0,133,0,31,0,11,0,195,0,0,0,28,0,144,0,0,0,0,0,75,0,96,0,147,0,196,0,99,0,0,0,141,0,35,0,129,0,0,0,241,0,26,0,186,0,0,0,0,0,223,0,249,0,112,0,0,0,0,0,147,0,0,0,9,0,93,0,230,0,170,0,84,0,206,0,8,0,216,0,147,0,147,0,199,0,76,0,54,0,73,0,223,0,0,0,190,0,0,0,97,0,173,0,239,0,169,0,204,0,178,0,0,0,202,0,221,0,43,0,97,0,0,0,0,0,126,0,192,0,1,0,0,0,44,0,238,0,0,0,220,0,0,0,26,0,0,0,2,0,143,0,52,0,0,0,157,0,0,0,239,0,189,0,147,0,0,0,0,0,0,0,252,0,0,0,199,0,187,0,0,0,236,0,105,0,251,0,234,0,172,0,0,0,189,0,0,0,60,0,0,0,170,0,0,0,211,0,113,0,240,0,82,0,186,0,191,0,48,0,41,0,0,0,15,0,132,0,248,0,221,0,116,0,0,0,0,0,75,0,201,0,35,0,94,0,0,0,115,0,102,0,0,0,244,0,82,0,171,0,172,0,13,0,135,0,82,0,0,0,215,0,0,0,0,0,0,0,230,0,201,0,34,0,11,0,12,0,204,0,65,0,157,0,114,0,6,0,159,0,17,0,42,0,241,0,80,0,0,0,241,0,233,0,12,0,40,0,183,0,145,0,62,0,168,0,81,0,0,0,0,0,180,0,208,0,242,0,25,0,0,0,214,0,0,0,75,0,0,0,165,0,251,0,21,0,189,0,215,0,78,0,208,0,208,0,72,0,179,0,31,0,239,0,0,0,111,0,241,0,128,0,172,0,41,0,249,0,63,0,0,0,198,0,203,0,171,0,153,0,61,0,49,0,26,0,206,0,0,0,235,0,108,0,154,0,245,0,104,0,19,0,255,0,118,0,2,0,211,0,201,0,0,0,0,0,118,0,79,0,200,0,43,0,0,0,0,0,111,0,183,0,191,0,149,0,0,0,124,0,0,0,170,0,89,0,161,0,125,0,4,0,0,0,219,0,185,0,240,0,0,0,197,0,0,0,231,0,214,0,0,0,0,0,183,0,124,0,61,0,69,0,246,0,139,0,156,0,123,0,0,0,60,0,150,0,135,0,0,0,153,0,0,0,228,0,137,0,197,0,40,0,0,0,0,0,210,0,93,0,222,0,183,0,0,0,177,0,215,0,7,0,9,0,0,0,125,0,21,0,124,0,251,0,42,0,51,0,204,0,23,0,156,0,117,0,238,0,0,0,228,0,0,0,101,0,0,0,102,0,29,0,218,0,122,0,195,0,185,0,71,0,103,0,208,0,61,0,238,0,134,0,252,0,0,0,0,0,27,0,59,0,149,0,162,0,208,0,78,0,0,0,0,0,172,0,198,0,33,0,84,0,151,0,0,0,203,0,220,0,53,0,101,0,153,0,160,0,99,0,96,0,0,0,248,0,16,0,199,0,0,0,0,0,122,0,80,0,60,0,205,0,186,0,96,0,68,0,7,0,29,0,236,0,235,0,1,0,0,0,0,0,215,0,44,0,0,0,0,0,18,0,0,0,75,0,205,0,240,0,78,0,59,0,31,0,67,0,78,0,210,0,162,0,249,0,135,0,133,0,107,0,118,0,3,0,84,0,0,0,33,0,0,0,62,0,229,0,28,0,54,0,103,0,66,0,0,0,29,0,211,0,44,0,215,0,46,0,173,0,0,0,0,0,124,0,133,0,0,0,246,0,0,0,0,0,136,0,165,0,0,0,119,0,54,0,7,0,75,0,209,0,213,0,69,0,20,0,54,0,0,0,4,0,0,0,31,0,44,0,0,0,1,0,16,0,138,0,34,0,162,0,0,0,246,0,104,0,89,0,237,0,0,0,21,0,0,0,0,0,184,0,0,0,129,0,0,0,127,0,142,0,150,0,72,0,105,0,77,0,23,0,51,0,0,0,0,0,0,0,56,0,189,0,171,0,175,0,207,0,0,0,232,0,94,0,188,0,138,0,207,0,237,0,125,0,87,0,0,0,0,0,87,0,50,0,230,0,66,0,137,0,0,0,46,0,140,0,0,0,0,0,24,0,247,0,139,0,27,0,15,0,47,0,124,0,241,0,34,0,240,0,146,0,174,0,97,0,158,0,153,0,243,0,228,0,123,0,199,0,165,0,98,0,0,0,95,0,238,0,0,0,248,0,85,0,91,0,119,0,205,0,184,0,0,0,28,0,250,0,19,0,0,0,111,0,173,0,0,0,174,0,38,0);
signal scenario_full  : scenario_type := (35,31,148,31,65,31,246,31,151,31,89,31,51,31,51,30,3,31,18,31,76,31,172,31,172,30,103,31,206,31,77,31,148,31,6,31,145,31,196,31,117,31,49,31,49,30,233,31,233,30,96,31,55,31,55,30,130,31,189,31,189,30,189,29,219,31,194,31,194,30,170,31,170,30,170,29,170,28,200,31,222,31,222,30,64,31,64,30,160,31,12,31,109,31,42,31,42,30,212,31,197,31,8,31,8,30,17,31,35,31,89,31,98,31,132,31,194,31,194,30,27,31,11,31,11,30,11,29,2,31,108,31,240,31,82,31,93,31,93,30,214,31,105,31,229,31,156,31,127,31,200,31,59,31,109,31,173,31,173,30,64,31,92,31,226,31,226,30,226,29,71,31,154,31,67,31,96,31,47,31,13,31,13,30,13,29,8,31,47,31,236,31,3,31,3,30,129,31,129,30,107,31,195,31,75,31,187,31,203,31,238,31,190,31,190,30,190,29,190,28,190,27,190,26,66,31,8,31,8,30,185,31,185,30,166,31,114,31,42,31,224,31,1,31,1,30,119,31,249,31,120,31,250,31,201,31,3,31,3,30,30,31,30,30,32,31,75,31,24,31,98,31,37,31,203,31,11,31,25,31,136,31,136,30,251,31,242,31,224,31,11,31,44,31,164,31,46,31,46,30,170,31,170,30,117,31,168,31,207,31,31,31,31,30,212,31,99,31,195,31,195,30,79,31,43,31,231,31,231,30,210,31,132,31,177,31,68,31,205,31,198,31,114,31,94,31,94,30,38,31,38,30,251,31,216,31,80,31,188,31,22,31,241,31,241,30,45,31,184,31,184,30,98,31,191,31,191,30,166,31,119,31,119,30,119,29,32,31,134,31,224,31,193,31,193,30,124,31,6,31,164,31,146,31,251,31,117,31,115,31,87,31,162,31,171,31,152,31,224,31,185,31,185,30,81,31,23,31,111,31,25,31,25,30,11,31,8,31,81,31,187,31,24,31,27,31,132,31,73,31,73,30,120,31,250,31,250,30,81,31,42,31,42,30,220,31,253,31,198,31,202,31,42,31,42,31,47,31,113,31,93,31,93,30,93,29,93,28,179,31,179,30,179,29,62,31,156,31,156,30,129,31,95,31,250,31,250,30,87,31,148,31,12,31,12,30,160,31,8,31,217,31,100,31,130,31,39,31,91,31,117,31,4,31,81,31,81,30,153,31,13,31,78,31,162,31,32,31,61,31,172,31,197,31,57,31,183,31,44,31,35,31,222,31,243,31,28,31,113,31,238,31,192,31,64,31,42,31,61,31,143,31,143,30,144,31,51,31,233,31,16,31,246,31,77,31,77,30,46,31,238,31,21,31,132,31,132,30,34,31,82,31,48,31,252,31,252,30,252,29,252,28,153,31,156,31,6,31,61,31,83,31,157,31,157,30,126,31,184,31,100,31,34,31,27,31,27,30,27,29,179,31,179,30,171,31,112,31,152,31,152,30,46,31,151,31,132,31,132,30,195,31,2,31,161,31,12,31,212,31,251,31,146,31,255,31,255,30,25,31,25,30,28,31,28,30,107,31,107,30,107,29,107,28,189,31,235,31,235,30,40,31,65,31,65,30,117,31,25,31,65,31,252,31,52,31,7,31,7,30,7,29,109,31,175,31,220,31,120,31,239,31,171,31,248,31,124,31,124,30,132,31,242,31,112,31,118,31,95,31,181,31,24,31,169,31,184,31,165,31,24,31,93,31,225,31,116,31,145,31,155,31,39,31,86,31,49,31,133,31,31,31,11,31,195,31,195,30,28,31,144,31,144,30,144,29,75,31,96,31,147,31,196,31,99,31,99,30,141,31,35,31,129,31,129,30,241,31,26,31,186,31,186,30,186,29,223,31,249,31,112,31,112,30,112,29,147,31,147,30,9,31,93,31,230,31,170,31,84,31,206,31,8,31,216,31,147,31,147,31,199,31,76,31,54,31,73,31,223,31,223,30,190,31,190,30,97,31,173,31,239,31,169,31,204,31,178,31,178,30,202,31,221,31,43,31,97,31,97,30,97,29,126,31,192,31,1,31,1,30,44,31,238,31,238,30,220,31,220,30,26,31,26,30,2,31,143,31,52,31,52,30,157,31,157,30,239,31,189,31,147,31,147,30,147,29,147,28,252,31,252,30,199,31,187,31,187,30,236,31,105,31,251,31,234,31,172,31,172,30,189,31,189,30,60,31,60,30,170,31,170,30,211,31,113,31,240,31,82,31,186,31,191,31,48,31,41,31,41,30,15,31,132,31,248,31,221,31,116,31,116,30,116,29,75,31,201,31,35,31,94,31,94,30,115,31,102,31,102,30,244,31,82,31,171,31,172,31,13,31,135,31,82,31,82,30,215,31,215,30,215,29,215,28,230,31,201,31,34,31,11,31,12,31,204,31,65,31,157,31,114,31,6,31,159,31,17,31,42,31,241,31,80,31,80,30,241,31,233,31,12,31,40,31,183,31,145,31,62,31,168,31,81,31,81,30,81,29,180,31,208,31,242,31,25,31,25,30,214,31,214,30,75,31,75,30,165,31,251,31,21,31,189,31,215,31,78,31,208,31,208,31,72,31,179,31,31,31,239,31,239,30,111,31,241,31,128,31,172,31,41,31,249,31,63,31,63,30,198,31,203,31,171,31,153,31,61,31,49,31,26,31,206,31,206,30,235,31,108,31,154,31,245,31,104,31,19,31,255,31,118,31,2,31,211,31,201,31,201,30,201,29,118,31,79,31,200,31,43,31,43,30,43,29,111,31,183,31,191,31,149,31,149,30,124,31,124,30,170,31,89,31,161,31,125,31,4,31,4,30,219,31,185,31,240,31,240,30,197,31,197,30,231,31,214,31,214,30,214,29,183,31,124,31,61,31,69,31,246,31,139,31,156,31,123,31,123,30,60,31,150,31,135,31,135,30,153,31,153,30,228,31,137,31,197,31,40,31,40,30,40,29,210,31,93,31,222,31,183,31,183,30,177,31,215,31,7,31,9,31,9,30,125,31,21,31,124,31,251,31,42,31,51,31,204,31,23,31,156,31,117,31,238,31,238,30,228,31,228,30,101,31,101,30,102,31,29,31,218,31,122,31,195,31,185,31,71,31,103,31,208,31,61,31,238,31,134,31,252,31,252,30,252,29,27,31,59,31,149,31,162,31,208,31,78,31,78,30,78,29,172,31,198,31,33,31,84,31,151,31,151,30,203,31,220,31,53,31,101,31,153,31,160,31,99,31,96,31,96,30,248,31,16,31,199,31,199,30,199,29,122,31,80,31,60,31,205,31,186,31,96,31,68,31,7,31,29,31,236,31,235,31,1,31,1,30,1,29,215,31,44,31,44,30,44,29,18,31,18,30,75,31,205,31,240,31,78,31,59,31,31,31,67,31,78,31,210,31,162,31,249,31,135,31,133,31,107,31,118,31,3,31,84,31,84,30,33,31,33,30,62,31,229,31,28,31,54,31,103,31,66,31,66,30,29,31,211,31,44,31,215,31,46,31,173,31,173,30,173,29,124,31,133,31,133,30,246,31,246,30,246,29,136,31,165,31,165,30,119,31,54,31,7,31,75,31,209,31,213,31,69,31,20,31,54,31,54,30,4,31,4,30,31,31,44,31,44,30,1,31,16,31,138,31,34,31,162,31,162,30,246,31,104,31,89,31,237,31,237,30,21,31,21,30,21,29,184,31,184,30,129,31,129,30,127,31,142,31,150,31,72,31,105,31,77,31,23,31,51,31,51,30,51,29,51,28,56,31,189,31,171,31,175,31,207,31,207,30,232,31,94,31,188,31,138,31,207,31,237,31,125,31,87,31,87,30,87,29,87,31,50,31,230,31,66,31,137,31,137,30,46,31,140,31,140,30,140,29,24,31,247,31,139,31,27,31,15,31,47,31,124,31,241,31,34,31,240,31,146,31,174,31,97,31,158,31,153,31,243,31,228,31,123,31,199,31,165,31,98,31,98,30,95,31,238,31,238,30,248,31,85,31,91,31,119,31,205,31,184,31,184,30,28,31,250,31,19,31,19,30,111,31,173,31,173,30,174,31,38,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
