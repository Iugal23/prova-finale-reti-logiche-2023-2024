-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_81 is
end project_tb_81;

architecture project_tb_arch_81 of project_tb_81 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 941;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,167,0,0,0,210,0,6,0,39,0,183,0,0,0,237,0,87,0,213,0,184,0,107,0,140,0,66,0,175,0,0,0,0,0,161,0,251,0,195,0,83,0,102,0,91,0,139,0,207,0,0,0,242,0,0,0,213,0,0,0,186,0,46,0,114,0,0,0,39,0,0,0,142,0,0,0,52,0,131,0,0,0,251,0,0,0,0,0,175,0,240,0,0,0,144,0,66,0,0,0,245,0,77,0,0,0,0,0,6,0,157,0,23,0,137,0,65,0,0,0,116,0,37,0,26,0,223,0,176,0,154,0,90,0,82,0,54,0,63,0,0,0,217,0,0,0,0,0,0,0,0,0,120,0,176,0,236,0,84,0,40,0,56,0,47,0,1,0,234,0,20,0,4,0,0,0,0,0,235,0,21,0,0,0,252,0,138,0,0,0,0,0,80,0,0,0,154,0,109,0,179,0,20,0,0,0,179,0,68,0,225,0,58,0,122,0,55,0,46,0,4,0,187,0,27,0,229,0,0,0,158,0,0,0,13,0,18,0,0,0,126,0,25,0,240,0,209,0,0,0,148,0,52,0,164,0,153,0,0,0,48,0,129,0,206,0,202,0,44,0,0,0,236,0,131,0,61,0,66,0,141,0,145,0,200,0,45,0,97,0,205,0,0,0,0,0,206,0,11,0,144,0,248,0,67,0,0,0,84,0,14,0,83,0,19,0,195,0,152,0,28,0,122,0,0,0,181,0,161,0,15,0,0,0,34,0,0,0,170,0,0,0,196,0,253,0,80,0,196,0,243,0,173,0,0,0,194,0,102,0,71,0,233,0,66,0,207,0,164,0,32,0,98,0,188,0,172,0,171,0,0,0,141,0,58,0,116,0,103,0,0,0,235,0,70,0,0,0,170,0,227,0,190,0,201,0,124,0,127,0,102,0,231,0,236,0,0,0,255,0,226,0,0,0,132,0,15,0,211,0,0,0,83,0,207,0,215,0,35,0,224,0,125,0,0,0,23,0,71,0,98,0,20,0,0,0,43,0,177,0,81,0,46,0,199,0,0,0,116,0,0,0,52,0,97,0,171,0,173,0,0,0,97,0,0,0,5,0,0,0,0,0,199,0,137,0,0,0,93,0,93,0,0,0,47,0,234,0,185,0,52,0,175,0,0,0,0,0,95,0,0,0,210,0,54,0,204,0,71,0,111,0,0,0,67,0,0,0,0,0,18,0,44,0,212,0,193,0,0,0,241,0,0,0,72,0,44,0,244,0,121,0,37,0,168,0,65,0,199,0,197,0,108,0,0,0,151,0,17,0,110,0,0,0,64,0,20,0,211,0,169,0,165,0,160,0,92,0,235,0,16,0,0,0,0,0,32,0,178,0,162,0,0,0,177,0,86,0,79,0,141,0,219,0,134,0,0,0,88,0,31,0,188,0,210,0,0,0,0,0,231,0,227,0,27,0,35,0,0,0,0,0,33,0,43,0,60,0,0,0,7,0,0,0,84,0,0,0,135,0,248,0,93,0,151,0,224,0,57,0,215,0,249,0,186,0,44,0,117,0,218,0,47,0,75,0,46,0,110,0,18,0,142,0,187,0,0,0,182,0,0,0,254,0,84,0,0,0,194,0,50,0,44,0,47,0,179,0,172,0,251,0,0,0,138,0,247,0,118,0,10,0,1,0,224,0,208,0,104,0,112,0,176,0,104,0,246,0,194,0,124,0,12,0,158,0,0,0,18,0,0,0,127,0,11,0,252,0,114,0,165,0,0,0,179,0,0,0,245,0,65,0,91,0,0,0,0,0,158,0,209,0,199,0,0,0,148,0,118,0,105,0,193,0,244,0,190,0,0,0,0,0,0,0,28,0,170,0,193,0,0,0,111,0,0,0,0,0,0,0,116,0,89,0,127,0,131,0,11,0,0,0,5,0,130,0,0,0,117,0,0,0,203,0,190,0,37,0,214,0,105,0,15,0,204,0,229,0,14,0,0,0,61,0,163,0,239,0,99,0,0,0,146,0,221,0,68,0,193,0,73,0,100,0,13,0,125,0,0,0,0,0,0,0,71,0,120,0,110,0,65,0,113,0,66,0,101,0,143,0,214,0,84,0,16,0,225,0,0,0,91,0,76,0,251,0,156,0,132,0,232,0,40,0,0,0,245,0,108,0,0,0,108,0,110,0,208,0,0,0,0,0,204,0,250,0,27,0,64,0,163,0,39,0,192,0,240,0,205,0,84,0,120,0,124,0,228,0,198,0,127,0,0,0,0,0,182,0,166,0,0,0,203,0,90,0,166,0,166,0,94,0,0,0,250,0,227,0,153,0,198,0,42,0,105,0,19,0,0,0,10,0,234,0,84,0,102,0,0,0,170,0,195,0,174,0,0,0,212,0,0,0,54,0,202,0,68,0,0,0,156,0,238,0,3,0,154,0,25,0,176,0,55,0,0,0,142,0,49,0,0,0,0,0,47,0,50,0,222,0,87,0,0,0,216,0,0,0,59,0,182,0,0,0,51,0,41,0,49,0,203,0,23,0,185,0,7,0,107,0,0,0,93,0,0,0,0,0,0,0,232,0,49,0,0,0,0,0,109,0,127,0,0,0,0,0,3,0,93,0,181,0,204,0,237,0,0,0,145,0,215,0,0,0,44,0,251,0,184,0,0,0,46,0,34,0,0,0,158,0,195,0,148,0,0,0,37,0,151,0,100,0,246,0,0,0,215,0,237,0,141,0,141,0,0,0,93,0,158,0,194,0,163,0,0,0,242,0,1,0,191,0,145,0,19,0,0,0,17,0,244,0,0,0,194,0,233,0,81,0,171,0,223,0,138,0,76,0,0,0,0,0,67,0,0,0,38,0,0,0,68,0,65,0,42,0,174,0,148,0,130,0,88,0,28,0,159,0,16,0,0,0,254,0,176,0,144,0,234,0,8,0,16,0,66,0,219,0,0,0,202,0,171,0,71,0,0,0,155,0,160,0,233,0,215,0,88,0,126,0,149,0,9,0,105,0,239,0,43,0,33,0,151,0,61,0,32,0,76,0,219,0,0,0,0,0,7,0,0,0,0,0,55,0,0,0,222,0,154,0,0,0,243,0,119,0,144,0,106,0,111,0,164,0,10,0,53,0,0,0,0,0,147,0,0,0,0,0,48,0,41,0,7,0,86,0,61,0,211,0,155,0,72,0,169,0,31,0,221,0,17,0,37,0,0,0,214,0,236,0,44,0,191,0,105,0,251,0,157,0,94,0,211,0,229,0,0,0,208,0,8,0,2,0,0,0,22,0,0,0,0,0,90,0,0,0,69,0,0,0,58,0,169,0,0,0,0,0,179,0,80,0,0,0,104,0,196,0,140,0,125,0,0,0,0,0,8,0,148,0,0,0,181,0,0,0,245,0,0,0,208,0,78,0,197,0,169,0,222,0,0,0,64,0,18,0,0,0,209,0,0,0,156,0,199,0,211,0,206,0,250,0,0,0,212,0,103,0,42,0,207,0,218,0,66,0,233,0,167,0,140,0,115,0,0,0,53,0,238,0,27,0,29,0,51,0,180,0,94,0,128,0,18,0,59,0,136,0,0,0,52,0,60,0,0,0,43,0,180,0,3,0,0,0,0,0,119,0,30,0,28,0,45,0,127,0,150,0,137,0,53,0,155,0,243,0,228,0,228,0,245,0,178,0,0,0,246,0,16,0,103,0,0,0,126,0,78,0,0,0,197,0,139,0,221,0,101,0,0,0,93,0,80,0,231,0,95,0,147,0,127,0,0,0,65,0,164,0,0,0,134,0,206,0,0,0,75,0,204,0,0,0,108,0,195,0,173,0,207,0,208,0,0,0,0,0,0,0,0,0,255,0,75,0,114,0,173,0,41,0,127,0,37,0,52,0,207,0,24,0,252,0,208,0,169,0,245,0,160,0,84,0,86,0,174,0,8,0,8,0,237,0,119,0,250,0,81,0,201,0,214,0,230,0,92,0,161,0,237,0,0,0,53,0,0,0,0,0,21,0,185,0,99,0,205,0,58,0,0,0,0,0,0,0,239,0,253,0,0,0,211,0,179,0,0,0,0,0,18,0,40,0,3,0,171,0,0,0,224,0,20,0,133,0,0,0,81,0,0,0,188,0,0,0,35,0,168,0,82,0,0,0,126,0,24,0,220,0,202,0,88,0,0,0,182,0,0,0,191,0,125,0,236,0,100,0,118,0,206,0,0,0,19,0,134,0,250,0,254,0);
signal scenario_full  : scenario_type := (0,0,167,31,167,30,210,31,6,31,39,31,183,31,183,30,237,31,87,31,213,31,184,31,107,31,140,31,66,31,175,31,175,30,175,29,161,31,251,31,195,31,83,31,102,31,91,31,139,31,207,31,207,30,242,31,242,30,213,31,213,30,186,31,46,31,114,31,114,30,39,31,39,30,142,31,142,30,52,31,131,31,131,30,251,31,251,30,251,29,175,31,240,31,240,30,144,31,66,31,66,30,245,31,77,31,77,30,77,29,6,31,157,31,23,31,137,31,65,31,65,30,116,31,37,31,26,31,223,31,176,31,154,31,90,31,82,31,54,31,63,31,63,30,217,31,217,30,217,29,217,28,217,27,120,31,176,31,236,31,84,31,40,31,56,31,47,31,1,31,234,31,20,31,4,31,4,30,4,29,235,31,21,31,21,30,252,31,138,31,138,30,138,29,80,31,80,30,154,31,109,31,179,31,20,31,20,30,179,31,68,31,225,31,58,31,122,31,55,31,46,31,4,31,187,31,27,31,229,31,229,30,158,31,158,30,13,31,18,31,18,30,126,31,25,31,240,31,209,31,209,30,148,31,52,31,164,31,153,31,153,30,48,31,129,31,206,31,202,31,44,31,44,30,236,31,131,31,61,31,66,31,141,31,145,31,200,31,45,31,97,31,205,31,205,30,205,29,206,31,11,31,144,31,248,31,67,31,67,30,84,31,14,31,83,31,19,31,195,31,152,31,28,31,122,31,122,30,181,31,161,31,15,31,15,30,34,31,34,30,170,31,170,30,196,31,253,31,80,31,196,31,243,31,173,31,173,30,194,31,102,31,71,31,233,31,66,31,207,31,164,31,32,31,98,31,188,31,172,31,171,31,171,30,141,31,58,31,116,31,103,31,103,30,235,31,70,31,70,30,170,31,227,31,190,31,201,31,124,31,127,31,102,31,231,31,236,31,236,30,255,31,226,31,226,30,132,31,15,31,211,31,211,30,83,31,207,31,215,31,35,31,224,31,125,31,125,30,23,31,71,31,98,31,20,31,20,30,43,31,177,31,81,31,46,31,199,31,199,30,116,31,116,30,52,31,97,31,171,31,173,31,173,30,97,31,97,30,5,31,5,30,5,29,199,31,137,31,137,30,93,31,93,31,93,30,47,31,234,31,185,31,52,31,175,31,175,30,175,29,95,31,95,30,210,31,54,31,204,31,71,31,111,31,111,30,67,31,67,30,67,29,18,31,44,31,212,31,193,31,193,30,241,31,241,30,72,31,44,31,244,31,121,31,37,31,168,31,65,31,199,31,197,31,108,31,108,30,151,31,17,31,110,31,110,30,64,31,20,31,211,31,169,31,165,31,160,31,92,31,235,31,16,31,16,30,16,29,32,31,178,31,162,31,162,30,177,31,86,31,79,31,141,31,219,31,134,31,134,30,88,31,31,31,188,31,210,31,210,30,210,29,231,31,227,31,27,31,35,31,35,30,35,29,33,31,43,31,60,31,60,30,7,31,7,30,84,31,84,30,135,31,248,31,93,31,151,31,224,31,57,31,215,31,249,31,186,31,44,31,117,31,218,31,47,31,75,31,46,31,110,31,18,31,142,31,187,31,187,30,182,31,182,30,254,31,84,31,84,30,194,31,50,31,44,31,47,31,179,31,172,31,251,31,251,30,138,31,247,31,118,31,10,31,1,31,224,31,208,31,104,31,112,31,176,31,104,31,246,31,194,31,124,31,12,31,158,31,158,30,18,31,18,30,127,31,11,31,252,31,114,31,165,31,165,30,179,31,179,30,245,31,65,31,91,31,91,30,91,29,158,31,209,31,199,31,199,30,148,31,118,31,105,31,193,31,244,31,190,31,190,30,190,29,190,28,28,31,170,31,193,31,193,30,111,31,111,30,111,29,111,28,116,31,89,31,127,31,131,31,11,31,11,30,5,31,130,31,130,30,117,31,117,30,203,31,190,31,37,31,214,31,105,31,15,31,204,31,229,31,14,31,14,30,61,31,163,31,239,31,99,31,99,30,146,31,221,31,68,31,193,31,73,31,100,31,13,31,125,31,125,30,125,29,125,28,71,31,120,31,110,31,65,31,113,31,66,31,101,31,143,31,214,31,84,31,16,31,225,31,225,30,91,31,76,31,251,31,156,31,132,31,232,31,40,31,40,30,245,31,108,31,108,30,108,31,110,31,208,31,208,30,208,29,204,31,250,31,27,31,64,31,163,31,39,31,192,31,240,31,205,31,84,31,120,31,124,31,228,31,198,31,127,31,127,30,127,29,182,31,166,31,166,30,203,31,90,31,166,31,166,31,94,31,94,30,250,31,227,31,153,31,198,31,42,31,105,31,19,31,19,30,10,31,234,31,84,31,102,31,102,30,170,31,195,31,174,31,174,30,212,31,212,30,54,31,202,31,68,31,68,30,156,31,238,31,3,31,154,31,25,31,176,31,55,31,55,30,142,31,49,31,49,30,49,29,47,31,50,31,222,31,87,31,87,30,216,31,216,30,59,31,182,31,182,30,51,31,41,31,49,31,203,31,23,31,185,31,7,31,107,31,107,30,93,31,93,30,93,29,93,28,232,31,49,31,49,30,49,29,109,31,127,31,127,30,127,29,3,31,93,31,181,31,204,31,237,31,237,30,145,31,215,31,215,30,44,31,251,31,184,31,184,30,46,31,34,31,34,30,158,31,195,31,148,31,148,30,37,31,151,31,100,31,246,31,246,30,215,31,237,31,141,31,141,31,141,30,93,31,158,31,194,31,163,31,163,30,242,31,1,31,191,31,145,31,19,31,19,30,17,31,244,31,244,30,194,31,233,31,81,31,171,31,223,31,138,31,76,31,76,30,76,29,67,31,67,30,38,31,38,30,68,31,65,31,42,31,174,31,148,31,130,31,88,31,28,31,159,31,16,31,16,30,254,31,176,31,144,31,234,31,8,31,16,31,66,31,219,31,219,30,202,31,171,31,71,31,71,30,155,31,160,31,233,31,215,31,88,31,126,31,149,31,9,31,105,31,239,31,43,31,33,31,151,31,61,31,32,31,76,31,219,31,219,30,219,29,7,31,7,30,7,29,55,31,55,30,222,31,154,31,154,30,243,31,119,31,144,31,106,31,111,31,164,31,10,31,53,31,53,30,53,29,147,31,147,30,147,29,48,31,41,31,7,31,86,31,61,31,211,31,155,31,72,31,169,31,31,31,221,31,17,31,37,31,37,30,214,31,236,31,44,31,191,31,105,31,251,31,157,31,94,31,211,31,229,31,229,30,208,31,8,31,2,31,2,30,22,31,22,30,22,29,90,31,90,30,69,31,69,30,58,31,169,31,169,30,169,29,179,31,80,31,80,30,104,31,196,31,140,31,125,31,125,30,125,29,8,31,148,31,148,30,181,31,181,30,245,31,245,30,208,31,78,31,197,31,169,31,222,31,222,30,64,31,18,31,18,30,209,31,209,30,156,31,199,31,211,31,206,31,250,31,250,30,212,31,103,31,42,31,207,31,218,31,66,31,233,31,167,31,140,31,115,31,115,30,53,31,238,31,27,31,29,31,51,31,180,31,94,31,128,31,18,31,59,31,136,31,136,30,52,31,60,31,60,30,43,31,180,31,3,31,3,30,3,29,119,31,30,31,28,31,45,31,127,31,150,31,137,31,53,31,155,31,243,31,228,31,228,31,245,31,178,31,178,30,246,31,16,31,103,31,103,30,126,31,78,31,78,30,197,31,139,31,221,31,101,31,101,30,93,31,80,31,231,31,95,31,147,31,127,31,127,30,65,31,164,31,164,30,134,31,206,31,206,30,75,31,204,31,204,30,108,31,195,31,173,31,207,31,208,31,208,30,208,29,208,28,208,27,255,31,75,31,114,31,173,31,41,31,127,31,37,31,52,31,207,31,24,31,252,31,208,31,169,31,245,31,160,31,84,31,86,31,174,31,8,31,8,31,237,31,119,31,250,31,81,31,201,31,214,31,230,31,92,31,161,31,237,31,237,30,53,31,53,30,53,29,21,31,185,31,99,31,205,31,58,31,58,30,58,29,58,28,239,31,253,31,253,30,211,31,179,31,179,30,179,29,18,31,40,31,3,31,171,31,171,30,224,31,20,31,133,31,133,30,81,31,81,30,188,31,188,30,35,31,168,31,82,31,82,30,126,31,24,31,220,31,202,31,88,31,88,30,182,31,182,30,191,31,125,31,236,31,100,31,118,31,206,31,206,30,19,31,134,31,250,31,254,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
