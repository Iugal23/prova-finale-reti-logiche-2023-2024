-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 340;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,178,0,171,0,156,0,84,0,124,0,0,0,19,0,95,0,173,0,0,0,125,0,40,0,30,0,111,0,0,0,32,0,132,0,141,0,214,0,142,0,228,0,25,0,0,0,163,0,114,0,0,0,101,0,30,0,181,0,146,0,7,0,89,0,171,0,54,0,0,0,34,0,0,0,125,0,203,0,212,0,0,0,139,0,120,0,207,0,113,0,22,0,179,0,219,0,210,0,181,0,87,0,124,0,0,0,125,0,11,0,25,0,194,0,0,0,91,0,156,0,78,0,186,0,0,0,0,0,4,0,200,0,92,0,128,0,134,0,19,0,78,0,113,0,81,0,0,0,74,0,0,0,202,0,0,0,248,0,166,0,169,0,123,0,167,0,209,0,83,0,176,0,220,0,0,0,0,0,0,0,105,0,145,0,180,0,53,0,112,0,86,0,0,0,14,0,244,0,130,0,216,0,158,0,112,0,112,0,50,0,0,0,89,0,80,0,163,0,50,0,0,0,202,0,0,0,112,0,224,0,29,0,122,0,226,0,109,0,198,0,181,0,108,0,150,0,186,0,192,0,13,0,1,0,17,0,34,0,51,0,65,0,188,0,204,0,208,0,40,0,135,0,222,0,236,0,7,0,111,0,13,0,0,0,246,0,56,0,59,0,215,0,184,0,20,0,172,0,0,0,218,0,85,0,133,0,229,0,105,0,141,0,14,0,78,0,61,0,21,0,198,0,114,0,244,0,171,0,0,0,0,0,0,0,2,0,38,0,138,0,133,0,90,0,198,0,93,0,94,0,14,0,198,0,145,0,206,0,14,0,111,0,188,0,65,0,0,0,48,0,119,0,42,0,40,0,0,0,174,0,202,0,166,0,0,0,237,0,217,0,12,0,0,0,23,0,0,0,189,0,246,0,83,0,31,0,189,0,66,0,0,0,213,0,0,0,98,0,155,0,0,0,193,0,40,0,244,0,180,0,85,0,80,0,120,0,240,0,0,0,94,0,154,0,66,0,0,0,119,0,109,0,128,0,201,0,0,0,172,0,148,0,40,0,0,0,139,0,209,0,0,0,47,0,37,0,156,0,246,0,205,0,180,0,189,0,119,0,111,0,210,0,207,0,196,0,121,0,236,0,78,0,46,0,209,0,57,0,71,0,191,0,0,0,219,0,37,0,69,0,0,0,199,0,230,0,145,0,213,0,222,0,0,0,188,0,0,0,81,0,110,0,184,0,61,0,245,0,166,0,104,0,0,0,0,0,115,0,172,0,0,0,169,0,82,0,23,0,93,0,185,0,124,0,0,0,181,0,0,0,233,0,188,0,0,0,186,0,42,0,89,0,0,0,219,0,25,0,217,0,134,0,175,0,6,0,0,0,37,0,250,0,217,0,179,0,39,0,184,0,126,0,91,0,59,0,70,0,212,0,125,0,66,0,150,0,35,0,213,0,0,0,0,0,246,0,140,0,34,0,41,0,50,0,102,0,149,0,80,0,35,0,137,0,39,0,169,0,202,0,153,0,249,0,53,0,243,0);
signal scenario_full  : scenario_type := (0,0,178,31,171,31,156,31,84,31,124,31,124,30,19,31,95,31,173,31,173,30,125,31,40,31,30,31,111,31,111,30,32,31,132,31,141,31,214,31,142,31,228,31,25,31,25,30,163,31,114,31,114,30,101,31,30,31,181,31,146,31,7,31,89,31,171,31,54,31,54,30,34,31,34,30,125,31,203,31,212,31,212,30,139,31,120,31,207,31,113,31,22,31,179,31,219,31,210,31,181,31,87,31,124,31,124,30,125,31,11,31,25,31,194,31,194,30,91,31,156,31,78,31,186,31,186,30,186,29,4,31,200,31,92,31,128,31,134,31,19,31,78,31,113,31,81,31,81,30,74,31,74,30,202,31,202,30,248,31,166,31,169,31,123,31,167,31,209,31,83,31,176,31,220,31,220,30,220,29,220,28,105,31,145,31,180,31,53,31,112,31,86,31,86,30,14,31,244,31,130,31,216,31,158,31,112,31,112,31,50,31,50,30,89,31,80,31,163,31,50,31,50,30,202,31,202,30,112,31,224,31,29,31,122,31,226,31,109,31,198,31,181,31,108,31,150,31,186,31,192,31,13,31,1,31,17,31,34,31,51,31,65,31,188,31,204,31,208,31,40,31,135,31,222,31,236,31,7,31,111,31,13,31,13,30,246,31,56,31,59,31,215,31,184,31,20,31,172,31,172,30,218,31,85,31,133,31,229,31,105,31,141,31,14,31,78,31,61,31,21,31,198,31,114,31,244,31,171,31,171,30,171,29,171,28,2,31,38,31,138,31,133,31,90,31,198,31,93,31,94,31,14,31,198,31,145,31,206,31,14,31,111,31,188,31,65,31,65,30,48,31,119,31,42,31,40,31,40,30,174,31,202,31,166,31,166,30,237,31,217,31,12,31,12,30,23,31,23,30,189,31,246,31,83,31,31,31,189,31,66,31,66,30,213,31,213,30,98,31,155,31,155,30,193,31,40,31,244,31,180,31,85,31,80,31,120,31,240,31,240,30,94,31,154,31,66,31,66,30,119,31,109,31,128,31,201,31,201,30,172,31,148,31,40,31,40,30,139,31,209,31,209,30,47,31,37,31,156,31,246,31,205,31,180,31,189,31,119,31,111,31,210,31,207,31,196,31,121,31,236,31,78,31,46,31,209,31,57,31,71,31,191,31,191,30,219,31,37,31,69,31,69,30,199,31,230,31,145,31,213,31,222,31,222,30,188,31,188,30,81,31,110,31,184,31,61,31,245,31,166,31,104,31,104,30,104,29,115,31,172,31,172,30,169,31,82,31,23,31,93,31,185,31,124,31,124,30,181,31,181,30,233,31,188,31,188,30,186,31,42,31,89,31,89,30,219,31,25,31,217,31,134,31,175,31,6,31,6,30,37,31,250,31,217,31,179,31,39,31,184,31,126,31,91,31,59,31,70,31,212,31,125,31,66,31,150,31,35,31,213,31,213,30,213,29,246,31,140,31,34,31,41,31,50,31,102,31,149,31,80,31,35,31,137,31,39,31,169,31,202,31,153,31,249,31,53,31,243,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
