-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1011;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (165,0,32,0,212,0,22,0,92,0,135,0,0,0,255,0,102,0,87,0,79,0,107,0,227,0,0,0,148,0,102,0,79,0,131,0,36,0,0,0,0,0,248,0,0,0,0,0,182,0,0,0,254,0,0,0,25,0,127,0,90,0,9,0,0,0,0,0,151,0,152,0,220,0,160,0,130,0,140,0,61,0,252,0,229,0,224,0,131,0,30,0,0,0,238,0,0,0,39,0,0,0,224,0,117,0,0,0,166,0,193,0,182,0,75,0,0,0,128,0,201,0,117,0,13,0,188,0,10,0,41,0,69,0,0,0,174,0,117,0,211,0,97,0,81,0,198,0,134,0,195,0,30,0,145,0,182,0,0,0,243,0,68,0,211,0,153,0,100,0,0,0,20,0,237,0,38,0,0,0,0,0,126,0,0,0,97,0,0,0,63,0,53,0,203,0,50,0,80,0,0,0,105,0,160,0,0,0,169,0,68,0,150,0,66,0,2,0,0,0,170,0,53,0,0,0,9,0,11,0,0,0,65,0,208,0,0,0,127,0,36,0,144,0,173,0,21,0,226,0,61,0,236,0,11,0,174,0,0,0,187,0,0,0,0,0,221,0,0,0,136,0,254,0,0,0,231,0,144,0,222,0,251,0,0,0,140,0,0,0,0,0,121,0,126,0,241,0,0,0,197,0,177,0,239,0,0,0,243,0,0,0,9,0,101,0,149,0,80,0,0,0,163,0,83,0,0,0,40,0,195,0,27,0,200,0,88,0,160,0,39,0,9,0,238,0,0,0,0,0,185,0,109,0,242,0,0,0,138,0,189,0,60,0,85,0,234,0,34,0,65,0,174,0,188,0,67,0,245,0,0,0,238,0,0,0,0,0,135,0,0,0,102,0,162,0,83,0,79,0,91,0,0,0,0,0,60,0,237,0,54,0,118,0,103,0,79,0,0,0,73,0,166,0,29,0,0,0,251,0,182,0,209,0,29,0,152,0,0,0,60,0,0,0,98,0,16,0,114,0,0,0,0,0,0,0,0,0,70,0,17,0,122,0,102,0,81,0,65,0,120,0,188,0,96,0,26,0,96,0,190,0,228,0,243,0,10,0,182,0,183,0,81,0,120,0,53,0,151,0,232,0,46,0,254,0,0,0,0,0,0,0,151,0,0,0,98,0,206,0,250,0,8,0,250,0,95,0,19,0,0,0,128,0,61,0,0,0,0,0,181,0,219,0,0,0,48,0,84,0,107,0,0,0,164,0,45,0,0,0,158,0,6,0,97,0,0,0,204,0,6,0,0,0,4,0,9,0,63,0,0,0,191,0,36,0,244,0,230,0,184,0,74,0,195,0,128,0,162,0,160,0,22,0,162,0,108,0,124,0,133,0,226,0,194,0,209,0,161,0,146,0,209,0,85,0,153,0,239,0,0,0,0,0,0,0,70,0,7,0,238,0,254,0,83,0,211,0,165,0,215,0,114,0,0,0,242,0,159,0,135,0,198,0,208,0,167,0,75,0,0,0,179,0,243,0,97,0,0,0,0,0,174,0,121,0,41,0,63,0,225,0,168,0,156,0,0,0,0,0,0,0,8,0,0,0,90,0,146,0,33,0,173,0,31,0,53,0,0,0,0,0,0,0,25,0,180,0,128,0,232,0,147,0,200,0,118,0,246,0,115,0,22,0,130,0,219,0,107,0,109,0,153,0,171,0,0,0,137,0,209,0,76,0,168,0,220,0,36,0,215,0,51,0,195,0,0,0,247,0,0,0,107,0,75,0,213,0,47,0,150,0,54,0,4,0,0,0,142,0,44,0,0,0,199,0,203,0,128,0,72,0,68,0,0,0,152,0,6,0,141,0,27,0,0,0,154,0,0,0,165,0,0,0,0,0,53,0,231,0,0,0,0,0,82,0,76,0,144,0,0,0,201,0,35,0,0,0,155,0,23,0,101,0,78,0,205,0,0,0,253,0,137,0,130,0,1,0,68,0,0,0,168,0,8,0,0,0,182,0,0,0,149,0,33,0,240,0,145,0,0,0,0,0,43,0,231,0,0,0,0,0,73,0,83,0,110,0,0,0,91,0,220,0,117,0,0,0,185,0,0,0,130,0,159,0,32,0,107,0,115,0,159,0,232,0,232,0,9,0,0,0,107,0,35,0,0,0,79,0,123,0,174,0,80,0,7,0,237,0,186,0,15,0,186,0,40,0,90,0,0,0,185,0,222,0,249,0,161,0,194,0,156,0,246,0,191,0,122,0,179,0,151,0,0,0,77,0,218,0,31,0,185,0,192,0,103,0,219,0,74,0,186,0,173,0,0,0,148,0,107,0,118,0,7,0,0,0,156,0,146,0,0,0,201,0,27,0,93,0,21,0,129,0,75,0,132,0,239,0,210,0,163,0,231,0,53,0,171,0,184,0,126,0,0,0,235,0,242,0,169,0,173,0,149,0,142,0,0,0,0,0,0,0,141,0,155,0,41,0,145,0,220,0,221,0,86,0,247,0,162,0,226,0,147,0,230,0,64,0,0,0,0,0,129,0,196,0,0,0,100,0,0,0,36,0,0,0,88,0,1,0,0,0,156,0,171,0,201,0,121,0,64,0,171,0,153,0,184,0,89,0,202,0,67,0,193,0,52,0,196,0,127,0,231,0,92,0,122,0,37,0,247,0,184,0,126,0,0,0,241,0,157,0,124,0,221,0,157,0,67,0,0,0,204,0,106,0,0,0,38,0,170,0,117,0,1,0,63,0,231,0,97,0,100,0,0,0,165,0,66,0,44,0,81,0,8,0,0,0,25,0,247,0,113,0,251,0,7,0,182,0,0,0,165,0,192,0,251,0,67,0,153,0,233,0,47,0,19,0,28,0,102,0,239,0,182,0,0,0,32,0,225,0,17,0,4,0,218,0,238,0,17,0,99,0,210,0,129,0,9,0,83,0,0,0,152,0,56,0,24,0,121,0,115,0,251,0,247,0,57,0,0,0,29,0,191,0,110,0,219,0,145,0,6,0,0,0,51,0,73,0,100,0,0,0,0,0,245,0,152,0,122,0,57,0,76,0,191,0,55,0,58,0,39,0,24,0,74,0,187,0,229,0,113,0,0,0,111,0,3,0,40,0,109,0,67,0,167,0,81,0,172,0,231,0,246,0,0,0,0,0,76,0,11,0,0,0,155,0,68,0,112,0,68,0,55,0,152,0,219,0,0,0,0,0,54,0,2,0,0,0,171,0,0,0,255,0,194,0,57,0,235,0,97,0,213,0,0,0,0,0,0,0,4,0,193,0,21,0,0,0,0,0,77,0,82,0,0,0,205,0,77,0,0,0,0,0,200,0,30,0,0,0,0,0,255,0,209,0,247,0,244,0,49,0,147,0,167,0,0,0,0,0,231,0,0,0,38,0,189,0,36,0,40,0,145,0,205,0,96,0,0,0,14,0,243,0,62,0,0,0,0,0,102,0,162,0,55,0,209,0,0,0,2,0,220,0,114,0,0,0,0,0,211,0,204,0,60,0,227,0,188,0,31,0,85,0,55,0,97,0,245,0,187,0,5,0,163,0,155,0,176,0,0,0,235,0,0,0,90,0,217,0,146,0,122,0,127,0,156,0,184,0,53,0,160,0,172,0,56,0,0,0,247,0,7,0,0,0,167,0,117,0,94,0,62,0,26,0,244,0,96,0,62,0,0,0,146,0,43,0,214,0,37,0,42,0,243,0,224,0,208,0,0,0,221,0,163,0,189,0,13,0,228,0,69,0,0,0,253,0,0,0,140,0,63,0,208,0,0,0,0,0,227,0,54,0,0,0,211,0,25,0,160,0,76,0,87,0,88,0,21,0,252,0,166,0,176,0,0,0,0,0,43,0,3,0,2,0,206,0,0,0,123,0,140,0,54,0,11,0,131,0,0,0,57,0,118,0,0,0,0,0,100,0,53,0,242,0,177,0,0,0,129,0,2,0,0,0,145,0,139,0,123,0,248,0,72,0,26,0,99,0,227,0,0,0,0,0,236,0,0,0,0,0,0,0,41,0,8,0,183,0,65,0,79,0,0,0,229,0,175,0,105,0,195,0,91,0,141,0,132,0,0,0,84,0,0,0,78,0,0,0,229,0,0,0,13,0,53,0,45,0,6,0,0,0,115,0,114,0,105,0,48,0,28,0,225,0,102,0,92,0,209,0,6,0,118,0,231,0,0,0,131,0,43,0,0,0,42,0,9,0,68,0,64,0,84,0,193,0,0,0,108,0,0,0,68,0,178,0,0,0,34,0,217,0,234,0,255,0,79,0,0,0,170,0,113,0,73,0,152,0,60,0,12,0,30,0,135,0,34,0,161,0,132,0,29,0,75,0,112,0,0,0,121,0,102,0,0,0,229,0,57,0,229,0,92,0,0,0,121,0,197,0,5,0,26,0,0,0,140,0,0,0,50,0,48,0,74,0,168,0,0,0,232,0,49,0,187,0,18,0,32,0,3,0,137,0,153,0,0,0,14,0,0,0,0,0,0,0,0,0,0,0,219,0,196,0,68,0,226,0,202,0,0,0,0,0,0,0);
signal scenario_full  : scenario_type := (165,31,32,31,212,31,22,31,92,31,135,31,135,30,255,31,102,31,87,31,79,31,107,31,227,31,227,30,148,31,102,31,79,31,131,31,36,31,36,30,36,29,248,31,248,30,248,29,182,31,182,30,254,31,254,30,25,31,127,31,90,31,9,31,9,30,9,29,151,31,152,31,220,31,160,31,130,31,140,31,61,31,252,31,229,31,224,31,131,31,30,31,30,30,238,31,238,30,39,31,39,30,224,31,117,31,117,30,166,31,193,31,182,31,75,31,75,30,128,31,201,31,117,31,13,31,188,31,10,31,41,31,69,31,69,30,174,31,117,31,211,31,97,31,81,31,198,31,134,31,195,31,30,31,145,31,182,31,182,30,243,31,68,31,211,31,153,31,100,31,100,30,20,31,237,31,38,31,38,30,38,29,126,31,126,30,97,31,97,30,63,31,53,31,203,31,50,31,80,31,80,30,105,31,160,31,160,30,169,31,68,31,150,31,66,31,2,31,2,30,170,31,53,31,53,30,9,31,11,31,11,30,65,31,208,31,208,30,127,31,36,31,144,31,173,31,21,31,226,31,61,31,236,31,11,31,174,31,174,30,187,31,187,30,187,29,221,31,221,30,136,31,254,31,254,30,231,31,144,31,222,31,251,31,251,30,140,31,140,30,140,29,121,31,126,31,241,31,241,30,197,31,177,31,239,31,239,30,243,31,243,30,9,31,101,31,149,31,80,31,80,30,163,31,83,31,83,30,40,31,195,31,27,31,200,31,88,31,160,31,39,31,9,31,238,31,238,30,238,29,185,31,109,31,242,31,242,30,138,31,189,31,60,31,85,31,234,31,34,31,65,31,174,31,188,31,67,31,245,31,245,30,238,31,238,30,238,29,135,31,135,30,102,31,162,31,83,31,79,31,91,31,91,30,91,29,60,31,237,31,54,31,118,31,103,31,79,31,79,30,73,31,166,31,29,31,29,30,251,31,182,31,209,31,29,31,152,31,152,30,60,31,60,30,98,31,16,31,114,31,114,30,114,29,114,28,114,27,70,31,17,31,122,31,102,31,81,31,65,31,120,31,188,31,96,31,26,31,96,31,190,31,228,31,243,31,10,31,182,31,183,31,81,31,120,31,53,31,151,31,232,31,46,31,254,31,254,30,254,29,254,28,151,31,151,30,98,31,206,31,250,31,8,31,250,31,95,31,19,31,19,30,128,31,61,31,61,30,61,29,181,31,219,31,219,30,48,31,84,31,107,31,107,30,164,31,45,31,45,30,158,31,6,31,97,31,97,30,204,31,6,31,6,30,4,31,9,31,63,31,63,30,191,31,36,31,244,31,230,31,184,31,74,31,195,31,128,31,162,31,160,31,22,31,162,31,108,31,124,31,133,31,226,31,194,31,209,31,161,31,146,31,209,31,85,31,153,31,239,31,239,30,239,29,239,28,70,31,7,31,238,31,254,31,83,31,211,31,165,31,215,31,114,31,114,30,242,31,159,31,135,31,198,31,208,31,167,31,75,31,75,30,179,31,243,31,97,31,97,30,97,29,174,31,121,31,41,31,63,31,225,31,168,31,156,31,156,30,156,29,156,28,8,31,8,30,90,31,146,31,33,31,173,31,31,31,53,31,53,30,53,29,53,28,25,31,180,31,128,31,232,31,147,31,200,31,118,31,246,31,115,31,22,31,130,31,219,31,107,31,109,31,153,31,171,31,171,30,137,31,209,31,76,31,168,31,220,31,36,31,215,31,51,31,195,31,195,30,247,31,247,30,107,31,75,31,213,31,47,31,150,31,54,31,4,31,4,30,142,31,44,31,44,30,199,31,203,31,128,31,72,31,68,31,68,30,152,31,6,31,141,31,27,31,27,30,154,31,154,30,165,31,165,30,165,29,53,31,231,31,231,30,231,29,82,31,76,31,144,31,144,30,201,31,35,31,35,30,155,31,23,31,101,31,78,31,205,31,205,30,253,31,137,31,130,31,1,31,68,31,68,30,168,31,8,31,8,30,182,31,182,30,149,31,33,31,240,31,145,31,145,30,145,29,43,31,231,31,231,30,231,29,73,31,83,31,110,31,110,30,91,31,220,31,117,31,117,30,185,31,185,30,130,31,159,31,32,31,107,31,115,31,159,31,232,31,232,31,9,31,9,30,107,31,35,31,35,30,79,31,123,31,174,31,80,31,7,31,237,31,186,31,15,31,186,31,40,31,90,31,90,30,185,31,222,31,249,31,161,31,194,31,156,31,246,31,191,31,122,31,179,31,151,31,151,30,77,31,218,31,31,31,185,31,192,31,103,31,219,31,74,31,186,31,173,31,173,30,148,31,107,31,118,31,7,31,7,30,156,31,146,31,146,30,201,31,27,31,93,31,21,31,129,31,75,31,132,31,239,31,210,31,163,31,231,31,53,31,171,31,184,31,126,31,126,30,235,31,242,31,169,31,173,31,149,31,142,31,142,30,142,29,142,28,141,31,155,31,41,31,145,31,220,31,221,31,86,31,247,31,162,31,226,31,147,31,230,31,64,31,64,30,64,29,129,31,196,31,196,30,100,31,100,30,36,31,36,30,88,31,1,31,1,30,156,31,171,31,201,31,121,31,64,31,171,31,153,31,184,31,89,31,202,31,67,31,193,31,52,31,196,31,127,31,231,31,92,31,122,31,37,31,247,31,184,31,126,31,126,30,241,31,157,31,124,31,221,31,157,31,67,31,67,30,204,31,106,31,106,30,38,31,170,31,117,31,1,31,63,31,231,31,97,31,100,31,100,30,165,31,66,31,44,31,81,31,8,31,8,30,25,31,247,31,113,31,251,31,7,31,182,31,182,30,165,31,192,31,251,31,67,31,153,31,233,31,47,31,19,31,28,31,102,31,239,31,182,31,182,30,32,31,225,31,17,31,4,31,218,31,238,31,17,31,99,31,210,31,129,31,9,31,83,31,83,30,152,31,56,31,24,31,121,31,115,31,251,31,247,31,57,31,57,30,29,31,191,31,110,31,219,31,145,31,6,31,6,30,51,31,73,31,100,31,100,30,100,29,245,31,152,31,122,31,57,31,76,31,191,31,55,31,58,31,39,31,24,31,74,31,187,31,229,31,113,31,113,30,111,31,3,31,40,31,109,31,67,31,167,31,81,31,172,31,231,31,246,31,246,30,246,29,76,31,11,31,11,30,155,31,68,31,112,31,68,31,55,31,152,31,219,31,219,30,219,29,54,31,2,31,2,30,171,31,171,30,255,31,194,31,57,31,235,31,97,31,213,31,213,30,213,29,213,28,4,31,193,31,21,31,21,30,21,29,77,31,82,31,82,30,205,31,77,31,77,30,77,29,200,31,30,31,30,30,30,29,255,31,209,31,247,31,244,31,49,31,147,31,167,31,167,30,167,29,231,31,231,30,38,31,189,31,36,31,40,31,145,31,205,31,96,31,96,30,14,31,243,31,62,31,62,30,62,29,102,31,162,31,55,31,209,31,209,30,2,31,220,31,114,31,114,30,114,29,211,31,204,31,60,31,227,31,188,31,31,31,85,31,55,31,97,31,245,31,187,31,5,31,163,31,155,31,176,31,176,30,235,31,235,30,90,31,217,31,146,31,122,31,127,31,156,31,184,31,53,31,160,31,172,31,56,31,56,30,247,31,7,31,7,30,167,31,117,31,94,31,62,31,26,31,244,31,96,31,62,31,62,30,146,31,43,31,214,31,37,31,42,31,243,31,224,31,208,31,208,30,221,31,163,31,189,31,13,31,228,31,69,31,69,30,253,31,253,30,140,31,63,31,208,31,208,30,208,29,227,31,54,31,54,30,211,31,25,31,160,31,76,31,87,31,88,31,21,31,252,31,166,31,176,31,176,30,176,29,43,31,3,31,2,31,206,31,206,30,123,31,140,31,54,31,11,31,131,31,131,30,57,31,118,31,118,30,118,29,100,31,53,31,242,31,177,31,177,30,129,31,2,31,2,30,145,31,139,31,123,31,248,31,72,31,26,31,99,31,227,31,227,30,227,29,236,31,236,30,236,29,236,28,41,31,8,31,183,31,65,31,79,31,79,30,229,31,175,31,105,31,195,31,91,31,141,31,132,31,132,30,84,31,84,30,78,31,78,30,229,31,229,30,13,31,53,31,45,31,6,31,6,30,115,31,114,31,105,31,48,31,28,31,225,31,102,31,92,31,209,31,6,31,118,31,231,31,231,30,131,31,43,31,43,30,42,31,9,31,68,31,64,31,84,31,193,31,193,30,108,31,108,30,68,31,178,31,178,30,34,31,217,31,234,31,255,31,79,31,79,30,170,31,113,31,73,31,152,31,60,31,12,31,30,31,135,31,34,31,161,31,132,31,29,31,75,31,112,31,112,30,121,31,102,31,102,30,229,31,57,31,229,31,92,31,92,30,121,31,197,31,5,31,26,31,26,30,140,31,140,30,50,31,48,31,74,31,168,31,168,30,232,31,49,31,187,31,18,31,32,31,3,31,137,31,153,31,153,30,14,31,14,30,14,29,14,28,14,27,14,26,219,31,196,31,68,31,226,31,202,31,202,30,202,29,202,28);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
