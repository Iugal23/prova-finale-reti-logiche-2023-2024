-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_648 is
end project_tb_648;

architecture project_tb_arch_648 of project_tb_648 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 157;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (216,0,122,0,61,0,0,0,206,0,144,0,152,0,15,0,0,0,39,0,209,0,0,0,72,0,14,0,252,0,118,0,63,0,139,0,230,0,72,0,37,0,37,0,43,0,206,0,204,0,0,0,148,0,202,0,230,0,232,0,18,0,0,0,21,0,123,0,152,0,250,0,237,0,4,0,126,0,48,0,104,0,160,0,25,0,111,0,181,0,181,0,77,0,25,0,171,0,182,0,217,0,252,0,168,0,110,0,149,0,107,0,180,0,0,0,49,0,245,0,0,0,0,0,107,0,138,0,170,0,167,0,16,0,173,0,127,0,245,0,138,0,0,0,38,0,69,0,219,0,170,0,80,0,50,0,78,0,225,0,235,0,162,0,203,0,2,0,2,0,0,0,46,0,41,0,217,0,194,0,149,0,215,0,229,0,0,0,8,0,151,0,0,0,127,0,49,0,223,0,116,0,141,0,28,0,127,0,241,0,254,0,122,0,122,0,0,0,0,0,213,0,0,0,122,0,146,0,0,0,0,0,120,0,0,0,74,0,168,0,199,0,189,0,49,0,205,0,227,0,217,0,118,0,0,0,172,0,64,0,185,0,212,0,253,0,214,0,95,0,21,0,206,0,0,0,0,0,0,0,0,0,0,0,157,0,18,0,44,0,167,0,22,0,16,0,0,0,64,0,72,0,38,0,0,0,101,0,135,0,143,0,21,0);
signal scenario_full  : scenario_type := (216,31,122,31,61,31,61,30,206,31,144,31,152,31,15,31,15,30,39,31,209,31,209,30,72,31,14,31,252,31,118,31,63,31,139,31,230,31,72,31,37,31,37,31,43,31,206,31,204,31,204,30,148,31,202,31,230,31,232,31,18,31,18,30,21,31,123,31,152,31,250,31,237,31,4,31,126,31,48,31,104,31,160,31,25,31,111,31,181,31,181,31,77,31,25,31,171,31,182,31,217,31,252,31,168,31,110,31,149,31,107,31,180,31,180,30,49,31,245,31,245,30,245,29,107,31,138,31,170,31,167,31,16,31,173,31,127,31,245,31,138,31,138,30,38,31,69,31,219,31,170,31,80,31,50,31,78,31,225,31,235,31,162,31,203,31,2,31,2,31,2,30,46,31,41,31,217,31,194,31,149,31,215,31,229,31,229,30,8,31,151,31,151,30,127,31,49,31,223,31,116,31,141,31,28,31,127,31,241,31,254,31,122,31,122,31,122,30,122,29,213,31,213,30,122,31,146,31,146,30,146,29,120,31,120,30,74,31,168,31,199,31,189,31,49,31,205,31,227,31,217,31,118,31,118,30,172,31,64,31,185,31,212,31,253,31,214,31,95,31,21,31,206,31,206,30,206,29,206,28,206,27,206,26,157,31,18,31,44,31,167,31,22,31,16,31,16,30,64,31,72,31,38,31,38,30,101,31,135,31,143,31,21,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
