-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_741 is
end project_tb_741;

architecture project_tb_arch_741 of project_tb_741 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 713;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (120,0,0,0,127,0,241,0,144,0,178,0,166,0,127,0,9,0,67,0,36,0,0,0,103,0,180,0,0,0,0,0,209,0,0,0,72,0,0,0,240,0,251,0,0,0,144,0,239,0,68,0,0,0,21,0,7,0,163,0,5,0,67,0,13,0,28,0,218,0,0,0,149,0,129,0,100,0,15,0,0,0,45,0,174,0,234,0,85,0,217,0,188,0,61,0,0,0,104,0,178,0,18,0,0,0,109,0,54,0,163,0,248,0,121,0,6,0,164,0,11,0,199,0,0,0,132,0,164,0,81,0,20,0,9,0,149,0,84,0,164,0,128,0,124,0,113,0,0,0,65,0,10,0,142,0,58,0,2,0,0,0,51,0,243,0,177,0,81,0,217,0,221,0,251,0,55,0,123,0,234,0,241,0,61,0,29,0,89,0,0,0,218,0,126,0,171,0,95,0,41,0,0,0,53,0,65,0,137,0,0,0,120,0,115,0,246,0,70,0,192,0,94,0,0,0,89,0,188,0,140,0,47,0,0,0,201,0,78,0,114,0,17,0,233,0,216,0,0,0,0,0,77,0,75,0,106,0,130,0,252,0,32,0,34,0,235,0,21,0,0,0,39,0,0,0,111,0,31,0,248,0,66,0,176,0,0,0,87,0,117,0,103,0,59,0,217,0,195,0,0,0,7,0,139,0,105,0,3,0,55,0,193,0,0,0,65,0,152,0,6,0,0,0,16,0,150,0,122,0,22,0,0,0,142,0,171,0,191,0,95,0,222,0,26,0,130,0,0,0,15,0,154,0,102,0,41,0,45,0,209,0,0,0,232,0,112,0,34,0,0,0,14,0,0,0,170,0,190,0,232,0,212,0,231,0,2,0,1,0,73,0,76,0,81,0,126,0,0,0,127,0,0,0,0,0,26,0,38,0,231,0,123,0,43,0,100,0,0,0,206,0,188,0,220,0,168,0,72,0,140,0,153,0,162,0,0,0,124,0,218,0,237,0,254,0,232,0,177,0,0,0,81,0,3,0,222,0,0,0,208,0,142,0,222,0,43,0,50,0,199,0,175,0,0,0,49,0,212,0,210,0,134,0,202,0,98,0,48,0,243,0,255,0,0,0,0,0,66,0,0,0,48,0,234,0,177,0,207,0,0,0,87,0,166,0,158,0,198,0,153,0,216,0,63,0,18,0,39,0,0,0,172,0,0,0,0,0,0,0,169,0,2,0,234,0,10,0,0,0,239,0,5,0,42,0,120,0,220,0,124,0,218,0,75,0,172,0,188,0,0,0,211,0,97,0,221,0,94,0,88,0,113,0,0,0,234,0,0,0,146,0,36,0,124,0,194,0,0,0,0,0,173,0,67,0,42,0,78,0,225,0,0,0,0,0,0,0,0,0,136,0,249,0,0,0,0,0,29,0,241,0,148,0,44,0,122,0,148,0,9,0,212,0,121,0,0,0,169,0,0,0,174,0,45,0,35,0,6,0,179,0,0,0,109,0,148,0,164,0,71,0,211,0,170,0,190,0,106,0,200,0,30,0,0,0,148,0,127,0,0,0,202,0,39,0,0,0,122,0,84,0,0,0,108,0,16,0,0,0,229,0,0,0,93,0,0,0,35,0,0,0,76,0,0,0,9,0,127,0,95,0,13,0,225,0,0,0,220,0,179,0,5,0,249,0,47,0,174,0,70,0,201,0,144,0,56,0,217,0,150,0,0,0,137,0,75,0,194,0,0,0,215,0,0,0,16,0,137,0,27,0,74,0,246,0,250,0,0,0,0,0,0,0,171,0,0,0,209,0,140,0,220,0,0,0,108,0,25,0,144,0,33,0,143,0,67,0,0,0,244,0,0,0,102,0,132,0,0,0,73,0,91,0,189,0,254,0,0,0,88,0,0,0,33,0,15,0,212,0,237,0,0,0,73,0,118,0,66,0,233,0,157,0,3,0,162,0,153,0,0,0,145,0,226,0,0,0,0,0,0,0,0,0,0,0,0,0,72,0,0,0,0,0,0,0,240,0,11,0,96,0,235,0,225,0,0,0,206,0,0,0,139,0,171,0,105,0,228,0,43,0,0,0,152,0,232,0,121,0,193,0,0,0,24,0,0,0,58,0,58,0,214,0,153,0,139,0,207,0,248,0,148,0,143,0,114,0,199,0,159,0,255,0,143,0,134,0,253,0,184,0,146,0,200,0,208,0,0,0,211,0,0,0,95,0,141,0,196,0,221,0,208,0,125,0,237,0,0,0,185,0,0,0,174,0,34,0,214,0,94,0,227,0,0,0,218,0,172,0,0,0,0,0,42,0,94,0,9,0,0,0,149,0,188,0,85,0,0,0,112,0,213,0,0,0,0,0,0,0,166,0,118,0,231,0,20,0,81,0,14,0,144,0,20,0,237,0,130,0,229,0,0,0,65,0,170,0,0,0,146,0,254,0,205,0,119,0,150,0,1,0,248,0,175,0,151,0,184,0,144,0,60,0,210,0,149,0,75,0,69,0,195,0,206,0,234,0,119,0,26,0,47,0,0,0,0,0,45,0,234,0,156,0,121,0,214,0,8,0,225,0,55,0,175,0,24,0,208,0,16,0,250,0,0,0,62,0,227,0,238,0,113,0,136,0,127,0,18,0,0,0,89,0,158,0,227,0,38,0,129,0,114,0,160,0,248,0,0,0,89,0,226,0,127,0,96,0,209,0,154,0,190,0,2,0,245,0,23,0,241,0,243,0,132,0,237,0,0,0,0,0,134,0,31,0,0,0,96,0,173,0,6,0,160,0,245,0,194,0,122,0,0,0,0,0,34,0,71,0,102,0,81,0,232,0,172,0,211,0,250,0,0,0,0,0,161,0,0,0,156,0,180,0,233,0,40,0,111,0,229,0,101,0,223,0,30,0,219,0,116,0,197,0,0,0,250,0,101,0,17,0,27,0,0,0,14,0,156,0,88,0,161,0,77,0,162,0,116,0,31,0,146,0,107,0,100,0,183,0,77,0,0,0,59,0,132,0,156,0,99,0,0,0,187,0,52,0,0,0,0,0,0,0,240,0,0,0,159,0,226,0,0,0,182,0,0,0,161,0,0,0,210,0,126,0,110,0,161,0,25,0,0,0,21,0,136,0,40,0,0,0,146,0,138,0,62,0,74,0,175,0,226,0,0,0,43,0,118,0,39,0,186,0,0,0,20,0,120,0,0,0,20,0,123,0);
signal scenario_full  : scenario_type := (120,31,120,30,127,31,241,31,144,31,178,31,166,31,127,31,9,31,67,31,36,31,36,30,103,31,180,31,180,30,180,29,209,31,209,30,72,31,72,30,240,31,251,31,251,30,144,31,239,31,68,31,68,30,21,31,7,31,163,31,5,31,67,31,13,31,28,31,218,31,218,30,149,31,129,31,100,31,15,31,15,30,45,31,174,31,234,31,85,31,217,31,188,31,61,31,61,30,104,31,178,31,18,31,18,30,109,31,54,31,163,31,248,31,121,31,6,31,164,31,11,31,199,31,199,30,132,31,164,31,81,31,20,31,9,31,149,31,84,31,164,31,128,31,124,31,113,31,113,30,65,31,10,31,142,31,58,31,2,31,2,30,51,31,243,31,177,31,81,31,217,31,221,31,251,31,55,31,123,31,234,31,241,31,61,31,29,31,89,31,89,30,218,31,126,31,171,31,95,31,41,31,41,30,53,31,65,31,137,31,137,30,120,31,115,31,246,31,70,31,192,31,94,31,94,30,89,31,188,31,140,31,47,31,47,30,201,31,78,31,114,31,17,31,233,31,216,31,216,30,216,29,77,31,75,31,106,31,130,31,252,31,32,31,34,31,235,31,21,31,21,30,39,31,39,30,111,31,31,31,248,31,66,31,176,31,176,30,87,31,117,31,103,31,59,31,217,31,195,31,195,30,7,31,139,31,105,31,3,31,55,31,193,31,193,30,65,31,152,31,6,31,6,30,16,31,150,31,122,31,22,31,22,30,142,31,171,31,191,31,95,31,222,31,26,31,130,31,130,30,15,31,154,31,102,31,41,31,45,31,209,31,209,30,232,31,112,31,34,31,34,30,14,31,14,30,170,31,190,31,232,31,212,31,231,31,2,31,1,31,73,31,76,31,81,31,126,31,126,30,127,31,127,30,127,29,26,31,38,31,231,31,123,31,43,31,100,31,100,30,206,31,188,31,220,31,168,31,72,31,140,31,153,31,162,31,162,30,124,31,218,31,237,31,254,31,232,31,177,31,177,30,81,31,3,31,222,31,222,30,208,31,142,31,222,31,43,31,50,31,199,31,175,31,175,30,49,31,212,31,210,31,134,31,202,31,98,31,48,31,243,31,255,31,255,30,255,29,66,31,66,30,48,31,234,31,177,31,207,31,207,30,87,31,166,31,158,31,198,31,153,31,216,31,63,31,18,31,39,31,39,30,172,31,172,30,172,29,172,28,169,31,2,31,234,31,10,31,10,30,239,31,5,31,42,31,120,31,220,31,124,31,218,31,75,31,172,31,188,31,188,30,211,31,97,31,221,31,94,31,88,31,113,31,113,30,234,31,234,30,146,31,36,31,124,31,194,31,194,30,194,29,173,31,67,31,42,31,78,31,225,31,225,30,225,29,225,28,225,27,136,31,249,31,249,30,249,29,29,31,241,31,148,31,44,31,122,31,148,31,9,31,212,31,121,31,121,30,169,31,169,30,174,31,45,31,35,31,6,31,179,31,179,30,109,31,148,31,164,31,71,31,211,31,170,31,190,31,106,31,200,31,30,31,30,30,148,31,127,31,127,30,202,31,39,31,39,30,122,31,84,31,84,30,108,31,16,31,16,30,229,31,229,30,93,31,93,30,35,31,35,30,76,31,76,30,9,31,127,31,95,31,13,31,225,31,225,30,220,31,179,31,5,31,249,31,47,31,174,31,70,31,201,31,144,31,56,31,217,31,150,31,150,30,137,31,75,31,194,31,194,30,215,31,215,30,16,31,137,31,27,31,74,31,246,31,250,31,250,30,250,29,250,28,171,31,171,30,209,31,140,31,220,31,220,30,108,31,25,31,144,31,33,31,143,31,67,31,67,30,244,31,244,30,102,31,132,31,132,30,73,31,91,31,189,31,254,31,254,30,88,31,88,30,33,31,15,31,212,31,237,31,237,30,73,31,118,31,66,31,233,31,157,31,3,31,162,31,153,31,153,30,145,31,226,31,226,30,226,29,226,28,226,27,226,26,226,25,72,31,72,30,72,29,72,28,240,31,11,31,96,31,235,31,225,31,225,30,206,31,206,30,139,31,171,31,105,31,228,31,43,31,43,30,152,31,232,31,121,31,193,31,193,30,24,31,24,30,58,31,58,31,214,31,153,31,139,31,207,31,248,31,148,31,143,31,114,31,199,31,159,31,255,31,143,31,134,31,253,31,184,31,146,31,200,31,208,31,208,30,211,31,211,30,95,31,141,31,196,31,221,31,208,31,125,31,237,31,237,30,185,31,185,30,174,31,34,31,214,31,94,31,227,31,227,30,218,31,172,31,172,30,172,29,42,31,94,31,9,31,9,30,149,31,188,31,85,31,85,30,112,31,213,31,213,30,213,29,213,28,166,31,118,31,231,31,20,31,81,31,14,31,144,31,20,31,237,31,130,31,229,31,229,30,65,31,170,31,170,30,146,31,254,31,205,31,119,31,150,31,1,31,248,31,175,31,151,31,184,31,144,31,60,31,210,31,149,31,75,31,69,31,195,31,206,31,234,31,119,31,26,31,47,31,47,30,47,29,45,31,234,31,156,31,121,31,214,31,8,31,225,31,55,31,175,31,24,31,208,31,16,31,250,31,250,30,62,31,227,31,238,31,113,31,136,31,127,31,18,31,18,30,89,31,158,31,227,31,38,31,129,31,114,31,160,31,248,31,248,30,89,31,226,31,127,31,96,31,209,31,154,31,190,31,2,31,245,31,23,31,241,31,243,31,132,31,237,31,237,30,237,29,134,31,31,31,31,30,96,31,173,31,6,31,160,31,245,31,194,31,122,31,122,30,122,29,34,31,71,31,102,31,81,31,232,31,172,31,211,31,250,31,250,30,250,29,161,31,161,30,156,31,180,31,233,31,40,31,111,31,229,31,101,31,223,31,30,31,219,31,116,31,197,31,197,30,250,31,101,31,17,31,27,31,27,30,14,31,156,31,88,31,161,31,77,31,162,31,116,31,31,31,146,31,107,31,100,31,183,31,77,31,77,30,59,31,132,31,156,31,99,31,99,30,187,31,52,31,52,30,52,29,52,28,240,31,240,30,159,31,226,31,226,30,182,31,182,30,161,31,161,30,210,31,126,31,110,31,161,31,25,31,25,30,21,31,136,31,40,31,40,30,146,31,138,31,62,31,74,31,175,31,226,31,226,30,43,31,118,31,39,31,186,31,186,30,20,31,120,31,120,30,20,31,123,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
