-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_593 is
end project_tb_593;

architecture project_tb_arch_593 of project_tb_593 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 904;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (183,0,245,0,13,0,37,0,215,0,143,0,243,0,83,0,87,0,221,0,107,0,0,0,146,0,173,0,24,0,81,0,104,0,75,0,134,0,238,0,233,0,37,0,84,0,0,0,0,0,221,0,0,0,7,0,0,0,227,0,139,0,70,0,250,0,70,0,14,0,0,0,166,0,152,0,185,0,255,0,0,0,0,0,88,0,22,0,76,0,0,0,167,0,78,0,249,0,55,0,61,0,209,0,235,0,151,0,153,0,0,0,241,0,11,0,0,0,233,0,200,0,24,0,166,0,91,0,0,0,171,0,254,0,0,0,124,0,0,0,124,0,0,0,168,0,0,0,39,0,155,0,160,0,184,0,134,0,80,0,0,0,0,0,0,0,220,0,28,0,146,0,0,0,152,0,64,0,0,0,29,0,210,0,189,0,215,0,118,0,195,0,12,0,0,0,84,0,94,0,136,0,170,0,248,0,155,0,249,0,190,0,225,0,0,0,131,0,108,0,172,0,218,0,0,0,96,0,56,0,163,0,161,0,98,0,0,0,0,0,0,0,95,0,72,0,238,0,124,0,238,0,143,0,244,0,134,0,187,0,0,0,144,0,183,0,0,0,0,0,73,0,200,0,49,0,120,0,100,0,26,0,0,0,0,0,141,0,139,0,177,0,119,0,27,0,255,0,198,0,203,0,246,0,0,0,0,0,144,0,190,0,103,0,237,0,207,0,176,0,252,0,234,0,255,0,152,0,0,0,9,0,25,0,42,0,177,0,160,0,54,0,220,0,190,0,145,0,213,0,113,0,0,0,136,0,236,0,65,0,0,0,119,0,0,0,112,0,155,0,11,0,70,0,58,0,98,0,0,0,67,0,8,0,190,0,231,0,242,0,210,0,223,0,215,0,47,0,0,0,11,0,230,0,0,0,49,0,170,0,14,0,26,0,75,0,91,0,61,0,247,0,244,0,128,0,111,0,193,0,0,0,9,0,22,0,81,0,52,0,219,0,250,0,127,0,14,0,0,0,190,0,179,0,152,0,0,0,227,0,174,0,0,0,52,0,57,0,106,0,0,0,188,0,7,0,96,0,19,0,0,0,124,0,213,0,1,0,255,0,251,0,96,0,197,0,0,0,186,0,72,0,0,0,178,0,208,0,47,0,131,0,0,0,156,0,227,0,0,0,109,0,174,0,236,0,0,0,130,0,22,0,253,0,95,0,27,0,242,0,163,0,208,0,0,0,90,0,149,0,233,0,228,0,0,0,114,0,90,0,125,0,163,0,189,0,225,0,84,0,0,0,148,0,82,0,242,0,0,0,69,0,37,0,192,0,120,0,205,0,0,0,78,0,191,0,0,0,244,0,111,0,69,0,238,0,128,0,0,0,121,0,70,0,232,0,74,0,0,0,0,0,0,0,249,0,4,0,193,0,115,0,0,0,177,0,0,0,222,0,0,0,30,0,32,0,0,0,35,0,217,0,70,0,154,0,117,0,0,0,183,0,130,0,87,0,0,0,162,0,167,0,7,0,135,0,0,0,0,0,211,0,67,0,0,0,0,0,0,0,248,0,0,0,1,0,53,0,80,0,118,0,147,0,15,0,238,0,19,0,0,0,149,0,96,0,0,0,0,0,85,0,0,0,31,0,97,0,229,0,137,0,18,0,164,0,119,0,81,0,123,0,160,0,188,0,127,0,127,0,255,0,18,0,0,0,192,0,19,0,238,0,222,0,53,0,6,0,0,0,200,0,199,0,172,0,82,0,212,0,156,0,55,0,234,0,26,0,93,0,60,0,45,0,219,0,66,0,59,0,145,0,8,0,194,0,0,0,109,0,18,0,153,0,254,0,214,0,81,0,205,0,153,0,36,0,123,0,0,0,0,0,99,0,156,0,249,0,2,0,0,0,0,0,0,0,134,0,207,0,0,0,162,0,153,0,149,0,139,0,7,0,190,0,252,0,201,0,68,0,0,0,0,0,21,0,0,0,11,0,48,0,227,0,45,0,229,0,103,0,151,0,86,0,33,0,201,0,0,0,221,0,120,0,0,0,173,0,78,0,17,0,62,0,45,0,96,0,162,0,146,0,0,0,0,0,147,0,52,0,45,0,152,0,15,0,102,0,0,0,2,0,219,0,21,0,234,0,195,0,196,0,182,0,114,0,0,0,109,0,117,0,171,0,0,0,152,0,185,0,222,0,87,0,191,0,103,0,0,0,178,0,0,0,141,0,46,0,231,0,12,0,128,0,0,0,166,0,226,0,137,0,121,0,0,0,242,0,110,0,8,0,248,0,5,0,96,0,148,0,11,0,239,0,171,0,0,0,5,0,101,0,33,0,106,0,118,0,70,0,65,0,4,0,0,0,78,0,125,0,191,0,127,0,158,0,61,0,199,0,31,0,25,0,0,0,114,0,164,0,0,0,193,0,0,0,16,0,247,0,193,0,133,0,116,0,102,0,35,0,47,0,0,0,153,0,0,0,213,0,163,0,204,0,229,0,46,0,3,0,31,0,128,0,133,0,192,0,78,0,193,0,97,0,109,0,100,0,80,0,118,0,67,0,80,0,0,0,48,0,160,0,172,0,166,0,0,0,0,0,138,0,142,0,0,0,0,0,120,0,9,0,90,0,0,0,24,0,0,0,224,0,0,0,161,0,0,0,9,0,2,0,200,0,0,0,132,0,118,0,0,0,24,0,0,0,0,0,36,0,66,0,0,0,131,0,49,0,57,0,115,0,0,0,0,0,3,0,206,0,172,0,175,0,177,0,92,0,180,0,161,0,157,0,168,0,24,0,13,0,163,0,219,0,132,0,251,0,0,0,232,0,79,0,102,0,42,0,164,0,162,0,80,0,7,0,0,0,0,0,139,0,12,0,155,0,0,0,0,0,157,0,160,0,187,0,136,0,239,0,197,0,23,0,237,0,120,0,111,0,13,0,0,0,0,0,0,0,138,0,88,0,75,0,42,0,165,0,46,0,96,0,139,0,0,0,26,0,194,0,204,0,228,0,133,0,115,0,0,0,86,0,196,0,151,0,90,0,178,0,125,0,167,0,88,0,228,0,0,0,80,0,166,0,207,0,0,0,12,0,81,0,0,0,0,0,181,0,231,0,0,0,114,0,101,0,161,0,35,0,0,0,86,0,80,0,0,0,68,0,0,0,13,0,0,0,204,0,0,0,104,0,0,0,106,0,156,0,250,0,143,0,0,0,49,0,0,0,0,0,59,0,131,0,0,0,247,0,55,0,211,0,132,0,202,0,25,0,108,0,6,0,17,0,103,0,225,0,28,0,0,0,0,0,203,0,247,0,0,0,211,0,219,0,240,0,49,0,247,0,231,0,237,0,23,0,153,0,254,0,230,0,240,0,177,0,147,0,143,0,37,0,215,0,0,0,231,0,22,0,83,0,93,0,193,0,204,0,0,0,116,0,130,0,93,0,129,0,11,0,218,0,0,0,0,0,99,0,127,0,43,0,150,0,244,0,224,0,244,0,177,0,178,0,0,0,219,0,155,0,183,0,194,0,239,0,145,0,20,0,0,0,71,0,200,0,0,0,240,0,52,0,233,0,202,0,173,0,38,0,135,0,199,0,94,0,230,0,83,0,107,0,109,0,150,0,0,0,104,0,134,0,196,0,0,0,122,0,232,0,45,0,58,0,0,0,0,0,170,0,181,0,0,0,150,0,0,0,38,0,237,0,244,0,0,0,43,0,42,0,40,0,33,0,115,0,223,0,78,0,195,0,135,0,104,0,23,0,205,0,195,0,199,0,160,0,30,0,0,0,58,0,201,0,130,0,0,0,43,0,137,0,254,0,137,0,0,0,242,0,216,0,255,0,219,0,0,0,253,0,62,0,0,0,39,0,0,0,252,0,127,0,127,0,244,0,156,0,43,0,121,0,120,0,26,0,1,0,176,0,140,0,252,0,105,0,143,0,222,0,149,0,221,0,13,0,80,0,245,0,243,0,0,0,0,0,125,0,51,0,5,0,200,0,159,0,236,0,94,0,71,0,9,0,0,0,11,0,41,0,57,0,3,0,98,0,140,0,67,0,189,0,210,0,0,0,109,0);
signal scenario_full  : scenario_type := (183,31,245,31,13,31,37,31,215,31,143,31,243,31,83,31,87,31,221,31,107,31,107,30,146,31,173,31,24,31,81,31,104,31,75,31,134,31,238,31,233,31,37,31,84,31,84,30,84,29,221,31,221,30,7,31,7,30,227,31,139,31,70,31,250,31,70,31,14,31,14,30,166,31,152,31,185,31,255,31,255,30,255,29,88,31,22,31,76,31,76,30,167,31,78,31,249,31,55,31,61,31,209,31,235,31,151,31,153,31,153,30,241,31,11,31,11,30,233,31,200,31,24,31,166,31,91,31,91,30,171,31,254,31,254,30,124,31,124,30,124,31,124,30,168,31,168,30,39,31,155,31,160,31,184,31,134,31,80,31,80,30,80,29,80,28,220,31,28,31,146,31,146,30,152,31,64,31,64,30,29,31,210,31,189,31,215,31,118,31,195,31,12,31,12,30,84,31,94,31,136,31,170,31,248,31,155,31,249,31,190,31,225,31,225,30,131,31,108,31,172,31,218,31,218,30,96,31,56,31,163,31,161,31,98,31,98,30,98,29,98,28,95,31,72,31,238,31,124,31,238,31,143,31,244,31,134,31,187,31,187,30,144,31,183,31,183,30,183,29,73,31,200,31,49,31,120,31,100,31,26,31,26,30,26,29,141,31,139,31,177,31,119,31,27,31,255,31,198,31,203,31,246,31,246,30,246,29,144,31,190,31,103,31,237,31,207,31,176,31,252,31,234,31,255,31,152,31,152,30,9,31,25,31,42,31,177,31,160,31,54,31,220,31,190,31,145,31,213,31,113,31,113,30,136,31,236,31,65,31,65,30,119,31,119,30,112,31,155,31,11,31,70,31,58,31,98,31,98,30,67,31,8,31,190,31,231,31,242,31,210,31,223,31,215,31,47,31,47,30,11,31,230,31,230,30,49,31,170,31,14,31,26,31,75,31,91,31,61,31,247,31,244,31,128,31,111,31,193,31,193,30,9,31,22,31,81,31,52,31,219,31,250,31,127,31,14,31,14,30,190,31,179,31,152,31,152,30,227,31,174,31,174,30,52,31,57,31,106,31,106,30,188,31,7,31,96,31,19,31,19,30,124,31,213,31,1,31,255,31,251,31,96,31,197,31,197,30,186,31,72,31,72,30,178,31,208,31,47,31,131,31,131,30,156,31,227,31,227,30,109,31,174,31,236,31,236,30,130,31,22,31,253,31,95,31,27,31,242,31,163,31,208,31,208,30,90,31,149,31,233,31,228,31,228,30,114,31,90,31,125,31,163,31,189,31,225,31,84,31,84,30,148,31,82,31,242,31,242,30,69,31,37,31,192,31,120,31,205,31,205,30,78,31,191,31,191,30,244,31,111,31,69,31,238,31,128,31,128,30,121,31,70,31,232,31,74,31,74,30,74,29,74,28,249,31,4,31,193,31,115,31,115,30,177,31,177,30,222,31,222,30,30,31,32,31,32,30,35,31,217,31,70,31,154,31,117,31,117,30,183,31,130,31,87,31,87,30,162,31,167,31,7,31,135,31,135,30,135,29,211,31,67,31,67,30,67,29,67,28,248,31,248,30,1,31,53,31,80,31,118,31,147,31,15,31,238,31,19,31,19,30,149,31,96,31,96,30,96,29,85,31,85,30,31,31,97,31,229,31,137,31,18,31,164,31,119,31,81,31,123,31,160,31,188,31,127,31,127,31,255,31,18,31,18,30,192,31,19,31,238,31,222,31,53,31,6,31,6,30,200,31,199,31,172,31,82,31,212,31,156,31,55,31,234,31,26,31,93,31,60,31,45,31,219,31,66,31,59,31,145,31,8,31,194,31,194,30,109,31,18,31,153,31,254,31,214,31,81,31,205,31,153,31,36,31,123,31,123,30,123,29,99,31,156,31,249,31,2,31,2,30,2,29,2,28,134,31,207,31,207,30,162,31,153,31,149,31,139,31,7,31,190,31,252,31,201,31,68,31,68,30,68,29,21,31,21,30,11,31,48,31,227,31,45,31,229,31,103,31,151,31,86,31,33,31,201,31,201,30,221,31,120,31,120,30,173,31,78,31,17,31,62,31,45,31,96,31,162,31,146,31,146,30,146,29,147,31,52,31,45,31,152,31,15,31,102,31,102,30,2,31,219,31,21,31,234,31,195,31,196,31,182,31,114,31,114,30,109,31,117,31,171,31,171,30,152,31,185,31,222,31,87,31,191,31,103,31,103,30,178,31,178,30,141,31,46,31,231,31,12,31,128,31,128,30,166,31,226,31,137,31,121,31,121,30,242,31,110,31,8,31,248,31,5,31,96,31,148,31,11,31,239,31,171,31,171,30,5,31,101,31,33,31,106,31,118,31,70,31,65,31,4,31,4,30,78,31,125,31,191,31,127,31,158,31,61,31,199,31,31,31,25,31,25,30,114,31,164,31,164,30,193,31,193,30,16,31,247,31,193,31,133,31,116,31,102,31,35,31,47,31,47,30,153,31,153,30,213,31,163,31,204,31,229,31,46,31,3,31,31,31,128,31,133,31,192,31,78,31,193,31,97,31,109,31,100,31,80,31,118,31,67,31,80,31,80,30,48,31,160,31,172,31,166,31,166,30,166,29,138,31,142,31,142,30,142,29,120,31,9,31,90,31,90,30,24,31,24,30,224,31,224,30,161,31,161,30,9,31,2,31,200,31,200,30,132,31,118,31,118,30,24,31,24,30,24,29,36,31,66,31,66,30,131,31,49,31,57,31,115,31,115,30,115,29,3,31,206,31,172,31,175,31,177,31,92,31,180,31,161,31,157,31,168,31,24,31,13,31,163,31,219,31,132,31,251,31,251,30,232,31,79,31,102,31,42,31,164,31,162,31,80,31,7,31,7,30,7,29,139,31,12,31,155,31,155,30,155,29,157,31,160,31,187,31,136,31,239,31,197,31,23,31,237,31,120,31,111,31,13,31,13,30,13,29,13,28,138,31,88,31,75,31,42,31,165,31,46,31,96,31,139,31,139,30,26,31,194,31,204,31,228,31,133,31,115,31,115,30,86,31,196,31,151,31,90,31,178,31,125,31,167,31,88,31,228,31,228,30,80,31,166,31,207,31,207,30,12,31,81,31,81,30,81,29,181,31,231,31,231,30,114,31,101,31,161,31,35,31,35,30,86,31,80,31,80,30,68,31,68,30,13,31,13,30,204,31,204,30,104,31,104,30,106,31,156,31,250,31,143,31,143,30,49,31,49,30,49,29,59,31,131,31,131,30,247,31,55,31,211,31,132,31,202,31,25,31,108,31,6,31,17,31,103,31,225,31,28,31,28,30,28,29,203,31,247,31,247,30,211,31,219,31,240,31,49,31,247,31,231,31,237,31,23,31,153,31,254,31,230,31,240,31,177,31,147,31,143,31,37,31,215,31,215,30,231,31,22,31,83,31,93,31,193,31,204,31,204,30,116,31,130,31,93,31,129,31,11,31,218,31,218,30,218,29,99,31,127,31,43,31,150,31,244,31,224,31,244,31,177,31,178,31,178,30,219,31,155,31,183,31,194,31,239,31,145,31,20,31,20,30,71,31,200,31,200,30,240,31,52,31,233,31,202,31,173,31,38,31,135,31,199,31,94,31,230,31,83,31,107,31,109,31,150,31,150,30,104,31,134,31,196,31,196,30,122,31,232,31,45,31,58,31,58,30,58,29,170,31,181,31,181,30,150,31,150,30,38,31,237,31,244,31,244,30,43,31,42,31,40,31,33,31,115,31,223,31,78,31,195,31,135,31,104,31,23,31,205,31,195,31,199,31,160,31,30,31,30,30,58,31,201,31,130,31,130,30,43,31,137,31,254,31,137,31,137,30,242,31,216,31,255,31,219,31,219,30,253,31,62,31,62,30,39,31,39,30,252,31,127,31,127,31,244,31,156,31,43,31,121,31,120,31,26,31,1,31,176,31,140,31,252,31,105,31,143,31,222,31,149,31,221,31,13,31,80,31,245,31,243,31,243,30,243,29,125,31,51,31,5,31,200,31,159,31,236,31,94,31,71,31,9,31,9,30,11,31,41,31,57,31,3,31,98,31,140,31,67,31,189,31,210,31,210,30,109,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
