-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_719 is
end project_tb_719;

architecture project_tb_arch_719 of project_tb_719 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 865;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (115,0,247,0,146,0,0,0,176,0,50,0,129,0,134,0,253,0,11,0,10,0,0,0,172,0,7,0,109,0,14,0,154,0,121,0,131,0,47,0,142,0,0,0,133,0,201,0,192,0,0,0,0,0,252,0,19,0,33,0,154,0,221,0,2,0,201,0,0,0,73,0,75,0,164,0,229,0,68,0,213,0,58,0,224,0,136,0,0,0,159,0,13,0,133,0,45,0,193,0,69,0,172,0,54,0,11,0,0,0,206,0,0,0,103,0,0,0,0,0,77,0,0,0,68,0,0,0,252,0,207,0,241,0,112,0,92,0,72,0,199,0,140,0,222,0,55,0,236,0,136,0,167,0,208,0,0,0,223,0,151,0,24,0,4,0,157,0,0,0,180,0,0,0,0,0,195,0,53,0,184,0,149,0,0,0,109,0,85,0,27,0,142,0,214,0,0,0,118,0,0,0,0,0,168,0,0,0,58,0,39,0,5,0,232,0,231,0,115,0,86,0,112,0,106,0,249,0,0,0,0,0,62,0,78,0,104,0,238,0,0,0,133,0,186,0,108,0,124,0,0,0,125,0,198,0,252,0,32,0,0,0,0,0,88,0,0,0,153,0,234,0,27,0,27,0,181,0,153,0,118,0,240,0,179,0,5,0,0,0,200,0,137,0,0,0,23,0,82,0,145,0,39,0,212,0,135,0,0,0,8,0,134,0,12,0,153,0,102,0,134,0,202,0,245,0,0,0,0,0,213,0,0,0,141,0,190,0,137,0,0,0,204,0,253,0,0,0,159,0,179,0,135,0,163,0,0,0,94,0,124,0,126,0,98,0,181,0,53,0,152,0,57,0,141,0,83,0,189,0,118,0,193,0,55,0,0,0,0,0,0,0,106,0,12,0,72,0,127,0,68,0,7,0,173,0,29,0,0,0,14,0,171,0,208,0,211,0,137,0,0,0,203,0,51,0,240,0,234,0,186,0,0,0,159,0,142,0,0,0,12,0,78,0,133,0,0,0,175,0,39,0,32,0,124,0,0,0,129,0,189,0,176,0,0,0,0,0,7,0,58,0,0,0,236,0,35,0,191,0,231,0,58,0,98,0,0,0,33,0,0,0,184,0,0,0,28,0,0,0,37,0,114,0,119,0,154,0,105,0,0,0,203,0,41,0,55,0,234,0,0,0,103,0,135,0,166,0,138,0,0,0,50,0,0,0,93,0,118,0,169,0,212,0,29,0,0,0,75,0,0,0,0,0,191,0,92,0,200,0,216,0,232,0,98,0,101,0,30,0,63,0,170,0,208,0,144,0,0,0,7,0,107,0,0,0,213,0,68,0,237,0,222,0,96,0,85,0,207,0,79,0,120,0,46,0,72,0,164,0,0,0,51,0,77,0,0,0,107,0,93,0,72,0,196,0,183,0,106,0,148,0,234,0,173,0,53,0,201,0,212,0,146,0,0,0,52,0,69,0,188,0,68,0,0,0,255,0,103,0,86,0,148,0,109,0,71,0,167,0,97,0,176,0,24,0,0,0,203,0,144,0,0,0,110,0,23,0,160,0,0,0,50,0,171,0,158,0,208,0,248,0,155,0,171,0,0,0,79,0,155,0,30,0,103,0,0,0,201,0,156,0,84,0,83,0,208,0,202,0,31,0,222,0,0,0,214,0,0,0,44,0,216,0,0,0,58,0,75,0,55,0,127,0,219,0,161,0,48,0,202,0,123,0,162,0,187,0,143,0,0,0,168,0,158,0,62,0,89,0,188,0,121,0,0,0,0,0,131,0,0,0,30,0,127,0,0,0,52,0,95,0,76,0,0,0,0,0,200,0,0,0,51,0,0,0,199,0,164,0,120,0,14,0,52,0,4,0,163,0,207,0,116,0,145,0,0,0,12,0,210,0,0,0,95,0,163,0,184,0,0,0,146,0,156,0,140,0,146,0,96,0,121,0,188,0,18,0,170,0,0,0,5,0,0,0,0,0,211,0,30,0,136,0,55,0,0,0,51,0,204,0,132,0,255,0,48,0,97,0,0,0,197,0,18,0,57,0,117,0,23,0,53,0,111,0,0,0,159,0,198,0,23,0,181,0,55,0,0,0,116,0,31,0,246,0,178,0,0,0,124,0,13,0,124,0,155,0,22,0,18,0,0,0,188,0,178,0,11,0,9,0,118,0,223,0,132,0,29,0,11,0,236,0,75,0,4,0,0,0,187,0,28,0,12,0,0,0,0,0,0,0,73,0,174,0,118,0,215,0,14,0,3,0,86,0,159,0,34,0,169,0,73,0,61,0,235,0,200,0,0,0,248,0,248,0,101,0,0,0,239,0,223,0,50,0,102,0,216,0,88,0,162,0,111,0,118,0,90,0,63,0,177,0,0,0,2,0,85,0,102,0,82,0,0,0,216,0,50,0,50,0,142,0,48,0,156,0,206,0,165,0,114,0,246,0,57,0,215,0,201,0,1,0,75,0,213,0,106,0,191,0,144,0,102,0,110,0,30,0,65,0,113,0,0,0,0,0,157,0,145,0,239,0,191,0,99,0,160,0,0,0,0,0,0,0,211,0,129,0,97,0,207,0,212,0,228,0,86,0,18,0,132,0,195,0,0,0,194,0,121,0,76,0,9,0,79,0,10,0,194,0,93,0,11,0,95,0,82,0,31,0,244,0,7,0,250,0,0,0,130,0,130,0,207,0,0,0,253,0,89,0,25,0,0,0,58,0,46,0,75,0,149,0,153,0,52,0,26,0,17,0,202,0,181,0,0,0,54,0,0,0,239,0,73,0,192,0,118,0,0,0,0,0,0,0,162,0,156,0,0,0,77,0,0,0,56,0,55,0,192,0,114,0,0,0,23,0,0,0,92,0,176,0,0,0,187,0,20,0,186,0,0,0,132,0,232,0,247,0,0,0,30,0,0,0,162,0,48,0,195,0,87,0,252,0,126,0,236,0,136,0,0,0,0,0,0,0,0,0,167,0,219,0,159,0,197,0,131,0,255,0,0,0,10,0,209,0,198,0,179,0,247,0,118,0,195,0,117,0,61,0,23,0,154,0,117,0,0,0,128,0,49,0,52,0,0,0,0,0,0,0,73,0,220,0,34,0,0,0,0,0,93,0,214,0,242,0,184,0,61,0,192,0,137,0,0,0,45,0,43,0,186,0,146,0,48,0,158,0,139,0,157,0,130,0,225,0,181,0,237,0,180,0,0,0,15,0,227,0,133,0,154,0,105,0,236,0,127,0,245,0,144,0,218,0,248,0,223,0,0,0,79,0,232,0,131,0,166,0,163,0,251,0,133,0,242,0,114,0,238,0,148,0,177,0,33,0,220,0,50,0,60,0,156,0,42,0,147,0,209,0,150,0,55,0,0,0,254,0,78,0,118,0,0,0,211,0,0,0,13,0,174,0,88,0,218,0,0,0,0,0,234,0,53,0,234,0,0,0,221,0,66,0,89,0,2,0,185,0,0,0,189,0,198,0,104,0,57,0,92,0,226,0,235,0,0,0,223,0,166,0,241,0,0,0,175,0,252,0,0,0,220,0,221,0,155,0,215,0,136,0,47,0,179,0,39,0,178,0,119,0,0,0,227,0,96,0,51,0,247,0,114,0,166,0,238,0,226,0,57,0,143,0,0,0,49,0,187,0,86,0,0,0,0,0,132,0,59,0,0,0,0,0,111,0,206,0,204,0,118,0,232,0,89,0,0,0,216,0,0,0,130,0,217,0,0,0,103,0,156,0,187,0,148,0,242,0,120,0,180,0,249,0,0,0,105,0,109,0,200,0,83,0,231,0,68,0,115,0,229,0,228,0,34,0,55,0,0,0,156,0,131,0,109,0,32,0,19,0,0,0,18,0,224,0,22,0,0,0,86,0,0,0,138,0,223,0,74,0);
signal scenario_full  : scenario_type := (115,31,247,31,146,31,146,30,176,31,50,31,129,31,134,31,253,31,11,31,10,31,10,30,172,31,7,31,109,31,14,31,154,31,121,31,131,31,47,31,142,31,142,30,133,31,201,31,192,31,192,30,192,29,252,31,19,31,33,31,154,31,221,31,2,31,201,31,201,30,73,31,75,31,164,31,229,31,68,31,213,31,58,31,224,31,136,31,136,30,159,31,13,31,133,31,45,31,193,31,69,31,172,31,54,31,11,31,11,30,206,31,206,30,103,31,103,30,103,29,77,31,77,30,68,31,68,30,252,31,207,31,241,31,112,31,92,31,72,31,199,31,140,31,222,31,55,31,236,31,136,31,167,31,208,31,208,30,223,31,151,31,24,31,4,31,157,31,157,30,180,31,180,30,180,29,195,31,53,31,184,31,149,31,149,30,109,31,85,31,27,31,142,31,214,31,214,30,118,31,118,30,118,29,168,31,168,30,58,31,39,31,5,31,232,31,231,31,115,31,86,31,112,31,106,31,249,31,249,30,249,29,62,31,78,31,104,31,238,31,238,30,133,31,186,31,108,31,124,31,124,30,125,31,198,31,252,31,32,31,32,30,32,29,88,31,88,30,153,31,234,31,27,31,27,31,181,31,153,31,118,31,240,31,179,31,5,31,5,30,200,31,137,31,137,30,23,31,82,31,145,31,39,31,212,31,135,31,135,30,8,31,134,31,12,31,153,31,102,31,134,31,202,31,245,31,245,30,245,29,213,31,213,30,141,31,190,31,137,31,137,30,204,31,253,31,253,30,159,31,179,31,135,31,163,31,163,30,94,31,124,31,126,31,98,31,181,31,53,31,152,31,57,31,141,31,83,31,189,31,118,31,193,31,55,31,55,30,55,29,55,28,106,31,12,31,72,31,127,31,68,31,7,31,173,31,29,31,29,30,14,31,171,31,208,31,211,31,137,31,137,30,203,31,51,31,240,31,234,31,186,31,186,30,159,31,142,31,142,30,12,31,78,31,133,31,133,30,175,31,39,31,32,31,124,31,124,30,129,31,189,31,176,31,176,30,176,29,7,31,58,31,58,30,236,31,35,31,191,31,231,31,58,31,98,31,98,30,33,31,33,30,184,31,184,30,28,31,28,30,37,31,114,31,119,31,154,31,105,31,105,30,203,31,41,31,55,31,234,31,234,30,103,31,135,31,166,31,138,31,138,30,50,31,50,30,93,31,118,31,169,31,212,31,29,31,29,30,75,31,75,30,75,29,191,31,92,31,200,31,216,31,232,31,98,31,101,31,30,31,63,31,170,31,208,31,144,31,144,30,7,31,107,31,107,30,213,31,68,31,237,31,222,31,96,31,85,31,207,31,79,31,120,31,46,31,72,31,164,31,164,30,51,31,77,31,77,30,107,31,93,31,72,31,196,31,183,31,106,31,148,31,234,31,173,31,53,31,201,31,212,31,146,31,146,30,52,31,69,31,188,31,68,31,68,30,255,31,103,31,86,31,148,31,109,31,71,31,167,31,97,31,176,31,24,31,24,30,203,31,144,31,144,30,110,31,23,31,160,31,160,30,50,31,171,31,158,31,208,31,248,31,155,31,171,31,171,30,79,31,155,31,30,31,103,31,103,30,201,31,156,31,84,31,83,31,208,31,202,31,31,31,222,31,222,30,214,31,214,30,44,31,216,31,216,30,58,31,75,31,55,31,127,31,219,31,161,31,48,31,202,31,123,31,162,31,187,31,143,31,143,30,168,31,158,31,62,31,89,31,188,31,121,31,121,30,121,29,131,31,131,30,30,31,127,31,127,30,52,31,95,31,76,31,76,30,76,29,200,31,200,30,51,31,51,30,199,31,164,31,120,31,14,31,52,31,4,31,163,31,207,31,116,31,145,31,145,30,12,31,210,31,210,30,95,31,163,31,184,31,184,30,146,31,156,31,140,31,146,31,96,31,121,31,188,31,18,31,170,31,170,30,5,31,5,30,5,29,211,31,30,31,136,31,55,31,55,30,51,31,204,31,132,31,255,31,48,31,97,31,97,30,197,31,18,31,57,31,117,31,23,31,53,31,111,31,111,30,159,31,198,31,23,31,181,31,55,31,55,30,116,31,31,31,246,31,178,31,178,30,124,31,13,31,124,31,155,31,22,31,18,31,18,30,188,31,178,31,11,31,9,31,118,31,223,31,132,31,29,31,11,31,236,31,75,31,4,31,4,30,187,31,28,31,12,31,12,30,12,29,12,28,73,31,174,31,118,31,215,31,14,31,3,31,86,31,159,31,34,31,169,31,73,31,61,31,235,31,200,31,200,30,248,31,248,31,101,31,101,30,239,31,223,31,50,31,102,31,216,31,88,31,162,31,111,31,118,31,90,31,63,31,177,31,177,30,2,31,85,31,102,31,82,31,82,30,216,31,50,31,50,31,142,31,48,31,156,31,206,31,165,31,114,31,246,31,57,31,215,31,201,31,1,31,75,31,213,31,106,31,191,31,144,31,102,31,110,31,30,31,65,31,113,31,113,30,113,29,157,31,145,31,239,31,191,31,99,31,160,31,160,30,160,29,160,28,211,31,129,31,97,31,207,31,212,31,228,31,86,31,18,31,132,31,195,31,195,30,194,31,121,31,76,31,9,31,79,31,10,31,194,31,93,31,11,31,95,31,82,31,31,31,244,31,7,31,250,31,250,30,130,31,130,31,207,31,207,30,253,31,89,31,25,31,25,30,58,31,46,31,75,31,149,31,153,31,52,31,26,31,17,31,202,31,181,31,181,30,54,31,54,30,239,31,73,31,192,31,118,31,118,30,118,29,118,28,162,31,156,31,156,30,77,31,77,30,56,31,55,31,192,31,114,31,114,30,23,31,23,30,92,31,176,31,176,30,187,31,20,31,186,31,186,30,132,31,232,31,247,31,247,30,30,31,30,30,162,31,48,31,195,31,87,31,252,31,126,31,236,31,136,31,136,30,136,29,136,28,136,27,167,31,219,31,159,31,197,31,131,31,255,31,255,30,10,31,209,31,198,31,179,31,247,31,118,31,195,31,117,31,61,31,23,31,154,31,117,31,117,30,128,31,49,31,52,31,52,30,52,29,52,28,73,31,220,31,34,31,34,30,34,29,93,31,214,31,242,31,184,31,61,31,192,31,137,31,137,30,45,31,43,31,186,31,146,31,48,31,158,31,139,31,157,31,130,31,225,31,181,31,237,31,180,31,180,30,15,31,227,31,133,31,154,31,105,31,236,31,127,31,245,31,144,31,218,31,248,31,223,31,223,30,79,31,232,31,131,31,166,31,163,31,251,31,133,31,242,31,114,31,238,31,148,31,177,31,33,31,220,31,50,31,60,31,156,31,42,31,147,31,209,31,150,31,55,31,55,30,254,31,78,31,118,31,118,30,211,31,211,30,13,31,174,31,88,31,218,31,218,30,218,29,234,31,53,31,234,31,234,30,221,31,66,31,89,31,2,31,185,31,185,30,189,31,198,31,104,31,57,31,92,31,226,31,235,31,235,30,223,31,166,31,241,31,241,30,175,31,252,31,252,30,220,31,221,31,155,31,215,31,136,31,47,31,179,31,39,31,178,31,119,31,119,30,227,31,96,31,51,31,247,31,114,31,166,31,238,31,226,31,57,31,143,31,143,30,49,31,187,31,86,31,86,30,86,29,132,31,59,31,59,30,59,29,111,31,206,31,204,31,118,31,232,31,89,31,89,30,216,31,216,30,130,31,217,31,217,30,103,31,156,31,187,31,148,31,242,31,120,31,180,31,249,31,249,30,105,31,109,31,200,31,83,31,231,31,68,31,115,31,229,31,228,31,34,31,55,31,55,30,156,31,131,31,109,31,32,31,19,31,19,30,18,31,224,31,22,31,22,30,86,31,86,30,138,31,223,31,74,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
