-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_217 is
end project_tb_217;

architecture project_tb_arch_217 of project_tb_217 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 860;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (44,0,0,0,0,0,39,0,179,0,242,0,47,0,220,0,174,0,16,0,253,0,124,0,239,0,82,0,244,0,0,0,50,0,242,0,65,0,78,0,30,0,147,0,100,0,0,0,0,0,8,0,12,0,126,0,0,0,0,0,188,0,0,0,28,0,214,0,220,0,12,0,140,0,117,0,113,0,109,0,129,0,139,0,212,0,0,0,77,0,226,0,0,0,76,0,100,0,10,0,238,0,1,0,0,0,163,0,143,0,250,0,219,0,233,0,23,0,8,0,132,0,200,0,219,0,229,0,149,0,178,0,60,0,0,0,66,0,0,0,181,0,25,0,253,0,121,0,12,0,60,0,77,0,0,0,53,0,135,0,160,0,170,0,75,0,186,0,76,0,88,0,0,0,139,0,251,0,46,0,77,0,200,0,86,0,0,0,246,0,230,0,191,0,15,0,23,0,3,0,48,0,110,0,0,0,0,0,246,0,0,0,0,0,57,0,207,0,22,0,20,0,59,0,179,0,119,0,254,0,227,0,56,0,102,0,42,0,168,0,84,0,159,0,114,0,184,0,0,0,133,0,229,0,6,0,203,0,0,0,0,0,0,0,212,0,223,0,156,0,0,0,206,0,133,0,125,0,25,0,0,0,124,0,13,0,101,0,72,0,166,0,58,0,43,0,156,0,171,0,209,0,171,0,0,0,14,0,190,0,0,0,233,0,0,0,0,0,189,0,110,0,167,0,0,0,0,0,84,0,147,0,174,0,40,0,68,0,118,0,203,0,105,0,243,0,219,0,0,0,81,0,234,0,52,0,187,0,121,0,208,0,0,0,121,0,202,0,115,0,173,0,193,0,32,0,178,0,70,0,110,0,127,0,203,0,201,0,59,0,225,0,0,0,181,0,0,0,223,0,44,0,242,0,251,0,34,0,0,0,131,0,56,0,126,0,170,0,129,0,240,0,74,0,0,0,72,0,106,0,0,0,0,0,221,0,125,0,124,0,0,0,120,0,44,0,211,0,128,0,50,0,0,0,251,0,0,0,148,0,79,0,25,0,0,0,0,0,213,0,129,0,208,0,144,0,0,0,205,0,69,0,4,0,37,0,0,0,0,0,53,0,0,0,40,0,230,0,218,0,0,0,212,0,194,0,112,0,158,0,246,0,243,0,96,0,0,0,115,0,0,0,0,0,0,0,207,0,37,0,2,0,0,0,13,0,255,0,0,0,66,0,60,0,134,0,182,0,79,0,55,0,0,0,0,0,46,0,98,0,179,0,211,0,74,0,0,0,227,0,232,0,180,0,69,0,25,0,0,0,180,0,247,0,112,0,17,0,0,0,39,0,122,0,0,0,123,0,0,0,58,0,0,0,41,0,0,0,0,0,255,0,164,0,252,0,220,0,133,0,245,0,25,0,199,0,103,0,223,0,206,0,67,0,30,0,0,0,96,0,237,0,150,0,150,0,22,0,141,0,128,0,151,0,5,0,102,0,21,0,0,0,167,0,0,0,127,0,63,0,170,0,253,0,224,0,252,0,51,0,0,0,128,0,0,0,183,0,165,0,192,0,164,0,183,0,0,0,74,0,150,0,182,0,211,0,211,0,167,0,0,0,0,0,161,0,178,0,160,0,3,0,6,0,0,0,122,0,49,0,0,0,224,0,0,0,0,0,237,0,140,0,141,0,240,0,7,0,183,0,208,0,160,0,183,0,64,0,56,0,111,0,20,0,171,0,198,0,97,0,225,0,130,0,107,0,199,0,57,0,0,0,0,0,93,0,0,0,103,0,22,0,189,0,81,0,227,0,142,0,142,0,214,0,7,0,96,0,10,0,0,0,154,0,0,0,120,0,0,0,218,0,67,0,164,0,238,0,239,0,121,0,1,0,0,0,141,0,153,0,222,0,250,0,2,0,214,0,12,0,159,0,198,0,22,0,179,0,194,0,94,0,96,0,87,0,126,0,166,0,0,0,66,0,222,0,215,0,105,0,59,0,63,0,235,0,0,0,63,0,56,0,202,0,77,0,176,0,21,0,0,0,0,0,209,0,0,0,206,0,78,0,147,0,0,0,122,0,180,0,106,0,215,0,80,0,218,0,0,0,101,0,191,0,199,0,0,0,166,0,229,0,17,0,0,0,0,0,0,0,129,0,0,0,0,0,63,0,20,0,39,0,242,0,130,0,180,0,195,0,222,0,152,0,81,0,194,0,0,0,44,0,139,0,116,0,188,0,101,0,0,0,70,0,0,0,0,0,252,0,125,0,141,0,0,0,0,0,219,0,26,0,43,0,0,0,183,0,0,0,0,0,218,0,192,0,203,0,229,0,114,0,243,0,0,0,213,0,0,0,230,0,0,0,214,0,111,0,235,0,0,0,0,0,137,0,219,0,94,0,55,0,85,0,0,0,19,0,204,0,0,0,0,0,0,0,13,0,236,0,169,0,96,0,253,0,181,0,0,0,23,0,0,0,0,0,134,0,22,0,222,0,76,0,203,0,143,0,230,0,86,0,26,0,244,0,183,0,0,0,186,0,95,0,0,0,143,0,175,0,105,0,85,0,72,0,46,0,250,0,25,0,0,0,13,0,245,0,249,0,76,0,19,0,80,0,96,0,224,0,62,0,243,0,207,0,157,0,49,0,188,0,142,0,0,0,0,0,53,0,243,0,29,0,60,0,123,0,130,0,183,0,0,0,10,0,64,0,53,0,219,0,186,0,81,0,225,0,33,0,29,0,127,0,0,0,27,0,53,0,48,0,0,0,0,0,119,0,0,0,140,0,122,0,135,0,16,0,0,0,132,0,136,0,78,0,5,0,209,0,204,0,254,0,79,0,0,0,204,0,249,0,38,0,112,0,51,0,172,0,21,0,0,0,212,0,23,0,0,0,0,0,56,0,172,0,228,0,100,0,0,0,14,0,74,0,0,0,136,0,11,0,107,0,191,0,209,0,21,0,62,0,32,0,14,0,0,0,0,0,40,0,153,0,215,0,0,0,211,0,11,0,0,0,71,0,195,0,129,0,128,0,134,0,181,0,0,0,220,0,0,0,35,0,39,0,61,0,39,0,0,0,58,0,179,0,249,0,62,0,0,0,79,0,167,0,134,0,0,0,0,0,193,0,11,0,134,0,0,0,140,0,186,0,0,0,0,0,124,0,178,0,8,0,82,0,68,0,53,0,14,0,249,0,0,0,187,0,0,0,0,0,190,0,0,0,157,0,37,0,0,0,159,0,56,0,0,0,9,0,164,0,0,0,7,0,144,0,188,0,68,0,246,0,16,0,124,0,51,0,224,0,0,0,220,0,72,0,144,0,226,0,69,0,172,0,217,0,164,0,122,0,141,0,9,0,49,0,0,0,0,0,5,0,73,0,6,0,0,0,143,0,127,0,138,0,0,0,0,0,127,0,53,0,19,0,66,0,0,0,6,0,0,0,135,0,106,0,123,0,48,0,3,0,212,0,79,0,176,0,198,0,0,0,173,0,90,0,59,0,4,0,180,0,194,0,28,0,0,0,151,0,175,0,0,0,83,0,103,0,160,0,113,0,59,0,28,0,253,0,83,0,0,0,74,0,155,0,56,0,153,0,31,0,8,0,24,0,140,0,230,0,91,0,113,0,122,0,41,0,60,0,105,0,82,0,0,0,0,0,181,0,103,0,105,0,122,0,0,0,9,0,123,0,0,0,135,0,59,0,0,0,132,0,140,0,10,0,208,0,0,0,233,0,207,0,27,0,136,0,0,0,77,0,10,0,226,0,239,0,146,0,153,0,0,0,4,0,27,0,226,0,232,0,0,0,0,0,0,0,192,0,50,0,162,0,78,0,0,0,161,0,70,0,0,0,0,0,194,0,73,0,117,0,173,0,171,0,16,0);
signal scenario_full  : scenario_type := (44,31,44,30,44,29,39,31,179,31,242,31,47,31,220,31,174,31,16,31,253,31,124,31,239,31,82,31,244,31,244,30,50,31,242,31,65,31,78,31,30,31,147,31,100,31,100,30,100,29,8,31,12,31,126,31,126,30,126,29,188,31,188,30,28,31,214,31,220,31,12,31,140,31,117,31,113,31,109,31,129,31,139,31,212,31,212,30,77,31,226,31,226,30,76,31,100,31,10,31,238,31,1,31,1,30,163,31,143,31,250,31,219,31,233,31,23,31,8,31,132,31,200,31,219,31,229,31,149,31,178,31,60,31,60,30,66,31,66,30,181,31,25,31,253,31,121,31,12,31,60,31,77,31,77,30,53,31,135,31,160,31,170,31,75,31,186,31,76,31,88,31,88,30,139,31,251,31,46,31,77,31,200,31,86,31,86,30,246,31,230,31,191,31,15,31,23,31,3,31,48,31,110,31,110,30,110,29,246,31,246,30,246,29,57,31,207,31,22,31,20,31,59,31,179,31,119,31,254,31,227,31,56,31,102,31,42,31,168,31,84,31,159,31,114,31,184,31,184,30,133,31,229,31,6,31,203,31,203,30,203,29,203,28,212,31,223,31,156,31,156,30,206,31,133,31,125,31,25,31,25,30,124,31,13,31,101,31,72,31,166,31,58,31,43,31,156,31,171,31,209,31,171,31,171,30,14,31,190,31,190,30,233,31,233,30,233,29,189,31,110,31,167,31,167,30,167,29,84,31,147,31,174,31,40,31,68,31,118,31,203,31,105,31,243,31,219,31,219,30,81,31,234,31,52,31,187,31,121,31,208,31,208,30,121,31,202,31,115,31,173,31,193,31,32,31,178,31,70,31,110,31,127,31,203,31,201,31,59,31,225,31,225,30,181,31,181,30,223,31,44,31,242,31,251,31,34,31,34,30,131,31,56,31,126,31,170,31,129,31,240,31,74,31,74,30,72,31,106,31,106,30,106,29,221,31,125,31,124,31,124,30,120,31,44,31,211,31,128,31,50,31,50,30,251,31,251,30,148,31,79,31,25,31,25,30,25,29,213,31,129,31,208,31,144,31,144,30,205,31,69,31,4,31,37,31,37,30,37,29,53,31,53,30,40,31,230,31,218,31,218,30,212,31,194,31,112,31,158,31,246,31,243,31,96,31,96,30,115,31,115,30,115,29,115,28,207,31,37,31,2,31,2,30,13,31,255,31,255,30,66,31,60,31,134,31,182,31,79,31,55,31,55,30,55,29,46,31,98,31,179,31,211,31,74,31,74,30,227,31,232,31,180,31,69,31,25,31,25,30,180,31,247,31,112,31,17,31,17,30,39,31,122,31,122,30,123,31,123,30,58,31,58,30,41,31,41,30,41,29,255,31,164,31,252,31,220,31,133,31,245,31,25,31,199,31,103,31,223,31,206,31,67,31,30,31,30,30,96,31,237,31,150,31,150,31,22,31,141,31,128,31,151,31,5,31,102,31,21,31,21,30,167,31,167,30,127,31,63,31,170,31,253,31,224,31,252,31,51,31,51,30,128,31,128,30,183,31,165,31,192,31,164,31,183,31,183,30,74,31,150,31,182,31,211,31,211,31,167,31,167,30,167,29,161,31,178,31,160,31,3,31,6,31,6,30,122,31,49,31,49,30,224,31,224,30,224,29,237,31,140,31,141,31,240,31,7,31,183,31,208,31,160,31,183,31,64,31,56,31,111,31,20,31,171,31,198,31,97,31,225,31,130,31,107,31,199,31,57,31,57,30,57,29,93,31,93,30,103,31,22,31,189,31,81,31,227,31,142,31,142,31,214,31,7,31,96,31,10,31,10,30,154,31,154,30,120,31,120,30,218,31,67,31,164,31,238,31,239,31,121,31,1,31,1,30,141,31,153,31,222,31,250,31,2,31,214,31,12,31,159,31,198,31,22,31,179,31,194,31,94,31,96,31,87,31,126,31,166,31,166,30,66,31,222,31,215,31,105,31,59,31,63,31,235,31,235,30,63,31,56,31,202,31,77,31,176,31,21,31,21,30,21,29,209,31,209,30,206,31,78,31,147,31,147,30,122,31,180,31,106,31,215,31,80,31,218,31,218,30,101,31,191,31,199,31,199,30,166,31,229,31,17,31,17,30,17,29,17,28,129,31,129,30,129,29,63,31,20,31,39,31,242,31,130,31,180,31,195,31,222,31,152,31,81,31,194,31,194,30,44,31,139,31,116,31,188,31,101,31,101,30,70,31,70,30,70,29,252,31,125,31,141,31,141,30,141,29,219,31,26,31,43,31,43,30,183,31,183,30,183,29,218,31,192,31,203,31,229,31,114,31,243,31,243,30,213,31,213,30,230,31,230,30,214,31,111,31,235,31,235,30,235,29,137,31,219,31,94,31,55,31,85,31,85,30,19,31,204,31,204,30,204,29,204,28,13,31,236,31,169,31,96,31,253,31,181,31,181,30,23,31,23,30,23,29,134,31,22,31,222,31,76,31,203,31,143,31,230,31,86,31,26,31,244,31,183,31,183,30,186,31,95,31,95,30,143,31,175,31,105,31,85,31,72,31,46,31,250,31,25,31,25,30,13,31,245,31,249,31,76,31,19,31,80,31,96,31,224,31,62,31,243,31,207,31,157,31,49,31,188,31,142,31,142,30,142,29,53,31,243,31,29,31,60,31,123,31,130,31,183,31,183,30,10,31,64,31,53,31,219,31,186,31,81,31,225,31,33,31,29,31,127,31,127,30,27,31,53,31,48,31,48,30,48,29,119,31,119,30,140,31,122,31,135,31,16,31,16,30,132,31,136,31,78,31,5,31,209,31,204,31,254,31,79,31,79,30,204,31,249,31,38,31,112,31,51,31,172,31,21,31,21,30,212,31,23,31,23,30,23,29,56,31,172,31,228,31,100,31,100,30,14,31,74,31,74,30,136,31,11,31,107,31,191,31,209,31,21,31,62,31,32,31,14,31,14,30,14,29,40,31,153,31,215,31,215,30,211,31,11,31,11,30,71,31,195,31,129,31,128,31,134,31,181,31,181,30,220,31,220,30,35,31,39,31,61,31,39,31,39,30,58,31,179,31,249,31,62,31,62,30,79,31,167,31,134,31,134,30,134,29,193,31,11,31,134,31,134,30,140,31,186,31,186,30,186,29,124,31,178,31,8,31,82,31,68,31,53,31,14,31,249,31,249,30,187,31,187,30,187,29,190,31,190,30,157,31,37,31,37,30,159,31,56,31,56,30,9,31,164,31,164,30,7,31,144,31,188,31,68,31,246,31,16,31,124,31,51,31,224,31,224,30,220,31,72,31,144,31,226,31,69,31,172,31,217,31,164,31,122,31,141,31,9,31,49,31,49,30,49,29,5,31,73,31,6,31,6,30,143,31,127,31,138,31,138,30,138,29,127,31,53,31,19,31,66,31,66,30,6,31,6,30,135,31,106,31,123,31,48,31,3,31,212,31,79,31,176,31,198,31,198,30,173,31,90,31,59,31,4,31,180,31,194,31,28,31,28,30,151,31,175,31,175,30,83,31,103,31,160,31,113,31,59,31,28,31,253,31,83,31,83,30,74,31,155,31,56,31,153,31,31,31,8,31,24,31,140,31,230,31,91,31,113,31,122,31,41,31,60,31,105,31,82,31,82,30,82,29,181,31,103,31,105,31,122,31,122,30,9,31,123,31,123,30,135,31,59,31,59,30,132,31,140,31,10,31,208,31,208,30,233,31,207,31,27,31,136,31,136,30,77,31,10,31,226,31,239,31,146,31,153,31,153,30,4,31,27,31,226,31,232,31,232,30,232,29,232,28,192,31,50,31,162,31,78,31,78,30,161,31,70,31,70,30,70,29,194,31,73,31,117,31,173,31,171,31,16,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
