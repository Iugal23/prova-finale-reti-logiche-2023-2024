-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 286;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (191,0,233,0,0,0,156,0,135,0,56,0,103,0,231,0,85,0,25,0,0,0,137,0,124,0,170,0,163,0,11,0,209,0,0,0,175,0,37,0,109,0,90,0,185,0,207,0,86,0,116,0,252,0,164,0,238,0,6,0,14,0,202,0,62,0,178,0,24,0,174,0,86,0,51,0,100,0,0,0,242,0,43,0,0,0,0,0,165,0,80,0,69,0,190,0,67,0,172,0,22,0,27,0,73,0,0,0,194,0,0,0,218,0,251,0,14,0,101,0,153,0,245,0,33,0,169,0,204,0,103,0,239,0,0,0,116,0,0,0,59,0,66,0,91,0,189,0,0,0,194,0,105,0,171,0,92,0,139,0,144,0,207,0,211,0,0,0,230,0,109,0,94,0,174,0,134,0,12,0,220,0,218,0,0,0,202,0,162,0,15,0,0,0,254,0,0,0,0,0,185,0,150,0,77,0,137,0,199,0,109,0,59,0,0,0,170,0,60,0,126,0,0,0,157,0,4,0,28,0,49,0,0,0,133,0,250,0,63,0,3,0,0,0,253,0,64,0,132,0,79,0,0,0,0,0,247,0,230,0,0,0,109,0,105,0,99,0,6,0,166,0,196,0,55,0,212,0,0,0,210,0,0,0,0,0,0,0,88,0,0,0,142,0,223,0,0,0,136,0,231,0,253,0,0,0,51,0,101,0,133,0,0,0,52,0,0,0,16,0,222,0,117,0,0,0,56,0,84,0,54,0,145,0,0,0,248,0,101,0,4,0,146,0,0,0,0,0,236,0,252,0,145,0,0,0,252,0,189,0,160,0,230,0,48,0,148,0,219,0,155,0,107,0,113,0,173,0,28,0,214,0,152,0,246,0,141,0,186,0,63,0,29,0,0,0,141,0,0,0,181,0,70,0,254,0,0,0,201,0,113,0,173,0,0,0,0,0,0,0,0,0,167,0,67,0,29,0,191,0,49,0,22,0,50,0,0,0,143,0,8,0,86,0,190,0,202,0,162,0,56,0,0,0,163,0,90,0,69,0,175,0,56,0,62,0,112,0,52,0,0,0,206,0,0,0,4,0,4,0,147,0,124,0,35,0,130,0,118,0,42,0,82,0,96,0,0,0,206,0,0,0,13,0,0,0,0,0,0,0,104,0,0,0,58,0,98,0,148,0,0,0,0,0,219,0,0,0,12,0,0,0,33,0,0,0,135,0,248,0,1,0,242,0,45,0,0,0,164,0,200,0,183,0,135,0,201,0,223,0,239,0,157,0,0,0,254,0,192,0,72,0);
signal scenario_full  : scenario_type := (191,31,233,31,233,30,156,31,135,31,56,31,103,31,231,31,85,31,25,31,25,30,137,31,124,31,170,31,163,31,11,31,209,31,209,30,175,31,37,31,109,31,90,31,185,31,207,31,86,31,116,31,252,31,164,31,238,31,6,31,14,31,202,31,62,31,178,31,24,31,174,31,86,31,51,31,100,31,100,30,242,31,43,31,43,30,43,29,165,31,80,31,69,31,190,31,67,31,172,31,22,31,27,31,73,31,73,30,194,31,194,30,218,31,251,31,14,31,101,31,153,31,245,31,33,31,169,31,204,31,103,31,239,31,239,30,116,31,116,30,59,31,66,31,91,31,189,31,189,30,194,31,105,31,171,31,92,31,139,31,144,31,207,31,211,31,211,30,230,31,109,31,94,31,174,31,134,31,12,31,220,31,218,31,218,30,202,31,162,31,15,31,15,30,254,31,254,30,254,29,185,31,150,31,77,31,137,31,199,31,109,31,59,31,59,30,170,31,60,31,126,31,126,30,157,31,4,31,28,31,49,31,49,30,133,31,250,31,63,31,3,31,3,30,253,31,64,31,132,31,79,31,79,30,79,29,247,31,230,31,230,30,109,31,105,31,99,31,6,31,166,31,196,31,55,31,212,31,212,30,210,31,210,30,210,29,210,28,88,31,88,30,142,31,223,31,223,30,136,31,231,31,253,31,253,30,51,31,101,31,133,31,133,30,52,31,52,30,16,31,222,31,117,31,117,30,56,31,84,31,54,31,145,31,145,30,248,31,101,31,4,31,146,31,146,30,146,29,236,31,252,31,145,31,145,30,252,31,189,31,160,31,230,31,48,31,148,31,219,31,155,31,107,31,113,31,173,31,28,31,214,31,152,31,246,31,141,31,186,31,63,31,29,31,29,30,141,31,141,30,181,31,70,31,254,31,254,30,201,31,113,31,173,31,173,30,173,29,173,28,173,27,167,31,67,31,29,31,191,31,49,31,22,31,50,31,50,30,143,31,8,31,86,31,190,31,202,31,162,31,56,31,56,30,163,31,90,31,69,31,175,31,56,31,62,31,112,31,52,31,52,30,206,31,206,30,4,31,4,31,147,31,124,31,35,31,130,31,118,31,42,31,82,31,96,31,96,30,206,31,206,30,13,31,13,30,13,29,13,28,104,31,104,30,58,31,98,31,148,31,148,30,148,29,219,31,219,30,12,31,12,30,33,31,33,30,135,31,248,31,1,31,242,31,45,31,45,30,164,31,200,31,183,31,135,31,201,31,223,31,239,31,157,31,157,30,254,31,192,31,72,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
