-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_737 is
end project_tb_737;

architecture project_tb_arch_737 of project_tb_737 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 783;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (102,0,0,0,8,0,209,0,0,0,110,0,155,0,67,0,68,0,0,0,104,0,112,0,2,0,0,0,12,0,0,0,206,0,242,0,240,0,0,0,25,0,182,0,185,0,92,0,133,0,36,0,131,0,58,0,0,0,80,0,233,0,198,0,103,0,220,0,0,0,238,0,101,0,211,0,115,0,15,0,124,0,4,0,9,0,132,0,0,0,160,0,118,0,139,0,187,0,0,0,0,0,16,0,122,0,0,0,0,0,92,0,133,0,227,0,0,0,0,0,121,0,0,0,251,0,180,0,0,0,106,0,51,0,142,0,154,0,78,0,142,0,0,0,0,0,0,0,155,0,14,0,87,0,222,0,0,0,182,0,74,0,82,0,186,0,0,0,0,0,66,0,167,0,0,0,22,0,0,0,58,0,32,0,36,0,136,0,219,0,254,0,200,0,91,0,0,0,111,0,62,0,185,0,208,0,242,0,117,0,141,0,0,0,119,0,209,0,3,0,0,0,206,0,0,0,122,0,129,0,46,0,199,0,5,0,219,0,0,0,0,0,206,0,141,0,253,0,112,0,13,0,126,0,186,0,113,0,49,0,228,0,174,0,235,0,128,0,199,0,0,0,71,0,178,0,202,0,77,0,31,0,23,0,225,0,194,0,0,0,25,0,0,0,240,0,202,0,0,0,0,0,0,0,0,0,1,0,0,0,0,0,0,0,0,0,82,0,0,0,208,0,0,0,0,0,54,0,235,0,130,0,81,0,34,0,175,0,1,0,12,0,107,0,234,0,0,0,161,0,81,0,246,0,91,0,0,0,10,0,250,0,7,0,0,0,146,0,0,0,44,0,0,0,61,0,239,0,236,0,254,0,0,0,13,0,50,0,10,0,223,0,137,0,207,0,248,0,76,0,242,0,251,0,9,0,0,0,156,0,155,0,0,0,94,0,0,0,8,0,16,0,44,0,203,0,0,0,181,0,112,0,253,0,0,0,0,0,0,0,51,0,108,0,0,0,15,0,215,0,235,0,0,0,110,0,0,0,113,0,100,0,181,0,0,0,227,0,193,0,106,0,127,0,221,0,31,0,103,0,61,0,32,0,0,0,193,0,0,0,176,0,124,0,188,0,206,0,215,0,190,0,243,0,0,0,0,0,141,0,63,0,0,0,15,0,113,0,168,0,0,0,0,0,61,0,60,0,0,0,216,0,68,0,146,0,193,0,245,0,30,0,235,0,241,0,133,0,251,0,224,0,245,0,121,0,235,0,0,0,247,0,172,0,247,0,254,0,1,0,209,0,162,0,87,0,0,0,59,0,136,0,49,0,186,0,125,0,73,0,36,0,0,0,3,0,84,0,0,0,0,0,244,0,184,0,106,0,131,0,192,0,3,0,31,0,124,0,110,0,0,0,83,0,0,0,192,0,97,0,3,0,113,0,0,0,189,0,219,0,113,0,0,0,176,0,151,0,177,0,245,0,0,0,142,0,146,0,102,0,222,0,64,0,198,0,164,0,48,0,82,0,0,0,2,0,0,0,155,0,121,0,0,0,55,0,92,0,44,0,220,0,193,0,152,0,42,0,75,0,99,0,103,0,108,0,160,0,183,0,0,0,0,0,89,0,14,0,201,0,195,0,0,0,53,0,232,0,0,0,0,0,199,0,0,0,0,0,247,0,61,0,68,0,210,0,0,0,216,0,0,0,195,0,180,0,200,0,97,0,22,0,108,0,237,0,0,0,186,0,239,0,96,0,1,0,249,0,170,0,0,0,135,0,142,0,64,0,2,0,41,0,22,0,139,0,156,0,9,0,35,0,151,0,209,0,0,0,138,0,131,0,199,0,254,0,0,0,21,0,186,0,47,0,149,0,0,0,0,0,0,0,95,0,0,0,203,0,68,0,0,0,130,0,0,0,0,0,238,0,114,0,0,0,104,0,163,0,5,0,0,0,98,0,128,0,71,0,76,0,108,0,181,0,183,0,214,0,0,0,32,0,255,0,145,0,247,0,0,0,247,0,79,0,0,0,109,0,41,0,0,0,217,0,58,0,44,0,83,0,175,0,0,0,148,0,201,0,153,0,193,0,102,0,154,0,64,0,222,0,65,0,122,0,0,0,153,0,144,0,0,0,0,0,0,0,0,0,0,0,32,0,51,0,201,0,169,0,242,0,98,0,0,0,180,0,215,0,200,0,117,0,58,0,94,0,0,0,25,0,208,0,189,0,39,0,7,0,209,0,234,0,251,0,206,0,33,0,0,0,14,0,204,0,138,0,148,0,77,0,26,0,79,0,236,0,45,0,208,0,128,0,0,0,142,0,112,0,78,0,62,0,65,0,209,0,177,0,0,0,0,0,17,0,242,0,50,0,128,0,0,0,117,0,13,0,18,0,0,0,0,0,243,0,176,0,0,0,196,0,250,0,104,0,253,0,88,0,54,0,0,0,216,0,100,0,186,0,0,0,60,0,0,0,0,0,204,0,52,0,2,0,87,0,163,0,194,0,0,0,0,0,114,0,65,0,139,0,71,0,22,0,235,0,210,0,180,0,195,0,125,0,0,0,93,0,217,0,184,0,0,0,239,0,185,0,193,0,221,0,37,0,112,0,127,0,30,0,245,0,37,0,0,0,0,0,0,0,0,0,26,0,235,0,0,0,0,0,140,0,136,0,208,0,0,0,185,0,0,0,79,0,0,0,75,0,8,0,0,0,119,0,176,0,108,0,0,0,4,0,0,0,200,0,167,0,35,0,0,0,16,0,95,0,0,0,166,0,0,0,0,0,182,0,144,0,183,0,0,0,141,0,29,0,158,0,118,0,164,0,1,0,59,0,26,0,227,0,236,0,242,0,32,0,0,0,183,0,95,0,63,0,253,0,25,0,131,0,86,0,54,0,58,0,83,0,61,0,217,0,249,0,14,0,84,0,24,0,183,0,143,0,207,0,10,0,202,0,155,0,58,0,253,0,0,0,0,0,0,0,142,0,240,0,118,0,108,0,234,0,133,0,17,0,0,0,162,0,0,0,109,0,198,0,107,0,249,0,216,0,240,0,0,0,182,0,253,0,9,0,0,0,56,0,83,0,141,0,87,0,48,0,207,0,189,0,28,0,141,0,224,0,240,0,176,0,214,0,0,0,0,0,0,0,61,0,234,0,109,0,131,0,36,0,110,0,141,0,30,0,203,0,180,0,165,0,12,0,20,0,4,0,154,0,0,0,28,0,12,0,104,0,201,0,0,0,254,0,49,0,209,0,238,0,239,0,85,0,21,0,0,0,0,0,127,0,172,0,78,0,29,0,61,0,81,0,35,0,140,0,118,0,0,0,33,0,58,0,239,0,254,0,219,0,0,0,7,0,82,0,168,0,22,0,60,0,128,0,0,0,0,0,214,0,171,0,243,0,0,0,220,0,0,0,46,0,164,0,147,0,124,0,0,0,0,0,80,0,0,0,0,0,88,0,202,0,106,0,133,0,240,0,204,0,234,0,233,0,202,0,32,0,172,0,175,0,220,0,22,0,0,0,30,0,251,0);
signal scenario_full  : scenario_type := (102,31,102,30,8,31,209,31,209,30,110,31,155,31,67,31,68,31,68,30,104,31,112,31,2,31,2,30,12,31,12,30,206,31,242,31,240,31,240,30,25,31,182,31,185,31,92,31,133,31,36,31,131,31,58,31,58,30,80,31,233,31,198,31,103,31,220,31,220,30,238,31,101,31,211,31,115,31,15,31,124,31,4,31,9,31,132,31,132,30,160,31,118,31,139,31,187,31,187,30,187,29,16,31,122,31,122,30,122,29,92,31,133,31,227,31,227,30,227,29,121,31,121,30,251,31,180,31,180,30,106,31,51,31,142,31,154,31,78,31,142,31,142,30,142,29,142,28,155,31,14,31,87,31,222,31,222,30,182,31,74,31,82,31,186,31,186,30,186,29,66,31,167,31,167,30,22,31,22,30,58,31,32,31,36,31,136,31,219,31,254,31,200,31,91,31,91,30,111,31,62,31,185,31,208,31,242,31,117,31,141,31,141,30,119,31,209,31,3,31,3,30,206,31,206,30,122,31,129,31,46,31,199,31,5,31,219,31,219,30,219,29,206,31,141,31,253,31,112,31,13,31,126,31,186,31,113,31,49,31,228,31,174,31,235,31,128,31,199,31,199,30,71,31,178,31,202,31,77,31,31,31,23,31,225,31,194,31,194,30,25,31,25,30,240,31,202,31,202,30,202,29,202,28,202,27,1,31,1,30,1,29,1,28,1,27,82,31,82,30,208,31,208,30,208,29,54,31,235,31,130,31,81,31,34,31,175,31,1,31,12,31,107,31,234,31,234,30,161,31,81,31,246,31,91,31,91,30,10,31,250,31,7,31,7,30,146,31,146,30,44,31,44,30,61,31,239,31,236,31,254,31,254,30,13,31,50,31,10,31,223,31,137,31,207,31,248,31,76,31,242,31,251,31,9,31,9,30,156,31,155,31,155,30,94,31,94,30,8,31,16,31,44,31,203,31,203,30,181,31,112,31,253,31,253,30,253,29,253,28,51,31,108,31,108,30,15,31,215,31,235,31,235,30,110,31,110,30,113,31,100,31,181,31,181,30,227,31,193,31,106,31,127,31,221,31,31,31,103,31,61,31,32,31,32,30,193,31,193,30,176,31,124,31,188,31,206,31,215,31,190,31,243,31,243,30,243,29,141,31,63,31,63,30,15,31,113,31,168,31,168,30,168,29,61,31,60,31,60,30,216,31,68,31,146,31,193,31,245,31,30,31,235,31,241,31,133,31,251,31,224,31,245,31,121,31,235,31,235,30,247,31,172,31,247,31,254,31,1,31,209,31,162,31,87,31,87,30,59,31,136,31,49,31,186,31,125,31,73,31,36,31,36,30,3,31,84,31,84,30,84,29,244,31,184,31,106,31,131,31,192,31,3,31,31,31,124,31,110,31,110,30,83,31,83,30,192,31,97,31,3,31,113,31,113,30,189,31,219,31,113,31,113,30,176,31,151,31,177,31,245,31,245,30,142,31,146,31,102,31,222,31,64,31,198,31,164,31,48,31,82,31,82,30,2,31,2,30,155,31,121,31,121,30,55,31,92,31,44,31,220,31,193,31,152,31,42,31,75,31,99,31,103,31,108,31,160,31,183,31,183,30,183,29,89,31,14,31,201,31,195,31,195,30,53,31,232,31,232,30,232,29,199,31,199,30,199,29,247,31,61,31,68,31,210,31,210,30,216,31,216,30,195,31,180,31,200,31,97,31,22,31,108,31,237,31,237,30,186,31,239,31,96,31,1,31,249,31,170,31,170,30,135,31,142,31,64,31,2,31,41,31,22,31,139,31,156,31,9,31,35,31,151,31,209,31,209,30,138,31,131,31,199,31,254,31,254,30,21,31,186,31,47,31,149,31,149,30,149,29,149,28,95,31,95,30,203,31,68,31,68,30,130,31,130,30,130,29,238,31,114,31,114,30,104,31,163,31,5,31,5,30,98,31,128,31,71,31,76,31,108,31,181,31,183,31,214,31,214,30,32,31,255,31,145,31,247,31,247,30,247,31,79,31,79,30,109,31,41,31,41,30,217,31,58,31,44,31,83,31,175,31,175,30,148,31,201,31,153,31,193,31,102,31,154,31,64,31,222,31,65,31,122,31,122,30,153,31,144,31,144,30,144,29,144,28,144,27,144,26,32,31,51,31,201,31,169,31,242,31,98,31,98,30,180,31,215,31,200,31,117,31,58,31,94,31,94,30,25,31,208,31,189,31,39,31,7,31,209,31,234,31,251,31,206,31,33,31,33,30,14,31,204,31,138,31,148,31,77,31,26,31,79,31,236,31,45,31,208,31,128,31,128,30,142,31,112,31,78,31,62,31,65,31,209,31,177,31,177,30,177,29,17,31,242,31,50,31,128,31,128,30,117,31,13,31,18,31,18,30,18,29,243,31,176,31,176,30,196,31,250,31,104,31,253,31,88,31,54,31,54,30,216,31,100,31,186,31,186,30,60,31,60,30,60,29,204,31,52,31,2,31,87,31,163,31,194,31,194,30,194,29,114,31,65,31,139,31,71,31,22,31,235,31,210,31,180,31,195,31,125,31,125,30,93,31,217,31,184,31,184,30,239,31,185,31,193,31,221,31,37,31,112,31,127,31,30,31,245,31,37,31,37,30,37,29,37,28,37,27,26,31,235,31,235,30,235,29,140,31,136,31,208,31,208,30,185,31,185,30,79,31,79,30,75,31,8,31,8,30,119,31,176,31,108,31,108,30,4,31,4,30,200,31,167,31,35,31,35,30,16,31,95,31,95,30,166,31,166,30,166,29,182,31,144,31,183,31,183,30,141,31,29,31,158,31,118,31,164,31,1,31,59,31,26,31,227,31,236,31,242,31,32,31,32,30,183,31,95,31,63,31,253,31,25,31,131,31,86,31,54,31,58,31,83,31,61,31,217,31,249,31,14,31,84,31,24,31,183,31,143,31,207,31,10,31,202,31,155,31,58,31,253,31,253,30,253,29,253,28,142,31,240,31,118,31,108,31,234,31,133,31,17,31,17,30,162,31,162,30,109,31,198,31,107,31,249,31,216,31,240,31,240,30,182,31,253,31,9,31,9,30,56,31,83,31,141,31,87,31,48,31,207,31,189,31,28,31,141,31,224,31,240,31,176,31,214,31,214,30,214,29,214,28,61,31,234,31,109,31,131,31,36,31,110,31,141,31,30,31,203,31,180,31,165,31,12,31,20,31,4,31,154,31,154,30,28,31,12,31,104,31,201,31,201,30,254,31,49,31,209,31,238,31,239,31,85,31,21,31,21,30,21,29,127,31,172,31,78,31,29,31,61,31,81,31,35,31,140,31,118,31,118,30,33,31,58,31,239,31,254,31,219,31,219,30,7,31,82,31,168,31,22,31,60,31,128,31,128,30,128,29,214,31,171,31,243,31,243,30,220,31,220,30,46,31,164,31,147,31,124,31,124,30,124,29,80,31,80,30,80,29,88,31,202,31,106,31,133,31,240,31,204,31,234,31,233,31,202,31,32,31,172,31,175,31,220,31,22,31,22,30,30,31,251,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
