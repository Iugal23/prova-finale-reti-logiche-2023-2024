-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_880 is
end project_tb_880;

architecture project_tb_arch_880 of project_tb_880 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 668;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (65,0,0,0,192,0,86,0,63,0,31,0,15,0,66,0,217,0,36,0,229,0,0,0,101,0,14,0,165,0,214,0,0,0,0,0,189,0,61,0,219,0,0,0,54,0,0,0,61,0,24,0,217,0,127,0,51,0,232,0,0,0,134,0,182,0,172,0,139,0,37,0,0,0,139,0,8,0,245,0,180,0,138,0,111,0,0,0,17,0,115,0,93,0,82,0,91,0,0,0,253,0,238,0,6,0,162,0,116,0,232,0,232,0,219,0,0,0,112,0,244,0,233,0,210,0,127,0,0,0,208,0,243,0,172,0,147,0,0,0,142,0,0,0,68,0,32,0,45,0,85,0,41,0,206,0,179,0,35,0,100,0,184,0,0,0,130,0,102,0,238,0,194,0,124,0,231,0,0,0,0,0,214,0,211,0,204,0,239,0,0,0,76,0,0,0,0,0,47,0,130,0,48,0,0,0,125,0,12,0,100,0,13,0,247,0,254,0,201,0,0,0,159,0,208,0,0,0,68,0,138,0,180,0,25,0,119,0,218,0,238,0,36,0,75,0,0,0,0,0,208,0,0,0,90,0,0,0,239,0,230,0,52,0,149,0,38,0,241,0,182,0,152,0,0,0,184,0,136,0,212,0,0,0,112,0,193,0,181,0,196,0,0,0,0,0,139,0,53,0,150,0,14,0,3,0,27,0,91,0,234,0,118,0,156,0,10,0,144,0,120,0,0,0,80,0,187,0,102,0,234,0,64,0,14,0,24,0,199,0,159,0,43,0,180,0,0,0,169,0,8,0,99,0,67,0,0,0,0,0,126,0,89,0,90,0,24,0,6,0,231,0,0,0,111,0,172,0,149,0,0,0,58,0,49,0,167,0,24,0,37,0,0,0,112,0,83,0,92,0,179,0,0,0,176,0,36,0,0,0,0,0,172,0,254,0,14,0,175,0,221,0,162,0,62,0,0,0,133,0,188,0,0,0,0,0,0,0,93,0,49,0,121,0,0,0,140,0,67,0,146,0,0,0,245,0,0,0,53,0,0,0,3,0,31,0,78,0,236,0,40,0,108,0,0,0,0,0,0,0,67,0,159,0,180,0,101,0,85,0,33,0,0,0,62,0,115,0,115,0,255,0,182,0,0,0,150,0,180,0,9,0,11,0,15,0,0,0,154,0,216,0,57,0,159,0,161,0,0,0,230,0,0,0,80,0,0,0,12,0,0,0,85,0,60,0,0,0,60,0,22,0,53,0,245,0,0,0,207,0,247,0,235,0,0,0,0,0,244,0,147,0,25,0,0,0,173,0,59,0,130,0,0,0,0,0,0,0,93,0,0,0,0,0,188,0,45,0,242,0,135,0,161,0,71,0,0,0,161,0,98,0,135,0,104,0,245,0,17,0,49,0,114,0,86,0,96,0,157,0,38,0,142,0,207,0,96,0,244,0,81,0,254,0,0,0,159,0,69,0,0,0,5,0,0,0,145,0,255,0,24,0,100,0,137,0,45,0,0,0,0,0,236,0,248,0,0,0,0,0,89,0,121,0,0,0,111,0,0,0,0,0,79,0,63,0,69,0,165,0,184,0,21,0,91,0,249,0,0,0,53,0,94,0,0,0,0,0,75,0,0,0,178,0,1,0,0,0,90,0,76,0,207,0,118,0,97,0,112,0,0,0,81,0,61,0,47,0,170,0,116,0,49,0,189,0,80,0,40,0,102,0,138,0,57,0,106,0,43,0,120,0,218,0,134,0,0,0,5,0,70,0,192,0,39,0,0,0,180,0,0,0,54,0,188,0,122,0,50,0,0,0,55,0,42,0,53,0,48,0,74,0,179,0,226,0,56,0,0,0,238,0,0,0,220,0,238,0,231,0,234,0,114,0,111,0,71,0,0,0,52,0,0,0,153,0,244,0,0,0,0,0,178,0,98,0,0,0,199,0,236,0,0,0,128,0,0,0,98,0,48,0,40,0,198,0,0,0,0,0,212,0,0,0,167,0,78,0,117,0,106,0,0,0,242,0,247,0,0,0,71,0,48,0,94,0,169,0,126,0,12,0,28,0,138,0,248,0,43,0,228,0,235,0,113,0,164,0,163,0,167,0,227,0,0,0,119,0,169,0,40,0,89,0,0,0,75,0,67,0,17,0,38,0,0,0,101,0,45,0,0,0,228,0,0,0,0,0,163,0,0,0,8,0,5,0,129,0,170,0,0,0,55,0,44,0,56,0,230,0,31,0,241,0,0,0,239,0,86,0,168,0,179,0,209,0,103,0,64,0,0,0,252,0,135,0,219,0,104,0,197,0,0,0,10,0,0,0,179,0,36,0,30,0,162,0,0,0,208,0,29,0,179,0,16,0,136,0,83,0,118,0,101,0,31,0,71,0,59,0,63,0,0,0,79,0,0,0,83,0,52,0,3,0,0,0,181,0,65,0,19,0,0,0,0,0,0,0,0,0,14,0,144,0,88,0,0,0,74,0,30,0,151,0,0,0,108,0,49,0,0,0,221,0,0,0,227,0,64,0,183,0,195,0,0,0,249,0,0,0,219,0,242,0,0,0,119,0,0,0,50,0,113,0,55,0,116,0,0,0,7,0,112,0,0,0,0,0,0,0,202,0,154,0,57,0,184,0,0,0,72,0,129,0,160,0,0,0,79,0,241,0,41,0,238,0,73,0,0,0,230,0,118,0,170,0,92,0,0,0,0,0,234,0,182,0,47,0,151,0,219,0,130,0,0,0,206,0,76,0,82,0,29,0,134,0,4,0,91,0,15,0,46,0,111,0,194,0,64,0,132,0,36,0,82,0,168,0,126,0,0,0,205,0,159,0,108,0,95,0,0,0,188,0,0,0,37,0,0,0,124,0,254,0,96,0,49,0,19,0,132,0,142,0,163,0,0,0,112,0,217,0,119,0,237,0,171,0,39,0,220,0,0,0,12,0,198,0,254,0,0,0,214,0,15,0,77,0,153,0,233,0,236,0,41,0,118,0,74,0,0,0,241,0,19,0);
signal scenario_full  : scenario_type := (65,31,65,30,192,31,86,31,63,31,31,31,15,31,66,31,217,31,36,31,229,31,229,30,101,31,14,31,165,31,214,31,214,30,214,29,189,31,61,31,219,31,219,30,54,31,54,30,61,31,24,31,217,31,127,31,51,31,232,31,232,30,134,31,182,31,172,31,139,31,37,31,37,30,139,31,8,31,245,31,180,31,138,31,111,31,111,30,17,31,115,31,93,31,82,31,91,31,91,30,253,31,238,31,6,31,162,31,116,31,232,31,232,31,219,31,219,30,112,31,244,31,233,31,210,31,127,31,127,30,208,31,243,31,172,31,147,31,147,30,142,31,142,30,68,31,32,31,45,31,85,31,41,31,206,31,179,31,35,31,100,31,184,31,184,30,130,31,102,31,238,31,194,31,124,31,231,31,231,30,231,29,214,31,211,31,204,31,239,31,239,30,76,31,76,30,76,29,47,31,130,31,48,31,48,30,125,31,12,31,100,31,13,31,247,31,254,31,201,31,201,30,159,31,208,31,208,30,68,31,138,31,180,31,25,31,119,31,218,31,238,31,36,31,75,31,75,30,75,29,208,31,208,30,90,31,90,30,239,31,230,31,52,31,149,31,38,31,241,31,182,31,152,31,152,30,184,31,136,31,212,31,212,30,112,31,193,31,181,31,196,31,196,30,196,29,139,31,53,31,150,31,14,31,3,31,27,31,91,31,234,31,118,31,156,31,10,31,144,31,120,31,120,30,80,31,187,31,102,31,234,31,64,31,14,31,24,31,199,31,159,31,43,31,180,31,180,30,169,31,8,31,99,31,67,31,67,30,67,29,126,31,89,31,90,31,24,31,6,31,231,31,231,30,111,31,172,31,149,31,149,30,58,31,49,31,167,31,24,31,37,31,37,30,112,31,83,31,92,31,179,31,179,30,176,31,36,31,36,30,36,29,172,31,254,31,14,31,175,31,221,31,162,31,62,31,62,30,133,31,188,31,188,30,188,29,188,28,93,31,49,31,121,31,121,30,140,31,67,31,146,31,146,30,245,31,245,30,53,31,53,30,3,31,31,31,78,31,236,31,40,31,108,31,108,30,108,29,108,28,67,31,159,31,180,31,101,31,85,31,33,31,33,30,62,31,115,31,115,31,255,31,182,31,182,30,150,31,180,31,9,31,11,31,15,31,15,30,154,31,216,31,57,31,159,31,161,31,161,30,230,31,230,30,80,31,80,30,12,31,12,30,85,31,60,31,60,30,60,31,22,31,53,31,245,31,245,30,207,31,247,31,235,31,235,30,235,29,244,31,147,31,25,31,25,30,173,31,59,31,130,31,130,30,130,29,130,28,93,31,93,30,93,29,188,31,45,31,242,31,135,31,161,31,71,31,71,30,161,31,98,31,135,31,104,31,245,31,17,31,49,31,114,31,86,31,96,31,157,31,38,31,142,31,207,31,96,31,244,31,81,31,254,31,254,30,159,31,69,31,69,30,5,31,5,30,145,31,255,31,24,31,100,31,137,31,45,31,45,30,45,29,236,31,248,31,248,30,248,29,89,31,121,31,121,30,111,31,111,30,111,29,79,31,63,31,69,31,165,31,184,31,21,31,91,31,249,31,249,30,53,31,94,31,94,30,94,29,75,31,75,30,178,31,1,31,1,30,90,31,76,31,207,31,118,31,97,31,112,31,112,30,81,31,61,31,47,31,170,31,116,31,49,31,189,31,80,31,40,31,102,31,138,31,57,31,106,31,43,31,120,31,218,31,134,31,134,30,5,31,70,31,192,31,39,31,39,30,180,31,180,30,54,31,188,31,122,31,50,31,50,30,55,31,42,31,53,31,48,31,74,31,179,31,226,31,56,31,56,30,238,31,238,30,220,31,238,31,231,31,234,31,114,31,111,31,71,31,71,30,52,31,52,30,153,31,244,31,244,30,244,29,178,31,98,31,98,30,199,31,236,31,236,30,128,31,128,30,98,31,48,31,40,31,198,31,198,30,198,29,212,31,212,30,167,31,78,31,117,31,106,31,106,30,242,31,247,31,247,30,71,31,48,31,94,31,169,31,126,31,12,31,28,31,138,31,248,31,43,31,228,31,235,31,113,31,164,31,163,31,167,31,227,31,227,30,119,31,169,31,40,31,89,31,89,30,75,31,67,31,17,31,38,31,38,30,101,31,45,31,45,30,228,31,228,30,228,29,163,31,163,30,8,31,5,31,129,31,170,31,170,30,55,31,44,31,56,31,230,31,31,31,241,31,241,30,239,31,86,31,168,31,179,31,209,31,103,31,64,31,64,30,252,31,135,31,219,31,104,31,197,31,197,30,10,31,10,30,179,31,36,31,30,31,162,31,162,30,208,31,29,31,179,31,16,31,136,31,83,31,118,31,101,31,31,31,71,31,59,31,63,31,63,30,79,31,79,30,83,31,52,31,3,31,3,30,181,31,65,31,19,31,19,30,19,29,19,28,19,27,14,31,144,31,88,31,88,30,74,31,30,31,151,31,151,30,108,31,49,31,49,30,221,31,221,30,227,31,64,31,183,31,195,31,195,30,249,31,249,30,219,31,242,31,242,30,119,31,119,30,50,31,113,31,55,31,116,31,116,30,7,31,112,31,112,30,112,29,112,28,202,31,154,31,57,31,184,31,184,30,72,31,129,31,160,31,160,30,79,31,241,31,41,31,238,31,73,31,73,30,230,31,118,31,170,31,92,31,92,30,92,29,234,31,182,31,47,31,151,31,219,31,130,31,130,30,206,31,76,31,82,31,29,31,134,31,4,31,91,31,15,31,46,31,111,31,194,31,64,31,132,31,36,31,82,31,168,31,126,31,126,30,205,31,159,31,108,31,95,31,95,30,188,31,188,30,37,31,37,30,124,31,254,31,96,31,49,31,19,31,132,31,142,31,163,31,163,30,112,31,217,31,119,31,237,31,171,31,39,31,220,31,220,30,12,31,198,31,254,31,254,30,214,31,15,31,77,31,153,31,233,31,236,31,41,31,118,31,74,31,74,30,241,31,19,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
