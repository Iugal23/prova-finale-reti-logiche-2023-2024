-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 595;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (85,0,71,0,127,0,122,0,0,0,88,0,0,0,196,0,176,0,0,0,105,0,46,0,113,0,228,0,0,0,26,0,0,0,81,0,16,0,199,0,150,0,74,0,0,0,31,0,147,0,57,0,103,0,100,0,50,0,133,0,245,0,109,0,187,0,43,0,229,0,29,0,0,0,0,0,31,0,14,0,0,0,255,0,109,0,170,0,162,0,52,0,159,0,0,0,0,0,141,0,189,0,239,0,13,0,78,0,40,0,74,0,192,0,255,0,117,0,66,0,159,0,53,0,0,0,202,0,183,0,52,0,75,0,180,0,103,0,62,0,0,0,117,0,247,0,163,0,0,0,148,0,0,0,0,0,111,0,7,0,70,0,193,0,0,0,180,0,146,0,213,0,237,0,225,0,121,0,185,0,244,0,89,0,0,0,0,0,190,0,127,0,80,0,177,0,215,0,23,0,25,0,168,0,242,0,71,0,0,0,222,0,194,0,72,0,191,0,148,0,100,0,99,0,0,0,203,0,156,0,0,0,154,0,33,0,95,0,232,0,239,0,38,0,201,0,200,0,56,0,0,0,0,0,175,0,121,0,46,0,42,0,123,0,0,0,45,0,0,0,0,0,0,0,141,0,128,0,77,0,0,0,0,0,0,0,93,0,215,0,0,0,0,0,190,0,23,0,0,0,201,0,138,0,68,0,48,0,59,0,157,0,211,0,0,0,253,0,240,0,35,0,254,0,120,0,174,0,158,0,0,0,0,0,162,0,65,0,23,0,29,0,167,0,0,0,0,0,27,0,6,0,146,0,0,0,53,0,0,0,232,0,213,0,94,0,247,0,71,0,59,0,0,0,154,0,1,0,0,0,195,0,188,0,185,0,47,0,254,0,22,0,41,0,22,0,106,0,53,0,194,0,124,0,30,0,91,0,76,0,88,0,135,0,0,0,22,0,78,0,246,0,0,0,0,0,155,0,0,0,79,0,70,0,80,0,191,0,0,0,53,0,170,0,145,0,233,0,206,0,0,0,225,0,124,0,111,0,235,0,103,0,138,0,224,0,74,0,175,0,0,0,144,0,0,0,244,0,126,0,118,0,79,0,0,0,222,0,118,0,96,0,0,0,160,0,0,0,7,0,62,0,183,0,181,0,1,0,140,0,182,0,21,0,0,0,139,0,148,0,121,0,191,0,29,0,240,0,218,0,142,0,8,0,53,0,102,0,63,0,220,0,0,0,199,0,27,0,22,0,112,0,0,0,254,0,52,0,253,0,86,0,169,0,87,0,23,0,159,0,159,0,128,0,146,0,225,0,233,0,249,0,225,0,46,0,217,0,154,0,210,0,166,0,0,0,240,0,181,0,0,0,0,0,220,0,0,0,133,0,165,0,0,0,129,0,154,0,44,0,0,0,69,0,155,0,0,0,45,0,156,0,134,0,106,0,43,0,134,0,97,0,0,0,0,0,160,0,0,0,248,0,150,0,26,0,121,0,124,0,179,0,226,0,8,0,118,0,221,0,7,0,244,0,0,0,65,0,0,0,0,0,2,0,0,0,232,0,51,0,0,0,180,0,88,0,0,0,58,0,49,0,144,0,194,0,200,0,0,0,0,0,242,0,0,0,104,0,190,0,186,0,156,0,50,0,155,0,125,0,254,0,230,0,220,0,237,0,195,0,116,0,206,0,151,0,244,0,180,0,190,0,1,0,132,0,248,0,0,0,152,0,112,0,7,0,68,0,89,0,0,0,136,0,89,0,88,0,44,0,109,0,0,0,230,0,185,0,198,0,90,0,58,0,154,0,145,0,209,0,193,0,140,0,125,0,0,0,111,0,175,0,190,0,195,0,99,0,18,0,142,0,0,0,0,0,161,0,0,0,249,0,194,0,120,0,121,0,245,0,0,0,170,0,0,0,0,0,194,0,0,0,0,0,91,0,0,0,0,0,0,0,0,0,194,0,0,0,96,0,186,0,192,0,0,0,58,0,5,0,226,0,213,0,123,0,150,0,101,0,15,0,77,0,245,0,160,0,137,0,188,0,208,0,22,0,0,0,39,0,168,0,79,0,85,0,64,0,162,0,180,0,247,0,153,0,0,0,253,0,145,0,234,0,92,0,237,0,0,0,72,0,0,0,161,0,252,0,72,0,82,0,0,0,208,0,188,0,148,0,198,0,194,0,0,0,231,0,127,0,239,0,195,0,171,0,61,0,215,0,16,0,0,0,111,0,0,0,69,0,250,0,84,0,72,0,0,0,110,0,238,0,84,0,181,0,0,0,0,0,211,0,0,0,175,0,111,0,82,0,0,0,147,0,0,0,248,0,129,0,68,0,78,0,250,0,0,0,0,0,243,0,22,0,0,0,156,0,0,0,141,0,54,0,0,0,0,0,27,0,0,0,235,0,0,0,90,0,61,0,0,0,0,0,24,0,101,0,157,0,0,0,0,0,0,0,206,0,33,0,242,0,65,0,202,0,0,0,0,0,77,0,0,0,0,0,233,0,0,0,2,0,115,0,106,0,128,0,241,0,58,0,0,0,113,0,242,0,17,0,162,0,102,0,123,0,168,0,244,0,0,0,92,0,0,0,10,0,0,0,122,0,161,0,94,0,0,0,0,0,50,0,101,0,179,0,208,0,163,0,31,0,65,0,136,0,0,0,223,0,182,0,21,0,94,0,106,0,0,0);
signal scenario_full  : scenario_type := (85,31,71,31,127,31,122,31,122,30,88,31,88,30,196,31,176,31,176,30,105,31,46,31,113,31,228,31,228,30,26,31,26,30,81,31,16,31,199,31,150,31,74,31,74,30,31,31,147,31,57,31,103,31,100,31,50,31,133,31,245,31,109,31,187,31,43,31,229,31,29,31,29,30,29,29,31,31,14,31,14,30,255,31,109,31,170,31,162,31,52,31,159,31,159,30,159,29,141,31,189,31,239,31,13,31,78,31,40,31,74,31,192,31,255,31,117,31,66,31,159,31,53,31,53,30,202,31,183,31,52,31,75,31,180,31,103,31,62,31,62,30,117,31,247,31,163,31,163,30,148,31,148,30,148,29,111,31,7,31,70,31,193,31,193,30,180,31,146,31,213,31,237,31,225,31,121,31,185,31,244,31,89,31,89,30,89,29,190,31,127,31,80,31,177,31,215,31,23,31,25,31,168,31,242,31,71,31,71,30,222,31,194,31,72,31,191,31,148,31,100,31,99,31,99,30,203,31,156,31,156,30,154,31,33,31,95,31,232,31,239,31,38,31,201,31,200,31,56,31,56,30,56,29,175,31,121,31,46,31,42,31,123,31,123,30,45,31,45,30,45,29,45,28,141,31,128,31,77,31,77,30,77,29,77,28,93,31,215,31,215,30,215,29,190,31,23,31,23,30,201,31,138,31,68,31,48,31,59,31,157,31,211,31,211,30,253,31,240,31,35,31,254,31,120,31,174,31,158,31,158,30,158,29,162,31,65,31,23,31,29,31,167,31,167,30,167,29,27,31,6,31,146,31,146,30,53,31,53,30,232,31,213,31,94,31,247,31,71,31,59,31,59,30,154,31,1,31,1,30,195,31,188,31,185,31,47,31,254,31,22,31,41,31,22,31,106,31,53,31,194,31,124,31,30,31,91,31,76,31,88,31,135,31,135,30,22,31,78,31,246,31,246,30,246,29,155,31,155,30,79,31,70,31,80,31,191,31,191,30,53,31,170,31,145,31,233,31,206,31,206,30,225,31,124,31,111,31,235,31,103,31,138,31,224,31,74,31,175,31,175,30,144,31,144,30,244,31,126,31,118,31,79,31,79,30,222,31,118,31,96,31,96,30,160,31,160,30,7,31,62,31,183,31,181,31,1,31,140,31,182,31,21,31,21,30,139,31,148,31,121,31,191,31,29,31,240,31,218,31,142,31,8,31,53,31,102,31,63,31,220,31,220,30,199,31,27,31,22,31,112,31,112,30,254,31,52,31,253,31,86,31,169,31,87,31,23,31,159,31,159,31,128,31,146,31,225,31,233,31,249,31,225,31,46,31,217,31,154,31,210,31,166,31,166,30,240,31,181,31,181,30,181,29,220,31,220,30,133,31,165,31,165,30,129,31,154,31,44,31,44,30,69,31,155,31,155,30,45,31,156,31,134,31,106,31,43,31,134,31,97,31,97,30,97,29,160,31,160,30,248,31,150,31,26,31,121,31,124,31,179,31,226,31,8,31,118,31,221,31,7,31,244,31,244,30,65,31,65,30,65,29,2,31,2,30,232,31,51,31,51,30,180,31,88,31,88,30,58,31,49,31,144,31,194,31,200,31,200,30,200,29,242,31,242,30,104,31,190,31,186,31,156,31,50,31,155,31,125,31,254,31,230,31,220,31,237,31,195,31,116,31,206,31,151,31,244,31,180,31,190,31,1,31,132,31,248,31,248,30,152,31,112,31,7,31,68,31,89,31,89,30,136,31,89,31,88,31,44,31,109,31,109,30,230,31,185,31,198,31,90,31,58,31,154,31,145,31,209,31,193,31,140,31,125,31,125,30,111,31,175,31,190,31,195,31,99,31,18,31,142,31,142,30,142,29,161,31,161,30,249,31,194,31,120,31,121,31,245,31,245,30,170,31,170,30,170,29,194,31,194,30,194,29,91,31,91,30,91,29,91,28,91,27,194,31,194,30,96,31,186,31,192,31,192,30,58,31,5,31,226,31,213,31,123,31,150,31,101,31,15,31,77,31,245,31,160,31,137,31,188,31,208,31,22,31,22,30,39,31,168,31,79,31,85,31,64,31,162,31,180,31,247,31,153,31,153,30,253,31,145,31,234,31,92,31,237,31,237,30,72,31,72,30,161,31,252,31,72,31,82,31,82,30,208,31,188,31,148,31,198,31,194,31,194,30,231,31,127,31,239,31,195,31,171,31,61,31,215,31,16,31,16,30,111,31,111,30,69,31,250,31,84,31,72,31,72,30,110,31,238,31,84,31,181,31,181,30,181,29,211,31,211,30,175,31,111,31,82,31,82,30,147,31,147,30,248,31,129,31,68,31,78,31,250,31,250,30,250,29,243,31,22,31,22,30,156,31,156,30,141,31,54,31,54,30,54,29,27,31,27,30,235,31,235,30,90,31,61,31,61,30,61,29,24,31,101,31,157,31,157,30,157,29,157,28,206,31,33,31,242,31,65,31,202,31,202,30,202,29,77,31,77,30,77,29,233,31,233,30,2,31,115,31,106,31,128,31,241,31,58,31,58,30,113,31,242,31,17,31,162,31,102,31,123,31,168,31,244,31,244,30,92,31,92,30,10,31,10,30,122,31,161,31,94,31,94,30,94,29,50,31,101,31,179,31,208,31,163,31,31,31,65,31,136,31,136,30,223,31,182,31,21,31,94,31,106,31,106,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
