-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 641;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (168,0,255,0,172,0,150,0,234,0,0,0,128,0,62,0,105,0,221,0,0,0,183,0,254,0,208,0,183,0,134,0,0,0,25,0,6,0,37,0,138,0,42,0,224,0,0,0,17,0,0,0,0,0,212,0,128,0,0,0,2,0,92,0,132,0,179,0,186,0,205,0,62,0,104,0,79,0,0,0,179,0,226,0,192,0,81,0,5,0,75,0,0,0,0,0,5,0,20,0,173,0,232,0,197,0,126,0,190,0,118,0,125,0,0,0,234,0,52,0,207,0,7,0,111,0,143,0,113,0,20,0,100,0,137,0,88,0,15,0,99,0,198,0,41,0,164,0,75,0,76,0,133,0,147,0,0,0,33,0,246,0,0,0,89,0,166,0,106,0,244,0,0,0,163,0,134,0,139,0,170,0,0,0,107,0,228,0,0,0,228,0,0,0,0,0,15,0,0,0,178,0,0,0,227,0,123,0,222,0,0,0,126,0,108,0,241,0,19,0,39,0,36,0,0,0,111,0,190,0,222,0,112,0,58,0,0,0,123,0,21,0,127,0,151,0,76,0,66,0,11,0,151,0,0,0,117,0,38,0,0,0,28,0,0,0,75,0,157,0,0,0,0,0,179,0,174,0,25,0,14,0,177,0,155,0,224,0,41,0,86,0,158,0,24,0,180,0,93,0,0,0,31,0,175,0,0,0,62,0,0,0,54,0,204,0,101,0,0,0,125,0,254,0,89,0,0,0,93,0,166,0,232,0,227,0,110,0,0,0,223,0,43,0,16,0,0,0,169,0,73,0,196,0,231,0,175,0,0,0,0,0,169,0,36,0,6,0,243,0,30,0,18,0,221,0,1,0,0,0,63,0,0,0,178,0,211,0,225,0,187,0,0,0,176,0,211,0,39,0,67,0,109,0,150,0,82,0,50,0,4,0,148,0,63,0,191,0,38,0,171,0,7,0,5,0,188,0,35,0,120,0,200,0,0,0,89,0,1,0,231,0,0,0,100,0,195,0,99,0,160,0,234,0,2,0,64,0,251,0,163,0,103,0,0,0,57,0,160,0,175,0,16,0,13,0,0,0,0,0,11,0,214,0,203,0,0,0,91,0,194,0,145,0,255,0,0,0,72,0,20,0,61,0,0,0,198,0,167,0,152,0,130,0,229,0,0,0,1,0,0,0,0,0,49,0,177,0,173,0,44,0,60,0,250,0,2,0,226,0,0,0,135,0,247,0,125,0,157,0,234,0,106,0,197,0,61,0,203,0,139,0,175,0,0,0,145,0,207,0,0,0,227,0,116,0,213,0,0,0,107,0,25,0,0,0,141,0,180,0,241,0,77,0,169,0,50,0,0,0,183,0,253,0,0,0,32,0,145,0,91,0,238,0,165,0,206,0,134,0,62,0,59,0,62,0,79,0,111,0,121,0,12,0,107,0,6,0,0,0,207,0,194,0,172,0,0,0,169,0,0,0,112,0,46,0,96,0,169,0,21,0,199,0,0,0,160,0,6,0,118,0,0,0,29,0,151,0,81,0,112,0,63,0,4,0,0,0,118,0,162,0,107,0,178,0,203,0,134,0,195,0,220,0,9,0,103,0,60,0,29,0,23,0,177,0,209,0,0,0,0,0,122,0,0,0,232,0,121,0,35,0,220,0,58,0,195,0,125,0,237,0,116,0,20,0,0,0,161,0,17,0,0,0,173,0,131,0,10,0,166,0,214,0,54,0,153,0,74,0,114,0,105,0,108,0,128,0,0,0,0,0,0,0,105,0,176,0,0,0,72,0,36,0,165,0,135,0,48,0,131,0,40,0,0,0,93,0,0,0,55,0,39,0,0,0,175,0,221,0,37,0,227,0,183,0,117,0,140,0,0,0,196,0,0,0,0,0,0,0,75,0,0,0,0,0,212,0,127,0,218,0,0,0,0,0,154,0,241,0,127,0,121,0,68,0,113,0,210,0,0,0,70,0,178,0,204,0,73,0,0,0,135,0,2,0,84,0,3,0,107,0,123,0,160,0,221,0,0,0,179,0,35,0,56,0,57,0,152,0,183,0,165,0,130,0,0,0,243,0,66,0,171,0,16,0,53,0,106,0,230,0,214,0,54,0,183,0,161,0,39,0,34,0,95,0,183,0,0,0,237,0,0,0,106,0,0,0,177,0,143,0,0,0,59,0,71,0,38,0,152,0,117,0,212,0,144,0,216,0,238,0,0,0,115,0,178,0,243,0,210,0,183,0,190,0,3,0,0,0,136,0,134,0,152,0,113,0,0,0,159,0,0,0,175,0,214,0,92,0,146,0,182,0,232,0,0,0,198,0,0,0,149,0,154,0,243,0,116,0,62,0,0,0,86,0,116,0,0,0,0,0,21,0,0,0,19,0,152,0,136,0,186,0,232,0,123,0,252,0,0,0,123,0,24,0,0,0,115,0,79,0,91,0,170,0,116,0,147,0,83,0,78,0,0,0,0,0,120,0,15,0,0,0,16,0,206,0,212,0,0,0,82,0,252,0,252,0,149,0,236,0,0,0,171,0,82,0,117,0,150,0,0,0,206,0,63,0,111,0,170,0,174,0,47,0,110,0,200,0,251,0,0,0,163,0,151,0,88,0,125,0,97,0,18,0,172,0,60,0,132,0,0,0,0,0,0,0,151,0,0,0,0,0,108,0,30,0,5,0,191,0,45,0,0,0,15,0,127,0,224,0,104,0,72,0,93,0,125,0,136,0,180,0,38,0,155,0,13,0,0,0,140,0,142,0,23,0,255,0,164,0,185,0,0,0,0,0,131,0,234,0,80,0,111,0,220,0,111,0,141,0,187,0,94,0,60,0,39,0,211,0,132,0,40,0,120,0,58,0,95,0,228,0,182,0,168,0,190,0,55,0);
signal scenario_full  : scenario_type := (168,31,255,31,172,31,150,31,234,31,234,30,128,31,62,31,105,31,221,31,221,30,183,31,254,31,208,31,183,31,134,31,134,30,25,31,6,31,37,31,138,31,42,31,224,31,224,30,17,31,17,30,17,29,212,31,128,31,128,30,2,31,92,31,132,31,179,31,186,31,205,31,62,31,104,31,79,31,79,30,179,31,226,31,192,31,81,31,5,31,75,31,75,30,75,29,5,31,20,31,173,31,232,31,197,31,126,31,190,31,118,31,125,31,125,30,234,31,52,31,207,31,7,31,111,31,143,31,113,31,20,31,100,31,137,31,88,31,15,31,99,31,198,31,41,31,164,31,75,31,76,31,133,31,147,31,147,30,33,31,246,31,246,30,89,31,166,31,106,31,244,31,244,30,163,31,134,31,139,31,170,31,170,30,107,31,228,31,228,30,228,31,228,30,228,29,15,31,15,30,178,31,178,30,227,31,123,31,222,31,222,30,126,31,108,31,241,31,19,31,39,31,36,31,36,30,111,31,190,31,222,31,112,31,58,31,58,30,123,31,21,31,127,31,151,31,76,31,66,31,11,31,151,31,151,30,117,31,38,31,38,30,28,31,28,30,75,31,157,31,157,30,157,29,179,31,174,31,25,31,14,31,177,31,155,31,224,31,41,31,86,31,158,31,24,31,180,31,93,31,93,30,31,31,175,31,175,30,62,31,62,30,54,31,204,31,101,31,101,30,125,31,254,31,89,31,89,30,93,31,166,31,232,31,227,31,110,31,110,30,223,31,43,31,16,31,16,30,169,31,73,31,196,31,231,31,175,31,175,30,175,29,169,31,36,31,6,31,243,31,30,31,18,31,221,31,1,31,1,30,63,31,63,30,178,31,211,31,225,31,187,31,187,30,176,31,211,31,39,31,67,31,109,31,150,31,82,31,50,31,4,31,148,31,63,31,191,31,38,31,171,31,7,31,5,31,188,31,35,31,120,31,200,31,200,30,89,31,1,31,231,31,231,30,100,31,195,31,99,31,160,31,234,31,2,31,64,31,251,31,163,31,103,31,103,30,57,31,160,31,175,31,16,31,13,31,13,30,13,29,11,31,214,31,203,31,203,30,91,31,194,31,145,31,255,31,255,30,72,31,20,31,61,31,61,30,198,31,167,31,152,31,130,31,229,31,229,30,1,31,1,30,1,29,49,31,177,31,173,31,44,31,60,31,250,31,2,31,226,31,226,30,135,31,247,31,125,31,157,31,234,31,106,31,197,31,61,31,203,31,139,31,175,31,175,30,145,31,207,31,207,30,227,31,116,31,213,31,213,30,107,31,25,31,25,30,141,31,180,31,241,31,77,31,169,31,50,31,50,30,183,31,253,31,253,30,32,31,145,31,91,31,238,31,165,31,206,31,134,31,62,31,59,31,62,31,79,31,111,31,121,31,12,31,107,31,6,31,6,30,207,31,194,31,172,31,172,30,169,31,169,30,112,31,46,31,96,31,169,31,21,31,199,31,199,30,160,31,6,31,118,31,118,30,29,31,151,31,81,31,112,31,63,31,4,31,4,30,118,31,162,31,107,31,178,31,203,31,134,31,195,31,220,31,9,31,103,31,60,31,29,31,23,31,177,31,209,31,209,30,209,29,122,31,122,30,232,31,121,31,35,31,220,31,58,31,195,31,125,31,237,31,116,31,20,31,20,30,161,31,17,31,17,30,173,31,131,31,10,31,166,31,214,31,54,31,153,31,74,31,114,31,105,31,108,31,128,31,128,30,128,29,128,28,105,31,176,31,176,30,72,31,36,31,165,31,135,31,48,31,131,31,40,31,40,30,93,31,93,30,55,31,39,31,39,30,175,31,221,31,37,31,227,31,183,31,117,31,140,31,140,30,196,31,196,30,196,29,196,28,75,31,75,30,75,29,212,31,127,31,218,31,218,30,218,29,154,31,241,31,127,31,121,31,68,31,113,31,210,31,210,30,70,31,178,31,204,31,73,31,73,30,135,31,2,31,84,31,3,31,107,31,123,31,160,31,221,31,221,30,179,31,35,31,56,31,57,31,152,31,183,31,165,31,130,31,130,30,243,31,66,31,171,31,16,31,53,31,106,31,230,31,214,31,54,31,183,31,161,31,39,31,34,31,95,31,183,31,183,30,237,31,237,30,106,31,106,30,177,31,143,31,143,30,59,31,71,31,38,31,152,31,117,31,212,31,144,31,216,31,238,31,238,30,115,31,178,31,243,31,210,31,183,31,190,31,3,31,3,30,136,31,134,31,152,31,113,31,113,30,159,31,159,30,175,31,214,31,92,31,146,31,182,31,232,31,232,30,198,31,198,30,149,31,154,31,243,31,116,31,62,31,62,30,86,31,116,31,116,30,116,29,21,31,21,30,19,31,152,31,136,31,186,31,232,31,123,31,252,31,252,30,123,31,24,31,24,30,115,31,79,31,91,31,170,31,116,31,147,31,83,31,78,31,78,30,78,29,120,31,15,31,15,30,16,31,206,31,212,31,212,30,82,31,252,31,252,31,149,31,236,31,236,30,171,31,82,31,117,31,150,31,150,30,206,31,63,31,111,31,170,31,174,31,47,31,110,31,200,31,251,31,251,30,163,31,151,31,88,31,125,31,97,31,18,31,172,31,60,31,132,31,132,30,132,29,132,28,151,31,151,30,151,29,108,31,30,31,5,31,191,31,45,31,45,30,15,31,127,31,224,31,104,31,72,31,93,31,125,31,136,31,180,31,38,31,155,31,13,31,13,30,140,31,142,31,23,31,255,31,164,31,185,31,185,30,185,29,131,31,234,31,80,31,111,31,220,31,111,31,141,31,187,31,94,31,60,31,39,31,211,31,132,31,40,31,120,31,58,31,95,31,228,31,182,31,168,31,190,31,55,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
