-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 772;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,245,0,90,0,0,0,0,0,0,0,174,0,0,0,44,0,25,0,163,0,177,0,141,0,251,0,2,0,32,0,168,0,0,0,227,0,0,0,145,0,80,0,208,0,105,0,72,0,234,0,0,0,174,0,174,0,156,0,0,0,0,0,236,0,62,0,0,0,217,0,0,0,37,0,0,0,12,0,146,0,133,0,173,0,34,0,22,0,105,0,182,0,199,0,157,0,4,0,0,0,0,0,18,0,185,0,0,0,0,0,137,0,208,0,250,0,0,0,16,0,124,0,0,0,29,0,138,0,67,0,38,0,145,0,203,0,21,0,52,0,88,0,0,0,236,0,0,0,195,0,167,0,0,0,0,0,175,0,0,0,196,0,0,0,99,0,27,0,22,0,142,0,111,0,241,0,31,0,53,0,165,0,239,0,75,0,71,0,72,0,21,0,26,0,21,0,184,0,159,0,53,0,0,0,4,0,96,0,0,0,241,0,0,0,126,0,14,0,202,0,212,0,9,0,156,0,0,0,26,0,247,0,139,0,7,0,106,0,181,0,26,0,0,0,235,0,126,0,13,0,82,0,0,0,227,0,124,0,239,0,0,0,0,0,236,0,0,0,209,0,44,0,137,0,0,0,0,0,39,0,74,0,131,0,245,0,20,0,14,0,241,0,0,0,0,0,117,0,194,0,6,0,0,0,106,0,0,0,127,0,191,0,0,0,46,0,0,0,10,0,153,0,0,0,0,0,210,0,125,0,90,0,101,0,1,0,0,0,0,0,223,0,2,0,214,0,0,0,22,0,178,0,36,0,28,0,242,0,128,0,121,0,0,0,0,0,0,0,31,0,230,0,0,0,0,0,183,0,228,0,202,0,143,0,0,0,152,0,229,0,0,0,26,0,245,0,0,0,73,0,247,0,92,0,20,0,93,0,0,0,24,0,220,0,0,0,52,0,188,0,0,0,33,0,226,0,152,0,251,0,154,0,172,0,191,0,108,0,31,0,229,0,51,0,150,0,146,0,94,0,22,0,0,0,47,0,10,0,143,0,43,0,101,0,80,0,251,0,200,0,161,0,216,0,194,0,194,0,207,0,115,0,190,0,100,0,184,0,154,0,0,0,0,0,0,0,208,0,0,0,70,0,215,0,224,0,0,0,60,0,48,0,26,0,0,0,56,0,24,0,28,0,8,0,89,0,72,0,129,0,83,0,32,0,11,0,50,0,0,0,225,0,194,0,27,0,81,0,228,0,114,0,117,0,159,0,0,0,69,0,0,0,0,0,57,0,251,0,173,0,46,0,0,0,159,0,60,0,0,0,223,0,214,0,46,0,0,0,83,0,187,0,250,0,0,0,178,0,177,0,31,0,170,0,223,0,113,0,244,0,204,0,156,0,209,0,249,0,105,0,124,0,53,0,177,0,64,0,0,0,212,0,225,0,160,0,157,0,175,0,229,0,0,0,126,0,13,0,188,0,248,0,117,0,0,0,0,0,0,0,76,0,6,0,118,0,0,0,3,0,175,0,132,0,192,0,161,0,218,0,82,0,78,0,25,0,65,0,101,0,137,0,0,0,0,0,162,0,0,0,13,0,0,0,0,0,0,0,202,0,167,0,0,0,10,0,99,0,80,0,135,0,69,0,0,0,39,0,181,0,48,0,131,0,18,0,6,0,2,0,0,0,23,0,0,0,0,0,42,0,0,0,0,0,172,0,173,0,0,0,149,0,93,0,90,0,0,0,33,0,225,0,106,0,179,0,0,0,44,0,55,0,104,0,26,0,175,0,57,0,0,0,217,0,160,0,62,0,207,0,67,0,0,0,0,0,248,0,2,0,0,0,53,0,0,0,0,0,103,0,0,0,205,0,21,0,157,0,206,0,90,0,84,0,193,0,238,0,193,0,0,0,0,0,0,0,125,0,173,0,11,0,130,0,168,0,0,0,169,0,185,0,13,0,47,0,206,0,13,0,0,0,48,0,169,0,97,0,212,0,165,0,0,0,208,0,118,0,249,0,147,0,222,0,0,0,0,0,114,0,15,0,211,0,104,0,32,0,117,0,135,0,37,0,123,0,224,0,127,0,221,0,0,0,1,0,199,0,237,0,209,0,0,0,0,0,0,0,229,0,233,0,33,0,75,0,42,0,247,0,250,0,15,0,147,0,0,0,99,0,129,0,212,0,63,0,99,0,117,0,100,0,98,0,167,0,13,0,249,0,48,0,11,0,168,0,27,0,109,0,0,0,172,0,176,0,234,0,106,0,2,0,143,0,0,0,113,0,0,0,0,0,0,0,237,0,37,0,0,0,239,0,127,0,9,0,102,0,46,0,64,0,181,0,122,0,252,0,98,0,62,0,82,0,0,0,125,0,0,0,253,0,31,0,54,0,0,0,100,0,76,0,51,0,66,0,213,0,33,0,58,0,0,0,227,0,203,0,14,0,157,0,0,0,130,0,9,0,187,0,204,0,0,0,254,0,34,0,128,0,253,0,176,0,0,0,196,0,0,0,229,0,247,0,126,0,18,0,0,0,139,0,172,0,155,0,57,0,0,0,0,0,204,0,88,0,222,0,51,0,88,0,34,0,242,0,172,0,0,0,42,0,114,0,207,0,90,0,92,0,178,0,183,0,251,0,36,0,0,0,0,0,205,0,55,0,41,0,190,0,221,0,124,0,0,0,111,0,129,0,105,0,11,0,0,0,126,0,0,0,145,0,23,0,0,0,0,0,10,0,46,0,143,0,11,0,21,0,96,0,195,0,186,0,43,0,0,0,6,0,0,0,0,0,147,0,180,0,0,0,0,0,1,0,123,0,54,0,9,0,0,0,197,0,202,0,149,0,4,0,99,0,192,0,23,0,6,0,106,0,250,0,109,0,182,0,127,0,0,0,227,0,17,0,223,0,221,0,159,0,87,0,0,0,51,0,0,0,41,0,231,0,0,0,80,0,46,0,44,0,130,0,75,0,230,0,81,0,0,0,15,0,196,0,150,0,206,0,0,0,162,0,159,0,0,0,224,0,0,0,192,0,5,0,96,0,160,0,0,0,239,0,2,0,234,0,0,0,206,0,18,0,0,0,232,0,3,0,171,0,240,0,32,0,226,0,150,0,134,0,237,0,214,0,1,0,205,0,1,0,117,0,28,0,1,0,135,0,0,0,0,0,229,0,0,0,137,0,92,0,0,0,100,0,0,0,254,0,103,0,0,0,147,0,86,0,0,0,99,0,1,0,0,0,36,0,0,0,163,0,131,0,174,0,171,0,215,0,139,0,130,0,97,0,54,0,105,0,118,0,201,0,186,0,26,0,119,0,0,0,37,0,155,0,61,0,0,0,157,0,0,0,143,0,170,0,58,0,198,0,180,0,189,0,38,0,118,0,0,0,28,0,60,0,77,0,183,0,19,0,56,0,192,0,170,0,198,0,147,0,237,0,11,0,0,0,86,0,149,0,213,0,248,0,117,0,61,0,53,0);
signal scenario_full  : scenario_type := (0,0,0,0,245,31,90,31,90,30,90,29,90,28,174,31,174,30,44,31,25,31,163,31,177,31,141,31,251,31,2,31,32,31,168,31,168,30,227,31,227,30,145,31,80,31,208,31,105,31,72,31,234,31,234,30,174,31,174,31,156,31,156,30,156,29,236,31,62,31,62,30,217,31,217,30,37,31,37,30,12,31,146,31,133,31,173,31,34,31,22,31,105,31,182,31,199,31,157,31,4,31,4,30,4,29,18,31,185,31,185,30,185,29,137,31,208,31,250,31,250,30,16,31,124,31,124,30,29,31,138,31,67,31,38,31,145,31,203,31,21,31,52,31,88,31,88,30,236,31,236,30,195,31,167,31,167,30,167,29,175,31,175,30,196,31,196,30,99,31,27,31,22,31,142,31,111,31,241,31,31,31,53,31,165,31,239,31,75,31,71,31,72,31,21,31,26,31,21,31,184,31,159,31,53,31,53,30,4,31,96,31,96,30,241,31,241,30,126,31,14,31,202,31,212,31,9,31,156,31,156,30,26,31,247,31,139,31,7,31,106,31,181,31,26,31,26,30,235,31,126,31,13,31,82,31,82,30,227,31,124,31,239,31,239,30,239,29,236,31,236,30,209,31,44,31,137,31,137,30,137,29,39,31,74,31,131,31,245,31,20,31,14,31,241,31,241,30,241,29,117,31,194,31,6,31,6,30,106,31,106,30,127,31,191,31,191,30,46,31,46,30,10,31,153,31,153,30,153,29,210,31,125,31,90,31,101,31,1,31,1,30,1,29,223,31,2,31,214,31,214,30,22,31,178,31,36,31,28,31,242,31,128,31,121,31,121,30,121,29,121,28,31,31,230,31,230,30,230,29,183,31,228,31,202,31,143,31,143,30,152,31,229,31,229,30,26,31,245,31,245,30,73,31,247,31,92,31,20,31,93,31,93,30,24,31,220,31,220,30,52,31,188,31,188,30,33,31,226,31,152,31,251,31,154,31,172,31,191,31,108,31,31,31,229,31,51,31,150,31,146,31,94,31,22,31,22,30,47,31,10,31,143,31,43,31,101,31,80,31,251,31,200,31,161,31,216,31,194,31,194,31,207,31,115,31,190,31,100,31,184,31,154,31,154,30,154,29,154,28,208,31,208,30,70,31,215,31,224,31,224,30,60,31,48,31,26,31,26,30,56,31,24,31,28,31,8,31,89,31,72,31,129,31,83,31,32,31,11,31,50,31,50,30,225,31,194,31,27,31,81,31,228,31,114,31,117,31,159,31,159,30,69,31,69,30,69,29,57,31,251,31,173,31,46,31,46,30,159,31,60,31,60,30,223,31,214,31,46,31,46,30,83,31,187,31,250,31,250,30,178,31,177,31,31,31,170,31,223,31,113,31,244,31,204,31,156,31,209,31,249,31,105,31,124,31,53,31,177,31,64,31,64,30,212,31,225,31,160,31,157,31,175,31,229,31,229,30,126,31,13,31,188,31,248,31,117,31,117,30,117,29,117,28,76,31,6,31,118,31,118,30,3,31,175,31,132,31,192,31,161,31,218,31,82,31,78,31,25,31,65,31,101,31,137,31,137,30,137,29,162,31,162,30,13,31,13,30,13,29,13,28,202,31,167,31,167,30,10,31,99,31,80,31,135,31,69,31,69,30,39,31,181,31,48,31,131,31,18,31,6,31,2,31,2,30,23,31,23,30,23,29,42,31,42,30,42,29,172,31,173,31,173,30,149,31,93,31,90,31,90,30,33,31,225,31,106,31,179,31,179,30,44,31,55,31,104,31,26,31,175,31,57,31,57,30,217,31,160,31,62,31,207,31,67,31,67,30,67,29,248,31,2,31,2,30,53,31,53,30,53,29,103,31,103,30,205,31,21,31,157,31,206,31,90,31,84,31,193,31,238,31,193,31,193,30,193,29,193,28,125,31,173,31,11,31,130,31,168,31,168,30,169,31,185,31,13,31,47,31,206,31,13,31,13,30,48,31,169,31,97,31,212,31,165,31,165,30,208,31,118,31,249,31,147,31,222,31,222,30,222,29,114,31,15,31,211,31,104,31,32,31,117,31,135,31,37,31,123,31,224,31,127,31,221,31,221,30,1,31,199,31,237,31,209,31,209,30,209,29,209,28,229,31,233,31,33,31,75,31,42,31,247,31,250,31,15,31,147,31,147,30,99,31,129,31,212,31,63,31,99,31,117,31,100,31,98,31,167,31,13,31,249,31,48,31,11,31,168,31,27,31,109,31,109,30,172,31,176,31,234,31,106,31,2,31,143,31,143,30,113,31,113,30,113,29,113,28,237,31,37,31,37,30,239,31,127,31,9,31,102,31,46,31,64,31,181,31,122,31,252,31,98,31,62,31,82,31,82,30,125,31,125,30,253,31,31,31,54,31,54,30,100,31,76,31,51,31,66,31,213,31,33,31,58,31,58,30,227,31,203,31,14,31,157,31,157,30,130,31,9,31,187,31,204,31,204,30,254,31,34,31,128,31,253,31,176,31,176,30,196,31,196,30,229,31,247,31,126,31,18,31,18,30,139,31,172,31,155,31,57,31,57,30,57,29,204,31,88,31,222,31,51,31,88,31,34,31,242,31,172,31,172,30,42,31,114,31,207,31,90,31,92,31,178,31,183,31,251,31,36,31,36,30,36,29,205,31,55,31,41,31,190,31,221,31,124,31,124,30,111,31,129,31,105,31,11,31,11,30,126,31,126,30,145,31,23,31,23,30,23,29,10,31,46,31,143,31,11,31,21,31,96,31,195,31,186,31,43,31,43,30,6,31,6,30,6,29,147,31,180,31,180,30,180,29,1,31,123,31,54,31,9,31,9,30,197,31,202,31,149,31,4,31,99,31,192,31,23,31,6,31,106,31,250,31,109,31,182,31,127,31,127,30,227,31,17,31,223,31,221,31,159,31,87,31,87,30,51,31,51,30,41,31,231,31,231,30,80,31,46,31,44,31,130,31,75,31,230,31,81,31,81,30,15,31,196,31,150,31,206,31,206,30,162,31,159,31,159,30,224,31,224,30,192,31,5,31,96,31,160,31,160,30,239,31,2,31,234,31,234,30,206,31,18,31,18,30,232,31,3,31,171,31,240,31,32,31,226,31,150,31,134,31,237,31,214,31,1,31,205,31,1,31,117,31,28,31,1,31,135,31,135,30,135,29,229,31,229,30,137,31,92,31,92,30,100,31,100,30,254,31,103,31,103,30,147,31,86,31,86,30,99,31,1,31,1,30,36,31,36,30,163,31,131,31,174,31,171,31,215,31,139,31,130,31,97,31,54,31,105,31,118,31,201,31,186,31,26,31,119,31,119,30,37,31,155,31,61,31,61,30,157,31,157,30,143,31,170,31,58,31,198,31,180,31,189,31,38,31,118,31,118,30,28,31,60,31,77,31,183,31,19,31,56,31,192,31,170,31,198,31,147,31,237,31,11,31,11,30,86,31,149,31,213,31,248,31,117,31,61,31,53,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
