-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_318 is
end project_tb_318;

architecture project_tb_arch_318 of project_tb_318 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 629;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (96,0,46,0,77,0,118,0,115,0,235,0,30,0,0,0,75,0,47,0,0,0,69,0,12,0,189,0,124,0,239,0,0,0,113,0,15,0,224,0,0,0,105,0,0,0,219,0,15,0,84,0,91,0,49,0,0,0,115,0,7,0,241,0,7,0,87,0,54,0,198,0,130,0,227,0,0,0,0,0,94,0,19,0,251,0,172,0,141,0,96,0,216,0,0,0,19,0,0,0,107,0,0,0,56,0,42,0,223,0,132,0,0,0,51,0,209,0,90,0,116,0,180,0,43,0,96,0,0,0,139,0,10,0,57,0,48,0,53,0,243,0,10,0,0,0,240,0,108,0,194,0,112,0,0,0,151,0,69,0,0,0,0,0,43,0,161,0,76,0,252,0,16,0,41,0,110,0,137,0,0,0,0,0,112,0,0,0,121,0,98,0,127,0,183,0,57,0,247,0,195,0,0,0,185,0,234,0,0,0,98,0,31,0,7,0,183,0,115,0,207,0,210,0,31,0,104,0,212,0,178,0,94,0,248,0,134,0,194,0,194,0,56,0,178,0,70,0,0,0,120,0,90,0,188,0,211,0,19,0,67,0,227,0,0,0,7,0,92,0,42,0,21,0,0,0,0,0,55,0,0,0,238,0,202,0,65,0,201,0,197,0,206,0,213,0,154,0,137,0,72,0,181,0,0,0,0,0,0,0,207,0,5,0,172,0,34,0,0,0,92,0,40,0,126,0,214,0,0,0,0,0,0,0,147,0,0,0,136,0,122,0,166,0,246,0,240,0,158,0,9,0,150,0,131,0,57,0,74,0,104,0,21,0,0,0,77,0,132,0,10,0,57,0,253,0,40,0,63,0,140,0,93,0,22,0,101,0,227,0,0,0,0,0,203,0,155,0,0,0,218,0,182,0,39,0,61,0,8,0,188,0,196,0,162,0,116,0,46,0,217,0,86,0,0,0,0,0,0,0,202,0,28,0,186,0,6,0,88,0,0,0,0,0,45,0,104,0,49,0,168,0,143,0,200,0,238,0,0,0,67,0,0,0,255,0,0,0,187,0,230,0,24,0,0,0,123,0,225,0,17,0,2,0,0,0,0,0,212,0,136,0,104,0,188,0,95,0,220,0,215,0,124,0,0,0,0,0,73,0,241,0,0,0,97,0,13,0,111,0,0,0,97,0,128,0,0,0,153,0,104,0,146,0,102,0,77,0,0,0,173,0,84,0,113,0,99,0,0,0,0,0,10,0,84,0,23,0,133,0,2,0,189,0,204,0,154,0,0,0,55,0,99,0,76,0,57,0,114,0,229,0,211,0,199,0,201,0,240,0,201,0,195,0,141,0,241,0,177,0,160,0,42,0,74,0,240,0,144,0,0,0,177,0,0,0,76,0,215,0,235,0,14,0,0,0,106,0,79,0,0,0,200,0,0,0,223,0,0,0,255,0,89,0,112,0,0,0,246,0,9,0,28,0,230,0,41,0,89,0,38,0,17,0,147,0,14,0,0,0,58,0,183,0,0,0,167,0,0,0,253,0,149,0,0,0,108,0,132,0,136,0,17,0,180,0,0,0,90,0,0,0,131,0,0,0,211,0,0,0,208,0,94,0,172,0,71,0,0,0,149,0,14,0,177,0,202,0,223,0,0,0,47,0,199,0,72,0,231,0,128,0,19,0,249,0,0,0,55,0,127,0,37,0,135,0,167,0,142,0,223,0,169,0,4,0,0,0,0,0,108,0,0,0,243,0,226,0,213,0,199,0,0,0,244,0,204,0,210,0,58,0,241,0,73,0,0,0,235,0,118,0,56,0,223,0,0,0,154,0,218,0,16,0,207,0,117,0,159,0,191,0,0,0,222,0,220,0,20,0,115,0,187,0,125,0,72,0,0,0,56,0,242,0,0,0,172,0,166,0,102,0,0,0,55,0,36,0,35,0,0,0,11,0,226,0,101,0,56,0,0,0,190,0,0,0,0,0,3,0,144,0,39,0,178,0,207,0,87,0,196,0,153,0,22,0,239,0,16,0,190,0,0,0,0,0,207,0,200,0,218,0,55,0,246,0,126,0,245,0,0,0,177,0,93,0,100,0,91,0,230,0,32,0,108,0,237,0,0,0,250,0,0,0,170,0,0,0,197,0,143,0,10,0,0,0,0,0,163,0,85,0,62,0,48,0,155,0,159,0,153,0,51,0,111,0,84,0,171,0,0,0,0,0,142,0,124,0,194,0,15,0,134,0,194,0,87,0,110,0,131,0,147,0,56,0,133,0,3,0,116,0,0,0,31,0,116,0,197,0,147,0,207,0,36,0,0,0,185,0,166,0,169,0,235,0,0,0,239,0,78,0,105,0,0,0,31,0,12,0,100,0,101,0,0,0,111,0,0,0,149,0,13,0,0,0,192,0,128,0,0,0,0,0,109,0,0,0,0,0,109,0,0,0,239,0,192,0,164,0,239,0,179,0,2,0,109,0,0,0,0,0,142,0,31,0,195,0,0,0,21,0,82,0,0,0,159,0,128,0,183,0,0,0,196,0,0,0,212,0,34,0,154,0,2,0,94,0,20,0,106,0,14,0,17,0,38,0,180,0,217,0,0,0,233,0,49,0,0,0,0,0,0,0,155,0,215,0,173,0,217,0,74,0,51,0,128,0,119,0,251,0,99,0,0,0,93,0,0,0,0,0,173,0,120,0,250,0,0,0,0,0,131,0,225,0,135,0,54,0,0,0,103,0,106,0,128,0,27,0,101,0,139,0,144,0,182,0,188,0,237,0,0,0,0,0,136,0,23,0,138,0,126,0,0,0,40,0,0,0,0,0,80,0,123,0,0,0);
signal scenario_full  : scenario_type := (96,31,46,31,77,31,118,31,115,31,235,31,30,31,30,30,75,31,47,31,47,30,69,31,12,31,189,31,124,31,239,31,239,30,113,31,15,31,224,31,224,30,105,31,105,30,219,31,15,31,84,31,91,31,49,31,49,30,115,31,7,31,241,31,7,31,87,31,54,31,198,31,130,31,227,31,227,30,227,29,94,31,19,31,251,31,172,31,141,31,96,31,216,31,216,30,19,31,19,30,107,31,107,30,56,31,42,31,223,31,132,31,132,30,51,31,209,31,90,31,116,31,180,31,43,31,96,31,96,30,139,31,10,31,57,31,48,31,53,31,243,31,10,31,10,30,240,31,108,31,194,31,112,31,112,30,151,31,69,31,69,30,69,29,43,31,161,31,76,31,252,31,16,31,41,31,110,31,137,31,137,30,137,29,112,31,112,30,121,31,98,31,127,31,183,31,57,31,247,31,195,31,195,30,185,31,234,31,234,30,98,31,31,31,7,31,183,31,115,31,207,31,210,31,31,31,104,31,212,31,178,31,94,31,248,31,134,31,194,31,194,31,56,31,178,31,70,31,70,30,120,31,90,31,188,31,211,31,19,31,67,31,227,31,227,30,7,31,92,31,42,31,21,31,21,30,21,29,55,31,55,30,238,31,202,31,65,31,201,31,197,31,206,31,213,31,154,31,137,31,72,31,181,31,181,30,181,29,181,28,207,31,5,31,172,31,34,31,34,30,92,31,40,31,126,31,214,31,214,30,214,29,214,28,147,31,147,30,136,31,122,31,166,31,246,31,240,31,158,31,9,31,150,31,131,31,57,31,74,31,104,31,21,31,21,30,77,31,132,31,10,31,57,31,253,31,40,31,63,31,140,31,93,31,22,31,101,31,227,31,227,30,227,29,203,31,155,31,155,30,218,31,182,31,39,31,61,31,8,31,188,31,196,31,162,31,116,31,46,31,217,31,86,31,86,30,86,29,86,28,202,31,28,31,186,31,6,31,88,31,88,30,88,29,45,31,104,31,49,31,168,31,143,31,200,31,238,31,238,30,67,31,67,30,255,31,255,30,187,31,230,31,24,31,24,30,123,31,225,31,17,31,2,31,2,30,2,29,212,31,136,31,104,31,188,31,95,31,220,31,215,31,124,31,124,30,124,29,73,31,241,31,241,30,97,31,13,31,111,31,111,30,97,31,128,31,128,30,153,31,104,31,146,31,102,31,77,31,77,30,173,31,84,31,113,31,99,31,99,30,99,29,10,31,84,31,23,31,133,31,2,31,189,31,204,31,154,31,154,30,55,31,99,31,76,31,57,31,114,31,229,31,211,31,199,31,201,31,240,31,201,31,195,31,141,31,241,31,177,31,160,31,42,31,74,31,240,31,144,31,144,30,177,31,177,30,76,31,215,31,235,31,14,31,14,30,106,31,79,31,79,30,200,31,200,30,223,31,223,30,255,31,89,31,112,31,112,30,246,31,9,31,28,31,230,31,41,31,89,31,38,31,17,31,147,31,14,31,14,30,58,31,183,31,183,30,167,31,167,30,253,31,149,31,149,30,108,31,132,31,136,31,17,31,180,31,180,30,90,31,90,30,131,31,131,30,211,31,211,30,208,31,94,31,172,31,71,31,71,30,149,31,14,31,177,31,202,31,223,31,223,30,47,31,199,31,72,31,231,31,128,31,19,31,249,31,249,30,55,31,127,31,37,31,135,31,167,31,142,31,223,31,169,31,4,31,4,30,4,29,108,31,108,30,243,31,226,31,213,31,199,31,199,30,244,31,204,31,210,31,58,31,241,31,73,31,73,30,235,31,118,31,56,31,223,31,223,30,154,31,218,31,16,31,207,31,117,31,159,31,191,31,191,30,222,31,220,31,20,31,115,31,187,31,125,31,72,31,72,30,56,31,242,31,242,30,172,31,166,31,102,31,102,30,55,31,36,31,35,31,35,30,11,31,226,31,101,31,56,31,56,30,190,31,190,30,190,29,3,31,144,31,39,31,178,31,207,31,87,31,196,31,153,31,22,31,239,31,16,31,190,31,190,30,190,29,207,31,200,31,218,31,55,31,246,31,126,31,245,31,245,30,177,31,93,31,100,31,91,31,230,31,32,31,108,31,237,31,237,30,250,31,250,30,170,31,170,30,197,31,143,31,10,31,10,30,10,29,163,31,85,31,62,31,48,31,155,31,159,31,153,31,51,31,111,31,84,31,171,31,171,30,171,29,142,31,124,31,194,31,15,31,134,31,194,31,87,31,110,31,131,31,147,31,56,31,133,31,3,31,116,31,116,30,31,31,116,31,197,31,147,31,207,31,36,31,36,30,185,31,166,31,169,31,235,31,235,30,239,31,78,31,105,31,105,30,31,31,12,31,100,31,101,31,101,30,111,31,111,30,149,31,13,31,13,30,192,31,128,31,128,30,128,29,109,31,109,30,109,29,109,31,109,30,239,31,192,31,164,31,239,31,179,31,2,31,109,31,109,30,109,29,142,31,31,31,195,31,195,30,21,31,82,31,82,30,159,31,128,31,183,31,183,30,196,31,196,30,212,31,34,31,154,31,2,31,94,31,20,31,106,31,14,31,17,31,38,31,180,31,217,31,217,30,233,31,49,31,49,30,49,29,49,28,155,31,215,31,173,31,217,31,74,31,51,31,128,31,119,31,251,31,99,31,99,30,93,31,93,30,93,29,173,31,120,31,250,31,250,30,250,29,131,31,225,31,135,31,54,31,54,30,103,31,106,31,128,31,27,31,101,31,139,31,144,31,182,31,188,31,237,31,237,30,237,29,136,31,23,31,138,31,126,31,126,30,40,31,40,30,40,29,80,31,123,31,123,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
