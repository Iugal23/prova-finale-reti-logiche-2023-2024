-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_142 is
end project_tb_142;

architecture project_tb_arch_142 of project_tb_142 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 712;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (105,0,195,0,238,0,146,0,176,0,208,0,4,0,18,0,40,0,0,0,94,0,238,0,31,0,131,0,145,0,153,0,199,0,9,0,215,0,27,0,78,0,44,0,138,0,169,0,175,0,173,0,32,0,0,0,182,0,0,0,172,0,211,0,8,0,157,0,241,0,93,0,74,0,80,0,107,0,232,0,0,0,14,0,0,0,177,0,66,0,0,0,95,0,138,0,0,0,147,0,0,0,180,0,238,0,68,0,141,0,154,0,0,0,241,0,150,0,44,0,91,0,241,0,114,0,135,0,157,0,180,0,67,0,115,0,173,0,9,0,0,0,0,0,111,0,113,0,24,0,0,0,0,0,32,0,74,0,159,0,232,0,149,0,248,0,92,0,44,0,5,0,64,0,0,0,21,0,143,0,34,0,176,0,102,0,1,0,0,0,101,0,0,0,0,0,193,0,198,0,188,0,239,0,215,0,99,0,145,0,36,0,113,0,0,0,223,0,0,0,0,0,123,0,103,0,0,0,199,0,0,0,22,0,234,0,140,0,85,0,35,0,55,0,39,0,0,0,216,0,15,0,0,0,0,0,156,0,165,0,109,0,239,0,0,0,142,0,170,0,14,0,27,0,88,0,203,0,23,0,43,0,159,0,0,0,25,0,38,0,31,0,0,0,5,0,217,0,91,0,0,0,0,0,110,0,206,0,144,0,62,0,0,0,35,0,146,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,63,0,225,0,179,0,0,0,0,0,121,0,44,0,0,0,10,0,116,0,219,0,123,0,242,0,40,0,0,0,62,0,177,0,204,0,42,0,143,0,106,0,187,0,50,0,205,0,54,0,65,0,203,0,35,0,18,0,142,0,76,0,204,0,92,0,159,0,230,0,145,0,180,0,0,0,152,0,30,0,61,0,198,0,152,0,173,0,42,0,64,0,194,0,227,0,25,0,85,0,225,0,0,0,0,0,182,0,166,0,148,0,174,0,0,0,30,0,0,0,29,0,146,0,125,0,0,0,31,0,0,0,0,0,55,0,100,0,0,0,209,0,126,0,235,0,162,0,156,0,152,0,73,0,52,0,38,0,0,0,140,0,251,0,0,0,181,0,0,0,0,0,176,0,23,0,128,0,101,0,0,0,107,0,11,0,112,0,0,0,102,0,214,0,224,0,218,0,90,0,111,0,24,0,0,0,0,0,0,0,0,0,247,0,250,0,118,0,0,0,8,0,196,0,28,0,195,0,127,0,223,0,166,0,111,0,114,0,126,0,143,0,15,0,231,0,165,0,0,0,129,0,117,0,0,0,0,0,188,0,208,0,65,0,108,0,51,0,106,0,0,0,0,0,232,0,254,0,0,0,32,0,0,0,243,0,47,0,0,0,0,0,129,0,83,0,0,0,243,0,47,0,146,0,0,0,28,0,180,0,113,0,235,0,61,0,170,0,0,0,170,0,166,0,200,0,0,0,110,0,208,0,197,0,144,0,0,0,183,0,0,0,47,0,41,0,70,0,0,0,0,0,212,0,0,0,133,0,39,0,54,0,148,0,106,0,75,0,42,0,228,0,0,0,208,0,0,0,0,0,191,0,67,0,111,0,152,0,59,0,2,0,71,0,0,0,156,0,0,0,86,0,0,0,221,0,113,0,156,0,0,0,221,0,190,0,162,0,141,0,215,0,60,0,40,0,84,0,0,0,59,0,218,0,3,0,84,0,87,0,0,0,162,0,77,0,50,0,99,0,248,0,21,0,73,0,138,0,6,0,159,0,0,0,66,0,241,0,19,0,74,0,0,0,163,0,123,0,220,0,68,0,204,0,91,0,0,0,0,0,143,0,227,0,147,0,175,0,45,0,249,0,135,0,54,0,81,0,49,0,136,0,0,0,68,0,202,0,208,0,36,0,213,0,216,0,230,0,143,0,92,0,223,0,142,0,0,0,86,0,68,0,144,0,82,0,68,0,229,0,109,0,64,0,0,0,0,0,210,0,92,0,201,0,54,0,74,0,16,0,0,0,133,0,206,0,198,0,252,0,20,0,0,0,0,0,178,0,72,0,138,0,58,0,152,0,6,0,211,0,130,0,80,0,232,0,37,0,132,0,219,0,94,0,209,0,253,0,68,0,108,0,0,0,35,0,140,0,248,0,135,0,201,0,0,0,207,0,0,0,234,0,129,0,0,0,182,0,25,0,4,0,190,0,137,0,252,0,132,0,201,0,187,0,0,0,150,0,0,0,97,0,189,0,111,0,29,0,91,0,131,0,125,0,0,0,49,0,0,0,132,0,0,0,136,0,0,0,0,0,26,0,83,0,0,0,124,0,120,0,29,0,249,0,0,0,36,0,28,0,38,0,0,0,5,0,86,0,127,0,45,0,218,0,212,0,223,0,252,0,173,0,216,0,0,0,7,0,151,0,96,0,199,0,44,0,22,0,0,0,67,0,147,0,80,0,37,0,107,0,102,0,31,0,0,0,59,0,125,0,221,0,64,0,119,0,121,0,62,0,31,0,200,0,46,0,0,0,179,0,44,0,0,0,0,0,0,0,0,0,255,0,148,0,231,0,23,0,0,0,34,0,179,0,244,0,165,0,33,0,12,0,188,0,0,0,198,0,2,0,113,0,126,0,105,0,240,0,123,0,169,0,0,0,78,0,142,0,180,0,253,0,0,0,0,0,168,0,200,0,249,0,194,0,0,0,232,0,169,0,0,0,97,0,86,0,173,0,64,0,40,0,202,0,216,0,179,0,90,0,48,0,210,0,39,0,108,0,0,0,151,0,129,0,143,0,233,0,91,0,0,0,122,0,15,0,140,0,149,0,0,0,235,0,0,0,173,0,171,0,33,0,48,0,193,0,59,0,22,0,126,0,0,0,107,0,0,0,11,0,241,0,79,0,96,0,0,0,11,0,140,0,0,0,87,0,76,0,158,0,97,0,68,0,0,0,54,0,0,0,0,0,190,0,108,0,171,0,151,0,0,0,27,0,207,0,174,0,51,0,161,0,0,0,49,0,0,0,0,0,211,0,183,0,56,0,249,0,150,0,0,0,5,0,98,0,0,0,0,0,169,0,182,0,32,0,75,0,99,0,61,0,151,0,133,0,57,0,139,0,0,0,176,0,164,0,0,0,0,0,243,0,184,0,4,0,0,0,106,0,0,0,71,0,252,0,163,0,102,0);
signal scenario_full  : scenario_type := (105,31,195,31,238,31,146,31,176,31,208,31,4,31,18,31,40,31,40,30,94,31,238,31,31,31,131,31,145,31,153,31,199,31,9,31,215,31,27,31,78,31,44,31,138,31,169,31,175,31,173,31,32,31,32,30,182,31,182,30,172,31,211,31,8,31,157,31,241,31,93,31,74,31,80,31,107,31,232,31,232,30,14,31,14,30,177,31,66,31,66,30,95,31,138,31,138,30,147,31,147,30,180,31,238,31,68,31,141,31,154,31,154,30,241,31,150,31,44,31,91,31,241,31,114,31,135,31,157,31,180,31,67,31,115,31,173,31,9,31,9,30,9,29,111,31,113,31,24,31,24,30,24,29,32,31,74,31,159,31,232,31,149,31,248,31,92,31,44,31,5,31,64,31,64,30,21,31,143,31,34,31,176,31,102,31,1,31,1,30,101,31,101,30,101,29,193,31,198,31,188,31,239,31,215,31,99,31,145,31,36,31,113,31,113,30,223,31,223,30,223,29,123,31,103,31,103,30,199,31,199,30,22,31,234,31,140,31,85,31,35,31,55,31,39,31,39,30,216,31,15,31,15,30,15,29,156,31,165,31,109,31,239,31,239,30,142,31,170,31,14,31,27,31,88,31,203,31,23,31,43,31,159,31,159,30,25,31,38,31,31,31,31,30,5,31,217,31,91,31,91,30,91,29,110,31,206,31,144,31,62,31,62,30,35,31,146,31,146,30,146,29,146,28,146,27,146,26,146,25,146,24,146,23,63,31,225,31,179,31,179,30,179,29,121,31,44,31,44,30,10,31,116,31,219,31,123,31,242,31,40,31,40,30,62,31,177,31,204,31,42,31,143,31,106,31,187,31,50,31,205,31,54,31,65,31,203,31,35,31,18,31,142,31,76,31,204,31,92,31,159,31,230,31,145,31,180,31,180,30,152,31,30,31,61,31,198,31,152,31,173,31,42,31,64,31,194,31,227,31,25,31,85,31,225,31,225,30,225,29,182,31,166,31,148,31,174,31,174,30,30,31,30,30,29,31,146,31,125,31,125,30,31,31,31,30,31,29,55,31,100,31,100,30,209,31,126,31,235,31,162,31,156,31,152,31,73,31,52,31,38,31,38,30,140,31,251,31,251,30,181,31,181,30,181,29,176,31,23,31,128,31,101,31,101,30,107,31,11,31,112,31,112,30,102,31,214,31,224,31,218,31,90,31,111,31,24,31,24,30,24,29,24,28,24,27,247,31,250,31,118,31,118,30,8,31,196,31,28,31,195,31,127,31,223,31,166,31,111,31,114,31,126,31,143,31,15,31,231,31,165,31,165,30,129,31,117,31,117,30,117,29,188,31,208,31,65,31,108,31,51,31,106,31,106,30,106,29,232,31,254,31,254,30,32,31,32,30,243,31,47,31,47,30,47,29,129,31,83,31,83,30,243,31,47,31,146,31,146,30,28,31,180,31,113,31,235,31,61,31,170,31,170,30,170,31,166,31,200,31,200,30,110,31,208,31,197,31,144,31,144,30,183,31,183,30,47,31,41,31,70,31,70,30,70,29,212,31,212,30,133,31,39,31,54,31,148,31,106,31,75,31,42,31,228,31,228,30,208,31,208,30,208,29,191,31,67,31,111,31,152,31,59,31,2,31,71,31,71,30,156,31,156,30,86,31,86,30,221,31,113,31,156,31,156,30,221,31,190,31,162,31,141,31,215,31,60,31,40,31,84,31,84,30,59,31,218,31,3,31,84,31,87,31,87,30,162,31,77,31,50,31,99,31,248,31,21,31,73,31,138,31,6,31,159,31,159,30,66,31,241,31,19,31,74,31,74,30,163,31,123,31,220,31,68,31,204,31,91,31,91,30,91,29,143,31,227,31,147,31,175,31,45,31,249,31,135,31,54,31,81,31,49,31,136,31,136,30,68,31,202,31,208,31,36,31,213,31,216,31,230,31,143,31,92,31,223,31,142,31,142,30,86,31,68,31,144,31,82,31,68,31,229,31,109,31,64,31,64,30,64,29,210,31,92,31,201,31,54,31,74,31,16,31,16,30,133,31,206,31,198,31,252,31,20,31,20,30,20,29,178,31,72,31,138,31,58,31,152,31,6,31,211,31,130,31,80,31,232,31,37,31,132,31,219,31,94,31,209,31,253,31,68,31,108,31,108,30,35,31,140,31,248,31,135,31,201,31,201,30,207,31,207,30,234,31,129,31,129,30,182,31,25,31,4,31,190,31,137,31,252,31,132,31,201,31,187,31,187,30,150,31,150,30,97,31,189,31,111,31,29,31,91,31,131,31,125,31,125,30,49,31,49,30,132,31,132,30,136,31,136,30,136,29,26,31,83,31,83,30,124,31,120,31,29,31,249,31,249,30,36,31,28,31,38,31,38,30,5,31,86,31,127,31,45,31,218,31,212,31,223,31,252,31,173,31,216,31,216,30,7,31,151,31,96,31,199,31,44,31,22,31,22,30,67,31,147,31,80,31,37,31,107,31,102,31,31,31,31,30,59,31,125,31,221,31,64,31,119,31,121,31,62,31,31,31,200,31,46,31,46,30,179,31,44,31,44,30,44,29,44,28,44,27,255,31,148,31,231,31,23,31,23,30,34,31,179,31,244,31,165,31,33,31,12,31,188,31,188,30,198,31,2,31,113,31,126,31,105,31,240,31,123,31,169,31,169,30,78,31,142,31,180,31,253,31,253,30,253,29,168,31,200,31,249,31,194,31,194,30,232,31,169,31,169,30,97,31,86,31,173,31,64,31,40,31,202,31,216,31,179,31,90,31,48,31,210,31,39,31,108,31,108,30,151,31,129,31,143,31,233,31,91,31,91,30,122,31,15,31,140,31,149,31,149,30,235,31,235,30,173,31,171,31,33,31,48,31,193,31,59,31,22,31,126,31,126,30,107,31,107,30,11,31,241,31,79,31,96,31,96,30,11,31,140,31,140,30,87,31,76,31,158,31,97,31,68,31,68,30,54,31,54,30,54,29,190,31,108,31,171,31,151,31,151,30,27,31,207,31,174,31,51,31,161,31,161,30,49,31,49,30,49,29,211,31,183,31,56,31,249,31,150,31,150,30,5,31,98,31,98,30,98,29,169,31,182,31,32,31,75,31,99,31,61,31,151,31,133,31,57,31,139,31,139,30,176,31,164,31,164,30,164,29,243,31,184,31,4,31,4,30,106,31,106,30,71,31,252,31,163,31,102,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
