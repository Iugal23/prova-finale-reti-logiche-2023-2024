-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_759 is
end project_tb_759;

architecture project_tb_arch_759 of project_tb_759 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 224;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (199,0,58,0,3,0,108,0,216,0,229,0,179,0,0,0,0,0,0,0,247,0,19,0,0,0,113,0,1,0,0,0,27,0,0,0,125,0,239,0,201,0,226,0,189,0,219,0,0,0,188,0,13,0,222,0,225,0,204,0,64,0,175,0,101,0,195,0,0,0,148,0,166,0,234,0,226,0,0,0,79,0,6,0,0,0,0,0,0,0,157,0,105,0,70,0,196,0,45,0,28,0,25,0,52,0,114,0,143,0,46,0,0,0,0,0,212,0,76,0,14,0,37,0,0,0,34,0,88,0,0,0,0,0,166,0,0,0,144,0,22,0,0,0,84,0,147,0,0,0,58,0,201,0,158,0,82,0,18,0,55,0,182,0,121,0,167,0,64,0,254,0,46,0,164,0,184,0,234,0,27,0,185,0,0,0,207,0,116,0,0,0,23,0,150,0,204,0,0,0,115,0,224,0,0,0,193,0,120,0,0,0,86,0,0,0,101,0,203,0,0,0,66,0,0,0,101,0,214,0,222,0,198,0,30,0,107,0,125,0,90,0,130,0,29,0,22,0,17,0,254,0,0,0,219,0,216,0,196,0,127,0,97,0,0,0,248,0,197,0,250,0,113,0,41,0,0,0,159,0,0,0,186,0,107,0,0,0,134,0,170,0,63,0,254,0,149,0,0,0,140,0,71,0,74,0,36,0,62,0,110,0,190,0,253,0,210,0,76,0,196,0,140,0,200,0,53,0,61,0,68,0,152,0,0,0,0,0,113,0,112,0,176,0,160,0,91,0,214,0,121,0,126,0,143,0,130,0,43,0,106,0,0,0,24,0,0,0,106,0,117,0,156,0,0,0,230,0,53,0,0,0,9,0,42,0,0,0,0,0,151,0,195,0,0,0,0,0,230,0,0,0,24,0,252,0,126,0,152,0,205,0,189,0,181,0,225,0,111,0,164,0,0,0,207,0,207,0,13,0,162,0,0,0,208,0,0,0,0,0,181,0,110,0,192,0,27,0);
signal scenario_full  : scenario_type := (199,31,58,31,3,31,108,31,216,31,229,31,179,31,179,30,179,29,179,28,247,31,19,31,19,30,113,31,1,31,1,30,27,31,27,30,125,31,239,31,201,31,226,31,189,31,219,31,219,30,188,31,13,31,222,31,225,31,204,31,64,31,175,31,101,31,195,31,195,30,148,31,166,31,234,31,226,31,226,30,79,31,6,31,6,30,6,29,6,28,157,31,105,31,70,31,196,31,45,31,28,31,25,31,52,31,114,31,143,31,46,31,46,30,46,29,212,31,76,31,14,31,37,31,37,30,34,31,88,31,88,30,88,29,166,31,166,30,144,31,22,31,22,30,84,31,147,31,147,30,58,31,201,31,158,31,82,31,18,31,55,31,182,31,121,31,167,31,64,31,254,31,46,31,164,31,184,31,234,31,27,31,185,31,185,30,207,31,116,31,116,30,23,31,150,31,204,31,204,30,115,31,224,31,224,30,193,31,120,31,120,30,86,31,86,30,101,31,203,31,203,30,66,31,66,30,101,31,214,31,222,31,198,31,30,31,107,31,125,31,90,31,130,31,29,31,22,31,17,31,254,31,254,30,219,31,216,31,196,31,127,31,97,31,97,30,248,31,197,31,250,31,113,31,41,31,41,30,159,31,159,30,186,31,107,31,107,30,134,31,170,31,63,31,254,31,149,31,149,30,140,31,71,31,74,31,36,31,62,31,110,31,190,31,253,31,210,31,76,31,196,31,140,31,200,31,53,31,61,31,68,31,152,31,152,30,152,29,113,31,112,31,176,31,160,31,91,31,214,31,121,31,126,31,143,31,130,31,43,31,106,31,106,30,24,31,24,30,106,31,117,31,156,31,156,30,230,31,53,31,53,30,9,31,42,31,42,30,42,29,151,31,195,31,195,30,195,29,230,31,230,30,24,31,252,31,126,31,152,31,205,31,189,31,181,31,225,31,111,31,164,31,164,30,207,31,207,31,13,31,162,31,162,30,208,31,208,30,208,29,181,31,110,31,192,31,27,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
