-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 155;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (191,0,204,0,50,0,0,0,0,0,54,0,154,0,47,0,28,0,163,0,0,0,214,0,241,0,152,0,0,0,2,0,4,0,217,0,148,0,173,0,111,0,132,0,0,0,244,0,115,0,250,0,73,0,227,0,233,0,199,0,242,0,183,0,167,0,0,0,129,0,0,0,198,0,194,0,180,0,190,0,1,0,0,0,10,0,125,0,0,0,155,0,88,0,0,0,0,0,2,0,85,0,0,0,236,0,189,0,117,0,161,0,229,0,0,0,0,0,178,0,0,0,55,0,170,0,254,0,56,0,181,0,72,0,37,0,84,0,0,0,103,0,206,0,201,0,114,0,22,0,139,0,30,0,206,0,0,0,0,0,220,0,31,0,141,0,110,0,0,0,126,0,13,0,0,0,0,0,0,0,0,0,99,0,189,0,0,0,221,0,1,0,111,0,45,0,244,0,0,0,184,0,0,0,240,0,163,0,248,0,77,0,169,0,197,0,205,0,111,0,246,0,85,0,151,0,202,0,227,0,99,0,89,0,53,0,49,0,92,0,125,0,151,0,50,0,0,0,189,0,194,0,174,0,0,0,64,0,214,0,190,0,0,0,0,0,201,0,174,0,147,0,6,0,15,0,172,0,138,0,200,0,253,0,222,0,66,0,182,0,146,0,117,0,255,0,0,0,0,0,161,0,59,0,205,0,177,0,0,0);
signal scenario_full  : scenario_type := (191,31,204,31,50,31,50,30,50,29,54,31,154,31,47,31,28,31,163,31,163,30,214,31,241,31,152,31,152,30,2,31,4,31,217,31,148,31,173,31,111,31,132,31,132,30,244,31,115,31,250,31,73,31,227,31,233,31,199,31,242,31,183,31,167,31,167,30,129,31,129,30,198,31,194,31,180,31,190,31,1,31,1,30,10,31,125,31,125,30,155,31,88,31,88,30,88,29,2,31,85,31,85,30,236,31,189,31,117,31,161,31,229,31,229,30,229,29,178,31,178,30,55,31,170,31,254,31,56,31,181,31,72,31,37,31,84,31,84,30,103,31,206,31,201,31,114,31,22,31,139,31,30,31,206,31,206,30,206,29,220,31,31,31,141,31,110,31,110,30,126,31,13,31,13,30,13,29,13,28,13,27,99,31,189,31,189,30,221,31,1,31,111,31,45,31,244,31,244,30,184,31,184,30,240,31,163,31,248,31,77,31,169,31,197,31,205,31,111,31,246,31,85,31,151,31,202,31,227,31,99,31,89,31,53,31,49,31,92,31,125,31,151,31,50,31,50,30,189,31,194,31,174,31,174,30,64,31,214,31,190,31,190,30,190,29,201,31,174,31,147,31,6,31,15,31,172,31,138,31,200,31,253,31,222,31,66,31,182,31,146,31,117,31,255,31,255,30,255,29,161,31,59,31,205,31,177,31,177,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
