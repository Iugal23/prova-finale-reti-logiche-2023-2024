-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 815;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (123,0,83,0,37,0,52,0,0,0,0,0,158,0,149,0,41,0,223,0,185,0,223,0,120,0,67,0,78,0,97,0,166,0,28,0,13,0,125,0,92,0,44,0,0,0,18,0,23,0,0,0,118,0,202,0,55,0,181,0,69,0,250,0,57,0,239,0,237,0,17,0,92,0,185,0,175,0,144,0,177,0,96,0,210,0,9,0,140,0,176,0,19,0,137,0,72,0,206,0,0,0,240,0,162,0,147,0,111,0,246,0,252,0,59,0,0,0,136,0,208,0,73,0,24,0,201,0,127,0,103,0,8,0,190,0,73,0,74,0,221,0,98,0,57,0,10,0,74,0,28,0,127,0,164,0,0,0,85,0,28,0,34,0,7,0,186,0,169,0,189,0,245,0,0,0,39,0,149,0,52,0,193,0,188,0,98,0,0,0,148,0,25,0,231,0,250,0,156,0,27,0,0,0,57,0,201,0,252,0,0,0,151,0,0,0,126,0,0,0,242,0,81,0,249,0,229,0,117,0,0,0,109,0,88,0,101,0,42,0,195,0,0,0,0,0,152,0,158,0,245,0,58,0,11,0,157,0,65,0,53,0,11,0,71,0,39,0,103,0,130,0,73,0,134,0,121,0,60,0,0,0,0,0,210,0,0,0,18,0,2,0,0,0,139,0,165,0,198,0,235,0,0,0,61,0,0,0,132,0,93,0,0,0,15,0,69,0,4,0,18,0,182,0,190,0,224,0,2,0,131,0,161,0,142,0,187,0,209,0,135,0,0,0,218,0,0,0,129,0,0,0,41,0,0,0,128,0,141,0,121,0,49,0,237,0,0,0,105,0,122,0,0,0,156,0,92,0,108,0,58,0,196,0,0,0,0,0,0,0,43,0,46,0,103,0,83,0,206,0,209,0,162,0,0,0,0,0,0,0,204,0,0,0,13,0,72,0,119,0,190,0,243,0,37,0,149,0,0,0,22,0,59,0,137,0,181,0,132,0,147,0,185,0,0,0,143,0,75,0,90,0,42,0,0,0,225,0,0,0,73,0,0,0,126,0,208,0,65,0,66,0,36,0,0,0,239,0,0,0,72,0,64,0,135,0,178,0,0,0,0,0,68,0,110,0,135,0,0,0,0,0,164,0,160,0,187,0,55,0,187,0,0,0,81,0,129,0,0,0,70,0,0,0,66,0,42,0,187,0,0,0,237,0,229,0,0,0,106,0,127,0,38,0,241,0,0,0,239,0,0,0,110,0,9,0,196,0,128,0,43,0,150,0,0,0,194,0,209,0,0,0,165,0,108,0,200,0,74,0,91,0,246,0,0,0,28,0,193,0,60,0,46,0,27,0,32,0,25,0,182,0,103,0,220,0,78,0,155,0,58,0,154,0,173,0,133,0,0,0,207,0,221,0,252,0,0,0,160,0,119,0,221,0,0,0,0,0,0,0,189,0,233,0,6,0,246,0,54,0,251,0,96,0,85,0,0,0,101,0,0,0,179,0,0,0,232,0,184,0,227,0,137,0,142,0,76,0,213,0,26,0,212,0,173,0,126,0,70,0,114,0,0,0,140,0,140,0,246,0,25,0,10,0,205,0,0,0,35,0,179,0,159,0,53,0,0,0,89,0,172,0,171,0,160,0,59,0,98,0,254,0,86,0,0,0,0,0,70,0,0,0,163,0,44,0,105,0,27,0,34,0,180,0,139,0,126,0,58,0,98,0,99,0,0,0,59,0,102,0,228,0,0,0,236,0,67,0,0,0,3,0,43,0,158,0,48,0,0,0,93,0,0,0,179,0,240,0,13,0,60,0,178,0,0,0,40,0,43,0,92,0,230,0,63,0,56,0,101,0,50,0,133,0,89,0,85,0,86,0,0,0,252,0,239,0,66,0,0,0,0,0,107,0,198,0,44,0,0,0,140,0,208,0,202,0,233,0,169,0,22,0,89,0,0,0,45,0,221,0,198,0,176,0,46,0,14,0,61,0,182,0,0,0,0,0,140,0,0,0,196,0,237,0,0,0,81,0,57,0,239,0,6,0,227,0,183,0,11,0,149,0,0,0,181,0,193,0,249,0,145,0,142,0,80,0,41,0,147,0,231,0,124,0,0,0,233,0,0,0,0,0,0,0,151,0,188,0,49,0,45,0,164,0,227,0,0,0,27,0,12,0,58,0,0,0,224,0,174,0,60,0,110,0,95,0,79,0,176,0,160,0,129,0,111,0,231,0,101,0,39,0,84,0,182,0,20,0,229,0,0,0,120,0,219,0,0,0,0,0,13,0,208,0,207,0,210,0,59,0,211,0,224,0,0,0,222,0,86,0,218,0,37,0,191,0,0,0,215,0,171,0,241,0,132,0,178,0,30,0,35,0,210,0,173,0,238,0,93,0,211,0,179,0,229,0,83,0,55,0,0,0,245,0,124,0,220,0,171,0,247,0,0,0,57,0,212,0,204,0,188,0,175,0,171,0,0,0,34,0,22,0,238,0,142,0,81,0,203,0,71,0,181,0,102,0,0,0,196,0,217,0,156,0,202,0,110,0,0,0,241,0,0,0,64,0,0,0,62,0,31,0,0,0,53,0,171,0,53,0,199,0,237,0,19,0,250,0,206,0,0,0,0,0,234,0,219,0,63,0,158,0,68,0,129,0,16,0,0,0,179,0,231,0,133,0,137,0,0,0,0,0,0,0,13,0,62,0,35,0,230,0,231,0,81,0,169,0,160,0,44,0,166,0,145,0,13,0,179,0,132,0,170,0,184,0,180,0,72,0,112,0,216,0,138,0,26,0,131,0,0,0,33,0,185,0,0,0,226,0,127,0,118,0,121,0,213,0,224,0,248,0,214,0,54,0,119,0,0,0,58,0,0,0,61,0,130,0,130,0,161,0,231,0,137,0,177,0,84,0,191,0,140,0,0,0,203,0,220,0,38,0,176,0,38,0,71,0,64,0,113,0,38,0,117,0,242,0,31,0,118,0,0,0,52,0,0,0,5,0,38,0,57,0,74,0,40,0,78,0,138,0,55,0,0,0,47,0,0,0,235,0,0,0,0,0,178,0,8,0,207,0,253,0,130,0,56,0,146,0,108,0,194,0,46,0,44,0,172,0,0,0,21,0,7,0,175,0,0,0,0,0,177,0,191,0,239,0,172,0,101,0,60,0,111,0,243,0,51,0,96,0,87,0,85,0,153,0,152,0,143,0,125,0,223,0,188,0,201,0,242,0,89,0,0,0,102,0,0,0,117,0,126,0,37,0,24,0,39,0,0,0,0,0,238,0,23,0,5,0,81,0,204,0,171,0,0,0,145,0,32,0,151,0,199,0,207,0,126,0,93,0,0,0,0,0,198,0,232,0,0,0,105,0,0,0,164,0,31,0,241,0,173,0,117,0,75,0,205,0,29,0,237,0,95,0,0,0,145,0,0,0,251,0,92,0,0,0,237,0,44,0,231,0,48,0,242,0,0,0,135,0,87,0,92,0,35,0,45,0,55,0,36,0,0,0,132,0,59,0,111,0,199,0,5,0,0,0,147,0,233,0,76,0,4,0,151,0,122,0,196,0,190,0,0,0,120,0,153,0,0,0,112,0,0,0,145,0,215,0,38,0,253,0,73,0,143,0,79,0,16,0,204,0,11,0,220,0,180,0,25,0,60,0,87,0,59,0,0,0);
signal scenario_full  : scenario_type := (123,31,83,31,37,31,52,31,52,30,52,29,158,31,149,31,41,31,223,31,185,31,223,31,120,31,67,31,78,31,97,31,166,31,28,31,13,31,125,31,92,31,44,31,44,30,18,31,23,31,23,30,118,31,202,31,55,31,181,31,69,31,250,31,57,31,239,31,237,31,17,31,92,31,185,31,175,31,144,31,177,31,96,31,210,31,9,31,140,31,176,31,19,31,137,31,72,31,206,31,206,30,240,31,162,31,147,31,111,31,246,31,252,31,59,31,59,30,136,31,208,31,73,31,24,31,201,31,127,31,103,31,8,31,190,31,73,31,74,31,221,31,98,31,57,31,10,31,74,31,28,31,127,31,164,31,164,30,85,31,28,31,34,31,7,31,186,31,169,31,189,31,245,31,245,30,39,31,149,31,52,31,193,31,188,31,98,31,98,30,148,31,25,31,231,31,250,31,156,31,27,31,27,30,57,31,201,31,252,31,252,30,151,31,151,30,126,31,126,30,242,31,81,31,249,31,229,31,117,31,117,30,109,31,88,31,101,31,42,31,195,31,195,30,195,29,152,31,158,31,245,31,58,31,11,31,157,31,65,31,53,31,11,31,71,31,39,31,103,31,130,31,73,31,134,31,121,31,60,31,60,30,60,29,210,31,210,30,18,31,2,31,2,30,139,31,165,31,198,31,235,31,235,30,61,31,61,30,132,31,93,31,93,30,15,31,69,31,4,31,18,31,182,31,190,31,224,31,2,31,131,31,161,31,142,31,187,31,209,31,135,31,135,30,218,31,218,30,129,31,129,30,41,31,41,30,128,31,141,31,121,31,49,31,237,31,237,30,105,31,122,31,122,30,156,31,92,31,108,31,58,31,196,31,196,30,196,29,196,28,43,31,46,31,103,31,83,31,206,31,209,31,162,31,162,30,162,29,162,28,204,31,204,30,13,31,72,31,119,31,190,31,243,31,37,31,149,31,149,30,22,31,59,31,137,31,181,31,132,31,147,31,185,31,185,30,143,31,75,31,90,31,42,31,42,30,225,31,225,30,73,31,73,30,126,31,208,31,65,31,66,31,36,31,36,30,239,31,239,30,72,31,64,31,135,31,178,31,178,30,178,29,68,31,110,31,135,31,135,30,135,29,164,31,160,31,187,31,55,31,187,31,187,30,81,31,129,31,129,30,70,31,70,30,66,31,42,31,187,31,187,30,237,31,229,31,229,30,106,31,127,31,38,31,241,31,241,30,239,31,239,30,110,31,9,31,196,31,128,31,43,31,150,31,150,30,194,31,209,31,209,30,165,31,108,31,200,31,74,31,91,31,246,31,246,30,28,31,193,31,60,31,46,31,27,31,32,31,25,31,182,31,103,31,220,31,78,31,155,31,58,31,154,31,173,31,133,31,133,30,207,31,221,31,252,31,252,30,160,31,119,31,221,31,221,30,221,29,221,28,189,31,233,31,6,31,246,31,54,31,251,31,96,31,85,31,85,30,101,31,101,30,179,31,179,30,232,31,184,31,227,31,137,31,142,31,76,31,213,31,26,31,212,31,173,31,126,31,70,31,114,31,114,30,140,31,140,31,246,31,25,31,10,31,205,31,205,30,35,31,179,31,159,31,53,31,53,30,89,31,172,31,171,31,160,31,59,31,98,31,254,31,86,31,86,30,86,29,70,31,70,30,163,31,44,31,105,31,27,31,34,31,180,31,139,31,126,31,58,31,98,31,99,31,99,30,59,31,102,31,228,31,228,30,236,31,67,31,67,30,3,31,43,31,158,31,48,31,48,30,93,31,93,30,179,31,240,31,13,31,60,31,178,31,178,30,40,31,43,31,92,31,230,31,63,31,56,31,101,31,50,31,133,31,89,31,85,31,86,31,86,30,252,31,239,31,66,31,66,30,66,29,107,31,198,31,44,31,44,30,140,31,208,31,202,31,233,31,169,31,22,31,89,31,89,30,45,31,221,31,198,31,176,31,46,31,14,31,61,31,182,31,182,30,182,29,140,31,140,30,196,31,237,31,237,30,81,31,57,31,239,31,6,31,227,31,183,31,11,31,149,31,149,30,181,31,193,31,249,31,145,31,142,31,80,31,41,31,147,31,231,31,124,31,124,30,233,31,233,30,233,29,233,28,151,31,188,31,49,31,45,31,164,31,227,31,227,30,27,31,12,31,58,31,58,30,224,31,174,31,60,31,110,31,95,31,79,31,176,31,160,31,129,31,111,31,231,31,101,31,39,31,84,31,182,31,20,31,229,31,229,30,120,31,219,31,219,30,219,29,13,31,208,31,207,31,210,31,59,31,211,31,224,31,224,30,222,31,86,31,218,31,37,31,191,31,191,30,215,31,171,31,241,31,132,31,178,31,30,31,35,31,210,31,173,31,238,31,93,31,211,31,179,31,229,31,83,31,55,31,55,30,245,31,124,31,220,31,171,31,247,31,247,30,57,31,212,31,204,31,188,31,175,31,171,31,171,30,34,31,22,31,238,31,142,31,81,31,203,31,71,31,181,31,102,31,102,30,196,31,217,31,156,31,202,31,110,31,110,30,241,31,241,30,64,31,64,30,62,31,31,31,31,30,53,31,171,31,53,31,199,31,237,31,19,31,250,31,206,31,206,30,206,29,234,31,219,31,63,31,158,31,68,31,129,31,16,31,16,30,179,31,231,31,133,31,137,31,137,30,137,29,137,28,13,31,62,31,35,31,230,31,231,31,81,31,169,31,160,31,44,31,166,31,145,31,13,31,179,31,132,31,170,31,184,31,180,31,72,31,112,31,216,31,138,31,26,31,131,31,131,30,33,31,185,31,185,30,226,31,127,31,118,31,121,31,213,31,224,31,248,31,214,31,54,31,119,31,119,30,58,31,58,30,61,31,130,31,130,31,161,31,231,31,137,31,177,31,84,31,191,31,140,31,140,30,203,31,220,31,38,31,176,31,38,31,71,31,64,31,113,31,38,31,117,31,242,31,31,31,118,31,118,30,52,31,52,30,5,31,38,31,57,31,74,31,40,31,78,31,138,31,55,31,55,30,47,31,47,30,235,31,235,30,235,29,178,31,8,31,207,31,253,31,130,31,56,31,146,31,108,31,194,31,46,31,44,31,172,31,172,30,21,31,7,31,175,31,175,30,175,29,177,31,191,31,239,31,172,31,101,31,60,31,111,31,243,31,51,31,96,31,87,31,85,31,153,31,152,31,143,31,125,31,223,31,188,31,201,31,242,31,89,31,89,30,102,31,102,30,117,31,126,31,37,31,24,31,39,31,39,30,39,29,238,31,23,31,5,31,81,31,204,31,171,31,171,30,145,31,32,31,151,31,199,31,207,31,126,31,93,31,93,30,93,29,198,31,232,31,232,30,105,31,105,30,164,31,31,31,241,31,173,31,117,31,75,31,205,31,29,31,237,31,95,31,95,30,145,31,145,30,251,31,92,31,92,30,237,31,44,31,231,31,48,31,242,31,242,30,135,31,87,31,92,31,35,31,45,31,55,31,36,31,36,30,132,31,59,31,111,31,199,31,5,31,5,30,147,31,233,31,76,31,4,31,151,31,122,31,196,31,190,31,190,30,120,31,153,31,153,30,112,31,112,30,145,31,215,31,38,31,253,31,73,31,143,31,79,31,16,31,204,31,11,31,220,31,180,31,25,31,60,31,87,31,59,31,59,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
