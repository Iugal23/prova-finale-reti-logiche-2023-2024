-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_733 is
end project_tb_733;

architecture project_tb_arch_733 of project_tb_733 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 424;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,235,0,252,0,13,0,95,0,0,0,0,0,254,0,211,0,5,0,196,0,34,0,224,0,0,0,137,0,0,0,247,0,0,0,231,0,114,0,246,0,10,0,74,0,69,0,164,0,104,0,86,0,0,0,0,0,70,0,119,0,168,0,26,0,175,0,64,0,239,0,239,0,205,0,0,0,176,0,167,0,82,0,84,0,0,0,229,0,180,0,0,0,219,0,161,0,53,0,240,0,250,0,41,0,224,0,157,0,0,0,192,0,120,0,78,0,135,0,7,0,0,0,106,0,53,0,179,0,0,0,198,0,116,0,94,0,95,0,244,0,143,0,242,0,192,0,214,0,186,0,196,0,95,0,75,0,206,0,20,0,164,0,62,0,140,0,9,0,33,0,131,0,220,0,132,0,0,0,56,0,0,0,40,0,44,0,202,0,0,0,137,0,60,0,173,0,210,0,6,0,0,0,120,0,147,0,0,0,79,0,20,0,30,0,139,0,210,0,22,0,46,0,110,0,0,0,188,0,5,0,125,0,0,0,182,0,18,0,148,0,0,0,117,0,223,0,204,0,118,0,161,0,0,0,195,0,4,0,36,0,101,0,0,0,167,0,0,0,112,0,159,0,119,0,253,0,74,0,12,0,205,0,0,0,183,0,6,0,0,0,0,0,114,0,205,0,0,0,78,0,0,0,216,0,31,0,205,0,0,0,11,0,215,0,203,0,130,0,45,0,238,0,152,0,63,0,161,0,221,0,0,0,55,0,119,0,0,0,241,0,88,0,0,0,47,0,210,0,178,0,255,0,189,0,0,0,250,0,159,0,97,0,0,0,76,0,202,0,238,0,56,0,45,0,60,0,118,0,139,0,0,0,56,0,41,0,144,0,214,0,139,0,50,0,163,0,189,0,152,0,5,0,123,0,0,0,0,0,136,0,62,0,1,0,129,0,132,0,69,0,234,0,156,0,12,0,62,0,12,0,46,0,0,0,212,0,176,0,10,0,71,0,97,0,36,0,241,0,222,0,118,0,245,0,46,0,236,0,0,0,2,0,161,0,86,0,144,0,77,0,78,0,132,0,196,0,255,0,150,0,185,0,247,0,76,0,166,0,9,0,30,0,0,0,30,0,230,0,0,0,54,0,143,0,100,0,252,0,23,0,6,0,248,0,42,0,42,0,32,0,208,0,222,0,64,0,174,0,36,0,235,0,90,0,102,0,145,0,211,0,192,0,73,0,230,0,195,0,4,0,190,0,225,0,0,0,162,0,222,0,4,0,222,0,169,0,0,0,213,0,203,0,0,0,51,0,49,0,0,0,141,0,0,0,195,0,85,0,125,0,0,0,70,0,134,0,189,0,132,0,71,0,15,0,223,0,0,0,33,0,35,0,174,0,247,0,0,0,0,0,70,0,182,0,75,0,255,0,132,0,176,0,251,0,124,0,0,0,203,0,146,0,224,0,178,0,56,0,0,0,64,0,153,0,234,0,190,0,0,0,149,0,0,0,0,0,143,0,177,0,9,0,0,0,213,0,133,0,227,0,0,0,0,0,230,0,49,0,32,0,76,0,23,0,195,0,234,0,175,0,253,0,122,0,102,0,175,0,193,0,136,0,242,0,230,0,110,0,222,0,72,0,0,0,0,0,146,0,177,0,0,0,50,0,196,0,174,0,0,0,85,0,47,0,188,0,55,0,111,0,94,0,29,0,2,0,0,0,161,0,220,0,121,0,8,0,58,0,239,0,135,0,74,0,115,0,230,0,0,0,0,0,233,0,0,0,0,0,236,0,0,0,24,0,188,0,37,0,221,0,148,0,179,0,192,0,126,0,212,0,0,0,251,0,166,0,4,0,122,0,161,0,169,0,0,0,187,0,42,0,83,0,128,0,235,0,57,0,111,0,229,0,125,0,0,0);
signal scenario_full  : scenario_type := (0,0,235,31,252,31,13,31,95,31,95,30,95,29,254,31,211,31,5,31,196,31,34,31,224,31,224,30,137,31,137,30,247,31,247,30,231,31,114,31,246,31,10,31,74,31,69,31,164,31,104,31,86,31,86,30,86,29,70,31,119,31,168,31,26,31,175,31,64,31,239,31,239,31,205,31,205,30,176,31,167,31,82,31,84,31,84,30,229,31,180,31,180,30,219,31,161,31,53,31,240,31,250,31,41,31,224,31,157,31,157,30,192,31,120,31,78,31,135,31,7,31,7,30,106,31,53,31,179,31,179,30,198,31,116,31,94,31,95,31,244,31,143,31,242,31,192,31,214,31,186,31,196,31,95,31,75,31,206,31,20,31,164,31,62,31,140,31,9,31,33,31,131,31,220,31,132,31,132,30,56,31,56,30,40,31,44,31,202,31,202,30,137,31,60,31,173,31,210,31,6,31,6,30,120,31,147,31,147,30,79,31,20,31,30,31,139,31,210,31,22,31,46,31,110,31,110,30,188,31,5,31,125,31,125,30,182,31,18,31,148,31,148,30,117,31,223,31,204,31,118,31,161,31,161,30,195,31,4,31,36,31,101,31,101,30,167,31,167,30,112,31,159,31,119,31,253,31,74,31,12,31,205,31,205,30,183,31,6,31,6,30,6,29,114,31,205,31,205,30,78,31,78,30,216,31,31,31,205,31,205,30,11,31,215,31,203,31,130,31,45,31,238,31,152,31,63,31,161,31,221,31,221,30,55,31,119,31,119,30,241,31,88,31,88,30,47,31,210,31,178,31,255,31,189,31,189,30,250,31,159,31,97,31,97,30,76,31,202,31,238,31,56,31,45,31,60,31,118,31,139,31,139,30,56,31,41,31,144,31,214,31,139,31,50,31,163,31,189,31,152,31,5,31,123,31,123,30,123,29,136,31,62,31,1,31,129,31,132,31,69,31,234,31,156,31,12,31,62,31,12,31,46,31,46,30,212,31,176,31,10,31,71,31,97,31,36,31,241,31,222,31,118,31,245,31,46,31,236,31,236,30,2,31,161,31,86,31,144,31,77,31,78,31,132,31,196,31,255,31,150,31,185,31,247,31,76,31,166,31,9,31,30,31,30,30,30,31,230,31,230,30,54,31,143,31,100,31,252,31,23,31,6,31,248,31,42,31,42,31,32,31,208,31,222,31,64,31,174,31,36,31,235,31,90,31,102,31,145,31,211,31,192,31,73,31,230,31,195,31,4,31,190,31,225,31,225,30,162,31,222,31,4,31,222,31,169,31,169,30,213,31,203,31,203,30,51,31,49,31,49,30,141,31,141,30,195,31,85,31,125,31,125,30,70,31,134,31,189,31,132,31,71,31,15,31,223,31,223,30,33,31,35,31,174,31,247,31,247,30,247,29,70,31,182,31,75,31,255,31,132,31,176,31,251,31,124,31,124,30,203,31,146,31,224,31,178,31,56,31,56,30,64,31,153,31,234,31,190,31,190,30,149,31,149,30,149,29,143,31,177,31,9,31,9,30,213,31,133,31,227,31,227,30,227,29,230,31,49,31,32,31,76,31,23,31,195,31,234,31,175,31,253,31,122,31,102,31,175,31,193,31,136,31,242,31,230,31,110,31,222,31,72,31,72,30,72,29,146,31,177,31,177,30,50,31,196,31,174,31,174,30,85,31,47,31,188,31,55,31,111,31,94,31,29,31,2,31,2,30,161,31,220,31,121,31,8,31,58,31,239,31,135,31,74,31,115,31,230,31,230,30,230,29,233,31,233,30,233,29,236,31,236,30,24,31,188,31,37,31,221,31,148,31,179,31,192,31,126,31,212,31,212,30,251,31,166,31,4,31,122,31,161,31,169,31,169,30,187,31,42,31,83,31,128,31,235,31,57,31,111,31,229,31,125,31,125,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
