-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 248;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,96,0,228,0,243,0,21,0,154,0,132,0,79,0,17,0,36,0,0,0,34,0,168,0,2,0,0,0,49,0,10,0,107,0,163,0,243,0,171,0,72,0,244,0,76,0,121,0,118,0,183,0,115,0,162,0,168,0,51,0,0,0,21,0,80,0,0,0,240,0,45,0,0,0,8,0,4,0,113,0,145,0,0,0,143,0,159,0,240,0,231,0,77,0,0,0,62,0,3,0,0,0,206,0,22,0,203,0,68,0,54,0,91,0,0,0,142,0,0,0,0,0,0,0,217,0,131,0,251,0,27,0,0,0,92,0,157,0,5,0,0,0,180,0,112,0,243,0,0,0,205,0,199,0,188,0,156,0,130,0,109,0,132,0,0,0,215,0,169,0,145,0,131,0,0,0,145,0,182,0,0,0,121,0,150,0,97,0,229,0,228,0,220,0,196,0,74,0,168,0,100,0,209,0,72,0,67,0,32,0,170,0,36,0,0,0,231,0,0,0,44,0,0,0,0,0,14,0,8,0,56,0,177,0,241,0,0,0,5,0,113,0,228,0,212,0,0,0,59,0,72,0,200,0,85,0,99,0,0,0,229,0,0,0,0,0,0,0,138,0,0,0,227,0,0,0,98,0,9,0,104,0,0,0,167,0,253,0,237,0,123,0,0,0,46,0,0,0,94,0,74,0,50,0,185,0,146,0,129,0,6,0,244,0,0,0,0,0,120,0,33,0,0,0,5,0,0,0,0,0,198,0,73,0,249,0,212,0,103,0,91,0,236,0,185,0,136,0,65,0,134,0,196,0,195,0,224,0,38,0,201,0,0,0,42,0,150,0,69,0,114,0,75,0,108,0,108,0,6,0,35,0,154,0,0,0,225,0,218,0,80,0,0,0,68,0,210,0,123,0,196,0,52,0,144,0,0,0,163,0,37,0,218,0,254,0,0,0,0,0,0,0,133,0,214,0,243,0,29,0,0,0,159,0,0,0,139,0,101,0,0,0,0,0,0,0,111,0,221,0,238,0,0,0,0,0,253,0,254,0,0,0,171,0,207,0,113,0,33,0,221,0,153,0,99,0,135,0,91,0,0,0,57,0,17,0,145,0,231,0,151,0);
signal scenario_full  : scenario_type := (0,0,0,0,96,31,228,31,243,31,21,31,154,31,132,31,79,31,17,31,36,31,36,30,34,31,168,31,2,31,2,30,49,31,10,31,107,31,163,31,243,31,171,31,72,31,244,31,76,31,121,31,118,31,183,31,115,31,162,31,168,31,51,31,51,30,21,31,80,31,80,30,240,31,45,31,45,30,8,31,4,31,113,31,145,31,145,30,143,31,159,31,240,31,231,31,77,31,77,30,62,31,3,31,3,30,206,31,22,31,203,31,68,31,54,31,91,31,91,30,142,31,142,30,142,29,142,28,217,31,131,31,251,31,27,31,27,30,92,31,157,31,5,31,5,30,180,31,112,31,243,31,243,30,205,31,199,31,188,31,156,31,130,31,109,31,132,31,132,30,215,31,169,31,145,31,131,31,131,30,145,31,182,31,182,30,121,31,150,31,97,31,229,31,228,31,220,31,196,31,74,31,168,31,100,31,209,31,72,31,67,31,32,31,170,31,36,31,36,30,231,31,231,30,44,31,44,30,44,29,14,31,8,31,56,31,177,31,241,31,241,30,5,31,113,31,228,31,212,31,212,30,59,31,72,31,200,31,85,31,99,31,99,30,229,31,229,30,229,29,229,28,138,31,138,30,227,31,227,30,98,31,9,31,104,31,104,30,167,31,253,31,237,31,123,31,123,30,46,31,46,30,94,31,74,31,50,31,185,31,146,31,129,31,6,31,244,31,244,30,244,29,120,31,33,31,33,30,5,31,5,30,5,29,198,31,73,31,249,31,212,31,103,31,91,31,236,31,185,31,136,31,65,31,134,31,196,31,195,31,224,31,38,31,201,31,201,30,42,31,150,31,69,31,114,31,75,31,108,31,108,31,6,31,35,31,154,31,154,30,225,31,218,31,80,31,80,30,68,31,210,31,123,31,196,31,52,31,144,31,144,30,163,31,37,31,218,31,254,31,254,30,254,29,254,28,133,31,214,31,243,31,29,31,29,30,159,31,159,30,139,31,101,31,101,30,101,29,101,28,111,31,221,31,238,31,238,30,238,29,253,31,254,31,254,30,171,31,207,31,113,31,33,31,221,31,153,31,99,31,135,31,91,31,91,30,57,31,17,31,145,31,231,31,151,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
