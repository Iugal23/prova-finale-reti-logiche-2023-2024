-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_870 is
end project_tb_870;

architecture project_tb_arch_870 of project_tb_870 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 340;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,159,0,12,0,0,0,87,0,43,0,106,0,50,0,0,0,101,0,178,0,0,0,0,0,144,0,149,0,221,0,0,0,187,0,87,0,191,0,218,0,157,0,159,0,11,0,224,0,127,0,248,0,199,0,14,0,196,0,159,0,148,0,156,0,172,0,63,0,234,0,182,0,245,0,0,0,104,0,130,0,143,0,0,0,0,0,168,0,47,0,0,0,0,0,196,0,41,0,0,0,206,0,142,0,0,0,0,0,47,0,45,0,50,0,94,0,0,0,255,0,179,0,116,0,227,0,195,0,169,0,60,0,234,0,253,0,0,0,143,0,243,0,129,0,197,0,4,0,9,0,250,0,196,0,60,0,0,0,204,0,13,0,128,0,0,0,208,0,33,0,181,0,0,0,0,0,87,0,73,0,234,0,0,0,0,0,137,0,227,0,204,0,255,0,32,0,0,0,0,0,61,0,65,0,4,0,231,0,67,0,40,0,79,0,93,0,245,0,143,0,105,0,0,0,135,0,248,0,0,0,183,0,0,0,47,0,236,0,169,0,75,0,197,0,102,0,119,0,209,0,73,0,39,0,0,0,173,0,63,0,0,0,0,0,92,0,70,0,181,0,0,0,0,0,0,0,132,0,163,0,253,0,127,0,27,0,239,0,194,0,181,0,206,0,25,0,6,0,1,0,136,0,22,0,105,0,204,0,113,0,109,0,154,0,2,0,233,0,40,0,190,0,162,0,107,0,130,0,138,0,94,0,139,0,0,0,106,0,253,0,253,0,97,0,42,0,208,0,62,0,0,0,22,0,171,0,22,0,241,0,189,0,0,0,130,0,0,0,0,0,0,0,220,0,67,0,235,0,31,0,0,0,9,0,164,0,189,0,237,0,132,0,0,0,244,0,150,0,253,0,146,0,66,0,0,0,251,0,110,0,105,0,168,0,0,0,79,0,226,0,5,0,10,0,137,0,188,0,0,0,0,0,203,0,193,0,90,0,31,0,4,0,230,0,212,0,21,0,222,0,0,0,209,0,223,0,63,0,108,0,60,0,22,0,128,0,39,0,0,0,0,0,11,0,93,0,0,0,114,0,230,0,112,0,128,0,46,0,0,0,83,0,66,0,10,0,161,0,196,0,6,0,59,0,188,0,191,0,253,0,0,0,255,0,0,0,193,0,145,0,6,0,123,0,124,0,0,0,178,0,37,0,160,0,235,0,120,0,0,0,71,0,0,0,230,0,111,0,0,0,200,0,53,0,91,0,132,0,178,0,210,0,130,0,117,0,0,0,147,0,136,0,174,0,143,0,29,0,0,0,106,0,77,0,58,0,41,0,81,0,201,0,169,0,206,0,112,0,207,0,0,0,4,0,224,0,200,0,0,0,40,0,243,0,40,0,31,0,106,0,193,0,94,0,15,0,0,0,0,0,86,0,76,0,37,0,29,0,0,0,0,0,103,0,182,0,0,0,253,0,188,0,212,0,159,0,216,0,83,0,31,0,101,0,87,0,175,0,119,0,247,0,240,0,39,0);
signal scenario_full  : scenario_type := (0,0,0,0,159,31,12,31,12,30,87,31,43,31,106,31,50,31,50,30,101,31,178,31,178,30,178,29,144,31,149,31,221,31,221,30,187,31,87,31,191,31,218,31,157,31,159,31,11,31,224,31,127,31,248,31,199,31,14,31,196,31,159,31,148,31,156,31,172,31,63,31,234,31,182,31,245,31,245,30,104,31,130,31,143,31,143,30,143,29,168,31,47,31,47,30,47,29,196,31,41,31,41,30,206,31,142,31,142,30,142,29,47,31,45,31,50,31,94,31,94,30,255,31,179,31,116,31,227,31,195,31,169,31,60,31,234,31,253,31,253,30,143,31,243,31,129,31,197,31,4,31,9,31,250,31,196,31,60,31,60,30,204,31,13,31,128,31,128,30,208,31,33,31,181,31,181,30,181,29,87,31,73,31,234,31,234,30,234,29,137,31,227,31,204,31,255,31,32,31,32,30,32,29,61,31,65,31,4,31,231,31,67,31,40,31,79,31,93,31,245,31,143,31,105,31,105,30,135,31,248,31,248,30,183,31,183,30,47,31,236,31,169,31,75,31,197,31,102,31,119,31,209,31,73,31,39,31,39,30,173,31,63,31,63,30,63,29,92,31,70,31,181,31,181,30,181,29,181,28,132,31,163,31,253,31,127,31,27,31,239,31,194,31,181,31,206,31,25,31,6,31,1,31,136,31,22,31,105,31,204,31,113,31,109,31,154,31,2,31,233,31,40,31,190,31,162,31,107,31,130,31,138,31,94,31,139,31,139,30,106,31,253,31,253,31,97,31,42,31,208,31,62,31,62,30,22,31,171,31,22,31,241,31,189,31,189,30,130,31,130,30,130,29,130,28,220,31,67,31,235,31,31,31,31,30,9,31,164,31,189,31,237,31,132,31,132,30,244,31,150,31,253,31,146,31,66,31,66,30,251,31,110,31,105,31,168,31,168,30,79,31,226,31,5,31,10,31,137,31,188,31,188,30,188,29,203,31,193,31,90,31,31,31,4,31,230,31,212,31,21,31,222,31,222,30,209,31,223,31,63,31,108,31,60,31,22,31,128,31,39,31,39,30,39,29,11,31,93,31,93,30,114,31,230,31,112,31,128,31,46,31,46,30,83,31,66,31,10,31,161,31,196,31,6,31,59,31,188,31,191,31,253,31,253,30,255,31,255,30,193,31,145,31,6,31,123,31,124,31,124,30,178,31,37,31,160,31,235,31,120,31,120,30,71,31,71,30,230,31,111,31,111,30,200,31,53,31,91,31,132,31,178,31,210,31,130,31,117,31,117,30,147,31,136,31,174,31,143,31,29,31,29,30,106,31,77,31,58,31,41,31,81,31,201,31,169,31,206,31,112,31,207,31,207,30,4,31,224,31,200,31,200,30,40,31,243,31,40,31,31,31,106,31,193,31,94,31,15,31,15,30,15,29,86,31,76,31,37,31,29,31,29,30,29,29,103,31,182,31,182,30,253,31,188,31,212,31,159,31,216,31,83,31,31,31,101,31,87,31,175,31,119,31,247,31,240,31,39,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
