-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 990;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (40,0,114,0,28,0,123,0,68,0,0,0,0,0,131,0,114,0,77,0,6,0,122,0,0,0,254,0,77,0,208,0,213,0,0,0,195,0,8,0,0,0,130,0,57,0,51,0,0,0,76,0,89,0,244,0,27,0,0,0,23,0,12,0,255,0,147,0,237,0,100,0,85,0,165,0,9,0,0,0,244,0,180,0,140,0,239,0,0,0,93,0,161,0,50,0,120,0,56,0,0,0,77,0,3,0,214,0,174,0,225,0,249,0,250,0,0,0,0,0,141,0,218,0,0,0,0,0,109,0,188,0,199,0,34,0,169,0,0,0,206,0,157,0,70,0,158,0,0,0,47,0,0,0,102,0,240,0,134,0,98,0,186,0,185,0,145,0,226,0,161,0,104,0,173,0,77,0,79,0,71,0,245,0,0,0,235,0,35,0,0,0,0,0,50,0,220,0,108,0,155,0,225,0,0,0,74,0,94,0,27,0,48,0,178,0,209,0,0,0,0,0,60,0,0,0,69,0,155,0,224,0,99,0,0,0,0,0,64,0,160,0,11,0,231,0,0,0,50,0,0,0,140,0,171,0,102,0,27,0,217,0,250,0,250,0,0,0,213,0,87,0,11,0,0,0,141,0,65,0,0,0,114,0,88,0,79,0,88,0,205,0,176,0,80,0,144,0,0,0,144,0,56,0,2,0,0,0,211,0,185,0,0,0,255,0,15,0,116,0,3,0,104,0,46,0,255,0,234,0,0,0,0,0,255,0,226,0,0,0,48,0,242,0,218,0,24,0,32,0,64,0,240,0,0,0,2,0,42,0,57,0,109,0,0,0,84,0,59,0,138,0,225,0,187,0,9,0,0,0,156,0,0,0,77,0,64,0,126,0,143,0,72,0,189,0,104,0,167,0,0,0,26,0,132,0,158,0,221,0,0,0,54,0,19,0,27,0,0,0,0,0,239,0,233,0,249,0,241,0,202,0,63,0,141,0,41,0,250,0,0,0,92,0,103,0,186,0,154,0,175,0,145,0,0,0,2,0,182,0,203,0,140,0,215,0,155,0,139,0,144,0,27,0,0,0,220,0,35,0,239,0,142,0,182,0,0,0,245,0,126,0,254,0,110,0,106,0,157,0,244,0,105,0,0,0,216,0,70,0,59,0,0,0,12,0,80,0,58,0,32,0,0,0,0,0,0,0,111,0,199,0,0,0,40,0,100,0,150,0,139,0,79,0,51,0,0,0,181,0,179,0,124,0,0,0,128,0,37,0,141,0,0,0,125,0,196,0,201,0,26,0,176,0,59,0,0,0,224,0,222,0,216,0,15,0,182,0,0,0,216,0,56,0,0,0,0,0,35,0,156,0,169,0,0,0,195,0,4,0,9,0,122,0,201,0,86,0,24,0,0,0,148,0,6,0,10,0,8,0,189,0,0,0,0,0,231,0,0,0,0,0,95,0,40,0,47,0,0,0,67,0,57,0,224,0,127,0,208,0,2,0,0,0,0,0,81,0,83,0,55,0,172,0,155,0,151,0,150,0,31,0,74,0,0,0,0,0,52,0,90,0,220,0,131,0,218,0,188,0,62,0,2,0,214,0,0,0,137,0,80,0,188,0,189,0,227,0,223,0,0,0,150,0,24,0,94,0,200,0,0,0,91,0,122,0,143,0,0,0,219,0,0,0,162,0,248,0,70,0,83,0,251,0,52,0,26,0,0,0,254,0,82,0,13,0,33,0,168,0,254,0,74,0,237,0,78,0,0,0,109,0,147,0,10,0,200,0,13,0,130,0,0,0,206,0,192,0,186,0,205,0,181,0,50,0,26,0,99,0,169,0,235,0,252,0,0,0,123,0,207,0,245,0,2,0,163,0,237,0,91,0,108,0,33,0,29,0,119,0,76,0,209,0,0,0,90,0,0,0,0,0,192,0,0,0,0,0,91,0,163,0,20,0,0,0,25,0,17,0,140,0,195,0,63,0,17,0,123,0,108,0,0,0,26,0,248,0,96,0,237,0,131,0,193,0,85,0,68,0,0,0,100,0,108,0,94,0,166,0,206,0,102,0,0,0,241,0,222,0,151,0,225,0,43,0,0,0,78,0,112,0,0,0,11,0,68,0,185,0,0,0,198,0,243,0,239,0,72,0,120,0,94,0,99,0,0,0,196,0,98,0,113,0,81,0,40,0,151,0,166,0,140,0,0,0,183,0,5,0,34,0,166,0,0,0,238,0,0,0,245,0,217,0,24,0,80,0,118,0,81,0,114,0,10,0,200,0,246,0,0,0,224,0,0,0,0,0,54,0,153,0,0,0,51,0,228,0,75,0,214,0,0,0,157,0,195,0,212,0,227,0,140,0,221,0,20,0,0,0,0,0,0,0,86,0,0,0,194,0,0,0,80,0,240,0,3,0,0,0,140,0,69,0,164,0,119,0,0,0,0,0,116,0,101,0,133,0,250,0,60,0,82,0,146,0,0,0,0,0,74,0,191,0,0,0,211,0,156,0,161,0,22,0,1,0,0,0,0,0,0,0,106,0,121,0,157,0,34,0,126,0,0,0,42,0,8,0,0,0,61,0,54,0,177,0,159,0,241,0,128,0,182,0,192,0,111,0,212,0,184,0,0,0,14,0,0,0,0,0,23,0,47,0,202,0,0,0,113,0,0,0,187,0,48,0,132,0,0,0,108,0,68,0,16,0,102,0,23,0,32,0,141,0,137,0,118,0,47,0,128,0,29,0,91,0,120,0,70,0,179,0,185,0,227,0,216,0,103,0,145,0,238,0,248,0,141,0,58,0,240,0,188,0,88,0,0,0,0,0,0,0,219,0,129,0,48,0,106,0,206,0,66,0,29,0,68,0,102,0,106,0,98,0,147,0,235,0,209,0,48,0,179,0,179,0,171,0,174,0,15,0,12,0,16,0,16,0,198,0,219,0,96,0,145,0,117,0,164,0,135,0,0,0,0,0,0,0,250,0,252,0,149,0,114,0,0,0,74,0,180,0,239,0,203,0,68,0,43,0,0,0,24,0,190,0,105,0,0,0,102,0,213,0,104,0,0,0,15,0,0,0,36,0,53,0,208,0,216,0,24,0,244,0,0,0,93,0,0,0,0,0,173,0,246,0,34,0,167,0,240,0,141,0,226,0,49,0,55,0,83,0,31,0,160,0,143,0,107,0,211,0,164,0,11,0,188,0,156,0,0,0,35,0,174,0,37,0,0,0,179,0,103,0,236,0,244,0,224,0,113,0,7,0,0,0,140,0,122,0,204,0,212,0,68,0,189,0,153,0,153,0,0,0,104,0,0,0,99,0,0,0,55,0,62,0,187,0,237,0,181,0,21,0,174,0,92,0,158,0,211,0,0,0,101,0,200,0,0,0,80,0,160,0,1,0,161,0,226,0,64,0,179,0,243,0,191,0,25,0,0,0,201,0,241,0,0,0,0,0,0,0,0,0,134,0,56,0,219,0,148,0,192,0,130,0,208,0,226,0,100,0,0,0,97,0,124,0,215,0,242,0,0,0,157,0,0,0,212,0,165,0,108,0,0,0,238,0,163,0,0,0,21,0,208,0,0,0,2,0,0,0,79,0,0,0,0,0,0,0,130,0,72,0,49,0,51,0,130,0,0,0,86,0,145,0,179,0,0,0,87,0,210,0,226,0,0,0,73,0,65,0,128,0,11,0,33,0,43,0,19,0,146,0,0,0,133,0,57,0,150,0,217,0,233,0,12,0,14,0,14,0,67,0,0,0,0,0,184,0,2,0,114,0,51,0,69,0,49,0,143,0,24,0,100,0,183,0,0,0,204,0,217,0,62,0,45,0,139,0,118,0,163,0,159,0,184,0,0,0,247,0,0,0,8,0,189,0,144,0,148,0,92,0,15,0,41,0,132,0,232,0,146,0,76,0,0,0,52,0,138,0,0,0,89,0,170,0,15,0,29,0,181,0,0,0,0,0,99,0,43,0,8,0,194,0,52,0,0,0,143,0,82,0,78,0,219,0,43,0,150,0,213,0,0,0,159,0,0,0,0,0,28,0,222,0,0,0,87,0,65,0,87,0,23,0,106,0,8,0,0,0,68,0,153,0,0,0,134,0,19,0,116,0,238,0,53,0,102,0,0,0,124,0,57,0,72,0,12,0,0,0,243,0,0,0,0,0,154,0,182,0,67,0,50,0,206,0,245,0,168,0,237,0,134,0,116,0,197,0,0,0,31,0,28,0,185,0,62,0,209,0,209,0,106,0,179,0,116,0,245,0,239,0,0,0,221,0,123,0,0,0,0,0,233,0,0,0,88,0,87,0,0,0,155,0,231,0,101,0,187,0,0,0,3,0,232,0,31,0,149,0,62,0,205,0,39,0,14,0,0,0,130,0,10,0,136,0,124,0,125,0,98,0,29,0,40,0,21,0,166,0,0,0,115,0,200,0,0,0,21,0,0,0,0,0,91,0,0,0);
signal scenario_full  : scenario_type := (40,31,114,31,28,31,123,31,68,31,68,30,68,29,131,31,114,31,77,31,6,31,122,31,122,30,254,31,77,31,208,31,213,31,213,30,195,31,8,31,8,30,130,31,57,31,51,31,51,30,76,31,89,31,244,31,27,31,27,30,23,31,12,31,255,31,147,31,237,31,100,31,85,31,165,31,9,31,9,30,244,31,180,31,140,31,239,31,239,30,93,31,161,31,50,31,120,31,56,31,56,30,77,31,3,31,214,31,174,31,225,31,249,31,250,31,250,30,250,29,141,31,218,31,218,30,218,29,109,31,188,31,199,31,34,31,169,31,169,30,206,31,157,31,70,31,158,31,158,30,47,31,47,30,102,31,240,31,134,31,98,31,186,31,185,31,145,31,226,31,161,31,104,31,173,31,77,31,79,31,71,31,245,31,245,30,235,31,35,31,35,30,35,29,50,31,220,31,108,31,155,31,225,31,225,30,74,31,94,31,27,31,48,31,178,31,209,31,209,30,209,29,60,31,60,30,69,31,155,31,224,31,99,31,99,30,99,29,64,31,160,31,11,31,231,31,231,30,50,31,50,30,140,31,171,31,102,31,27,31,217,31,250,31,250,31,250,30,213,31,87,31,11,31,11,30,141,31,65,31,65,30,114,31,88,31,79,31,88,31,205,31,176,31,80,31,144,31,144,30,144,31,56,31,2,31,2,30,211,31,185,31,185,30,255,31,15,31,116,31,3,31,104,31,46,31,255,31,234,31,234,30,234,29,255,31,226,31,226,30,48,31,242,31,218,31,24,31,32,31,64,31,240,31,240,30,2,31,42,31,57,31,109,31,109,30,84,31,59,31,138,31,225,31,187,31,9,31,9,30,156,31,156,30,77,31,64,31,126,31,143,31,72,31,189,31,104,31,167,31,167,30,26,31,132,31,158,31,221,31,221,30,54,31,19,31,27,31,27,30,27,29,239,31,233,31,249,31,241,31,202,31,63,31,141,31,41,31,250,31,250,30,92,31,103,31,186,31,154,31,175,31,145,31,145,30,2,31,182,31,203,31,140,31,215,31,155,31,139,31,144,31,27,31,27,30,220,31,35,31,239,31,142,31,182,31,182,30,245,31,126,31,254,31,110,31,106,31,157,31,244,31,105,31,105,30,216,31,70,31,59,31,59,30,12,31,80,31,58,31,32,31,32,30,32,29,32,28,111,31,199,31,199,30,40,31,100,31,150,31,139,31,79,31,51,31,51,30,181,31,179,31,124,31,124,30,128,31,37,31,141,31,141,30,125,31,196,31,201,31,26,31,176,31,59,31,59,30,224,31,222,31,216,31,15,31,182,31,182,30,216,31,56,31,56,30,56,29,35,31,156,31,169,31,169,30,195,31,4,31,9,31,122,31,201,31,86,31,24,31,24,30,148,31,6,31,10,31,8,31,189,31,189,30,189,29,231,31,231,30,231,29,95,31,40,31,47,31,47,30,67,31,57,31,224,31,127,31,208,31,2,31,2,30,2,29,81,31,83,31,55,31,172,31,155,31,151,31,150,31,31,31,74,31,74,30,74,29,52,31,90,31,220,31,131,31,218,31,188,31,62,31,2,31,214,31,214,30,137,31,80,31,188,31,189,31,227,31,223,31,223,30,150,31,24,31,94,31,200,31,200,30,91,31,122,31,143,31,143,30,219,31,219,30,162,31,248,31,70,31,83,31,251,31,52,31,26,31,26,30,254,31,82,31,13,31,33,31,168,31,254,31,74,31,237,31,78,31,78,30,109,31,147,31,10,31,200,31,13,31,130,31,130,30,206,31,192,31,186,31,205,31,181,31,50,31,26,31,99,31,169,31,235,31,252,31,252,30,123,31,207,31,245,31,2,31,163,31,237,31,91,31,108,31,33,31,29,31,119,31,76,31,209,31,209,30,90,31,90,30,90,29,192,31,192,30,192,29,91,31,163,31,20,31,20,30,25,31,17,31,140,31,195,31,63,31,17,31,123,31,108,31,108,30,26,31,248,31,96,31,237,31,131,31,193,31,85,31,68,31,68,30,100,31,108,31,94,31,166,31,206,31,102,31,102,30,241,31,222,31,151,31,225,31,43,31,43,30,78,31,112,31,112,30,11,31,68,31,185,31,185,30,198,31,243,31,239,31,72,31,120,31,94,31,99,31,99,30,196,31,98,31,113,31,81,31,40,31,151,31,166,31,140,31,140,30,183,31,5,31,34,31,166,31,166,30,238,31,238,30,245,31,217,31,24,31,80,31,118,31,81,31,114,31,10,31,200,31,246,31,246,30,224,31,224,30,224,29,54,31,153,31,153,30,51,31,228,31,75,31,214,31,214,30,157,31,195,31,212,31,227,31,140,31,221,31,20,31,20,30,20,29,20,28,86,31,86,30,194,31,194,30,80,31,240,31,3,31,3,30,140,31,69,31,164,31,119,31,119,30,119,29,116,31,101,31,133,31,250,31,60,31,82,31,146,31,146,30,146,29,74,31,191,31,191,30,211,31,156,31,161,31,22,31,1,31,1,30,1,29,1,28,106,31,121,31,157,31,34,31,126,31,126,30,42,31,8,31,8,30,61,31,54,31,177,31,159,31,241,31,128,31,182,31,192,31,111,31,212,31,184,31,184,30,14,31,14,30,14,29,23,31,47,31,202,31,202,30,113,31,113,30,187,31,48,31,132,31,132,30,108,31,68,31,16,31,102,31,23,31,32,31,141,31,137,31,118,31,47,31,128,31,29,31,91,31,120,31,70,31,179,31,185,31,227,31,216,31,103,31,145,31,238,31,248,31,141,31,58,31,240,31,188,31,88,31,88,30,88,29,88,28,219,31,129,31,48,31,106,31,206,31,66,31,29,31,68,31,102,31,106,31,98,31,147,31,235,31,209,31,48,31,179,31,179,31,171,31,174,31,15,31,12,31,16,31,16,31,198,31,219,31,96,31,145,31,117,31,164,31,135,31,135,30,135,29,135,28,250,31,252,31,149,31,114,31,114,30,74,31,180,31,239,31,203,31,68,31,43,31,43,30,24,31,190,31,105,31,105,30,102,31,213,31,104,31,104,30,15,31,15,30,36,31,53,31,208,31,216,31,24,31,244,31,244,30,93,31,93,30,93,29,173,31,246,31,34,31,167,31,240,31,141,31,226,31,49,31,55,31,83,31,31,31,160,31,143,31,107,31,211,31,164,31,11,31,188,31,156,31,156,30,35,31,174,31,37,31,37,30,179,31,103,31,236,31,244,31,224,31,113,31,7,31,7,30,140,31,122,31,204,31,212,31,68,31,189,31,153,31,153,31,153,30,104,31,104,30,99,31,99,30,55,31,62,31,187,31,237,31,181,31,21,31,174,31,92,31,158,31,211,31,211,30,101,31,200,31,200,30,80,31,160,31,1,31,161,31,226,31,64,31,179,31,243,31,191,31,25,31,25,30,201,31,241,31,241,30,241,29,241,28,241,27,134,31,56,31,219,31,148,31,192,31,130,31,208,31,226,31,100,31,100,30,97,31,124,31,215,31,242,31,242,30,157,31,157,30,212,31,165,31,108,31,108,30,238,31,163,31,163,30,21,31,208,31,208,30,2,31,2,30,79,31,79,30,79,29,79,28,130,31,72,31,49,31,51,31,130,31,130,30,86,31,145,31,179,31,179,30,87,31,210,31,226,31,226,30,73,31,65,31,128,31,11,31,33,31,43,31,19,31,146,31,146,30,133,31,57,31,150,31,217,31,233,31,12,31,14,31,14,31,67,31,67,30,67,29,184,31,2,31,114,31,51,31,69,31,49,31,143,31,24,31,100,31,183,31,183,30,204,31,217,31,62,31,45,31,139,31,118,31,163,31,159,31,184,31,184,30,247,31,247,30,8,31,189,31,144,31,148,31,92,31,15,31,41,31,132,31,232,31,146,31,76,31,76,30,52,31,138,31,138,30,89,31,170,31,15,31,29,31,181,31,181,30,181,29,99,31,43,31,8,31,194,31,52,31,52,30,143,31,82,31,78,31,219,31,43,31,150,31,213,31,213,30,159,31,159,30,159,29,28,31,222,31,222,30,87,31,65,31,87,31,23,31,106,31,8,31,8,30,68,31,153,31,153,30,134,31,19,31,116,31,238,31,53,31,102,31,102,30,124,31,57,31,72,31,12,31,12,30,243,31,243,30,243,29,154,31,182,31,67,31,50,31,206,31,245,31,168,31,237,31,134,31,116,31,197,31,197,30,31,31,28,31,185,31,62,31,209,31,209,31,106,31,179,31,116,31,245,31,239,31,239,30,221,31,123,31,123,30,123,29,233,31,233,30,88,31,87,31,87,30,155,31,231,31,101,31,187,31,187,30,3,31,232,31,31,31,149,31,62,31,205,31,39,31,14,31,14,30,130,31,10,31,136,31,124,31,125,31,98,31,29,31,40,31,21,31,166,31,166,30,115,31,200,31,200,30,21,31,21,30,21,29,91,31,91,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
