-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 750;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (139,0,0,0,113,0,12,0,234,0,0,0,85,0,157,0,118,0,27,0,62,0,0,0,0,0,47,0,0,0,0,0,250,0,146,0,63,0,115,0,20,0,0,0,49,0,66,0,136,0,142,0,0,0,64,0,43,0,242,0,82,0,10,0,247,0,52,0,12,0,187,0,207,0,78,0,0,0,220,0,251,0,228,0,192,0,169,0,0,0,114,0,39,0,134,0,0,0,112,0,200,0,196,0,0,0,16,0,186,0,0,0,102,0,21,0,227,0,99,0,77,0,89,0,199,0,136,0,27,0,0,0,166,0,0,0,0,0,142,0,104,0,77,0,0,0,106,0,203,0,223,0,0,0,255,0,63,0,64,0,92,0,227,0,213,0,188,0,47,0,0,0,0,0,1,0,135,0,182,0,37,0,5,0,0,0,68,0,57,0,244,0,181,0,223,0,237,0,244,0,166,0,0,0,57,0,233,0,215,0,149,0,158,0,144,0,195,0,24,0,0,0,231,0,124,0,89,0,52,0,0,0,191,0,0,0,212,0,100,0,213,0,0,0,0,0,220,0,146,0,34,0,153,0,129,0,27,0,125,0,146,0,121,0,197,0,31,0,135,0,165,0,182,0,200,0,71,0,159,0,183,0,90,0,0,0,82,0,161,0,8,0,244,0,151,0,173,0,214,0,206,0,0,0,247,0,0,0,200,0,69,0,14,0,182,0,37,0,45,0,0,0,180,0,74,0,83,0,32,0,37,0,48,0,162,0,110,0,218,0,93,0,138,0,170,0,113,0,230,0,0,0,244,0,0,0,40,0,196,0,11,0,48,0,0,0,250,0,6,0,120,0,32,0,156,0,175,0,182,0,0,0,167,0,207,0,0,0,0,0,72,0,76,0,176,0,0,0,30,0,131,0,4,0,226,0,186,0,212,0,98,0,63,0,0,0,199,0,0,0,101,0,80,0,155,0,107,0,193,0,0,0,71,0,92,0,15,0,209,0,52,0,57,0,219,0,38,0,127,0,164,0,38,0,221,0,128,0,230,0,123,0,231,0,167,0,45,0,106,0,0,0,0,0,201,0,0,0,122,0,216,0,254,0,115,0,109,0,0,0,135,0,61,0,245,0,85,0,0,0,77,0,115,0,246,0,204,0,244,0,114,0,196,0,0,0,227,0,175,0,247,0,0,0,0,0,25,0,73,0,130,0,14,0,89,0,30,0,124,0,87,0,184,0,96,0,0,0,61,0,0,0,47,0,36,0,227,0,27,0,84,0,0,0,10,0,95,0,90,0,99,0,171,0,9,0,189,0,217,0,28,0,212,0,175,0,207,0,253,0,5,0,188,0,0,0,61,0,21,0,83,0,86,0,188,0,0,0,0,0,0,0,239,0,0,0,229,0,250,0,192,0,48,0,252,0,216,0,0,0,128,0,22,0,21,0,76,0,16,0,112,0,101,0,107,0,0,0,92,0,204,0,63,0,176,0,171,0,0,0,50,0,81,0,118,0,56,0,160,0,248,0,0,0,51,0,0,0,251,0,185,0,0,0,87,0,50,0,235,0,57,0,63,0,140,0,0,0,75,0,0,0,7,0,99,0,218,0,98,0,188,0,36,0,116,0,104,0,77,0,99,0,81,0,0,0,39,0,190,0,203,0,0,0,235,0,133,0,91,0,130,0,0,0,197,0,190,0,0,0,0,0,40,0,33,0,72,0,220,0,23,0,0,0,21,0,161,0,0,0,198,0,0,0,171,0,160,0,0,0,125,0,31,0,59,0,162,0,210,0,170,0,223,0,177,0,93,0,137,0,109,0,0,0,11,0,0,0,49,0,0,0,0,0,209,0,31,0,0,0,109,0,228,0,54,0,165,0,250,0,26,0,0,0,43,0,149,0,35,0,249,0,157,0,253,0,181,0,90,0,75,0,0,0,87,0,42,0,52,0,233,0,107,0,184,0,106,0,150,0,63,0,0,0,222,0,8,0,0,0,181,0,0,0,249,0,183,0,17,0,253,0,104,0,0,0,95,0,183,0,175,0,4,0,206,0,161,0,225,0,233,0,175,0,195,0,0,0,172,0,191,0,0,0,57,0,0,0,71,0,0,0,0,0,0,0,203,0,68,0,95,0,106,0,237,0,0,0,149,0,255,0,0,0,207,0,0,0,125,0,188,0,242,0,0,0,0,0,101,0,240,0,92,0,20,0,222,0,103,0,0,0,72,0,50,0,92,0,113,0,104,0,24,0,40,0,223,0,0,0,0,0,242,0,0,0,200,0,82,0,189,0,164,0,108,0,6,0,255,0,0,0,0,0,155,0,232,0,0,0,0,0,23,0,200,0,0,0,67,0,232,0,161,0,202,0,22,0,207,0,238,0,37,0,0,0,0,0,73,0,158,0,224,0,168,0,144,0,103,0,170,0,217,0,0,0,76,0,176,0,28,0,57,0,117,0,61,0,151,0,177,0,35,0,92,0,0,0,106,0,206,0,113,0,8,0,0,0,149,0,142,0,66,0,0,0,37,0,96,0,97,0,37,0,28,0,230,0,27,0,197,0,196,0,216,0,220,0,64,0,209,0,50,0,33,0,1,0,0,0,218,0,63,0,9,0,150,0,201,0,135,0,63,0,11,0,97,0,219,0,212,0,52,0,85,0,105,0,0,0,217,0,16,0,0,0,0,0,92,0,202,0,0,0,0,0,218,0,143,0,78,0,122,0,0,0,112,0,169,0,0,0,179,0,0,0,120,0,129,0,22,0,0,0,168,0,129,0,189,0,27,0,53,0,118,0,0,0,21,0,0,0,0,0,0,0,48,0,219,0,94,0,0,0,120,0,169,0,168,0,0,0,19,0,0,0,77,0,15,0,0,0,146,0,0,0,7,0,206,0,209,0,11,0,0,0,0,0,225,0,46,0,16,0,11,0,231,0,51,0,62,0,8,0,0,0,135,0,106,0,33,0,0,0,5,0,0,0,144,0,32,0,0,0,124,0,33,0,95,0,10,0,3,0,11,0,0,0,253,0,202,0,139,0,242,0,0,0,0,0,249,0,210,0,25,0,158,0,255,0,84,0,0,0,0,0,78,0,0,0,215,0,189,0,99,0,0,0,108,0,212,0,194,0,195,0,225,0,0,0,62,0,20,0,2,0,0,0,113,0,90,0,0,0,253,0,112,0,154,0,142,0,0,0,0,0,181,0,176,0,134,0,124,0,15,0,0,0,216,0,120,0,0,0,255,0,141,0,0,0,69,0,215,0,221,0,28,0,72,0,169,0,237,0,9,0,38,0,0,0,0,0,57,0,142,0,0,0,99,0,115,0,0,0,3,0,63,0,56,0,61,0,143,0,0,0,110,0,0,0,43,0,208,0,180,0,220,0,99,0);
signal scenario_full  : scenario_type := (139,31,139,30,113,31,12,31,234,31,234,30,85,31,157,31,118,31,27,31,62,31,62,30,62,29,47,31,47,30,47,29,250,31,146,31,63,31,115,31,20,31,20,30,49,31,66,31,136,31,142,31,142,30,64,31,43,31,242,31,82,31,10,31,247,31,52,31,12,31,187,31,207,31,78,31,78,30,220,31,251,31,228,31,192,31,169,31,169,30,114,31,39,31,134,31,134,30,112,31,200,31,196,31,196,30,16,31,186,31,186,30,102,31,21,31,227,31,99,31,77,31,89,31,199,31,136,31,27,31,27,30,166,31,166,30,166,29,142,31,104,31,77,31,77,30,106,31,203,31,223,31,223,30,255,31,63,31,64,31,92,31,227,31,213,31,188,31,47,31,47,30,47,29,1,31,135,31,182,31,37,31,5,31,5,30,68,31,57,31,244,31,181,31,223,31,237,31,244,31,166,31,166,30,57,31,233,31,215,31,149,31,158,31,144,31,195,31,24,31,24,30,231,31,124,31,89,31,52,31,52,30,191,31,191,30,212,31,100,31,213,31,213,30,213,29,220,31,146,31,34,31,153,31,129,31,27,31,125,31,146,31,121,31,197,31,31,31,135,31,165,31,182,31,200,31,71,31,159,31,183,31,90,31,90,30,82,31,161,31,8,31,244,31,151,31,173,31,214,31,206,31,206,30,247,31,247,30,200,31,69,31,14,31,182,31,37,31,45,31,45,30,180,31,74,31,83,31,32,31,37,31,48,31,162,31,110,31,218,31,93,31,138,31,170,31,113,31,230,31,230,30,244,31,244,30,40,31,196,31,11,31,48,31,48,30,250,31,6,31,120,31,32,31,156,31,175,31,182,31,182,30,167,31,207,31,207,30,207,29,72,31,76,31,176,31,176,30,30,31,131,31,4,31,226,31,186,31,212,31,98,31,63,31,63,30,199,31,199,30,101,31,80,31,155,31,107,31,193,31,193,30,71,31,92,31,15,31,209,31,52,31,57,31,219,31,38,31,127,31,164,31,38,31,221,31,128,31,230,31,123,31,231,31,167,31,45,31,106,31,106,30,106,29,201,31,201,30,122,31,216,31,254,31,115,31,109,31,109,30,135,31,61,31,245,31,85,31,85,30,77,31,115,31,246,31,204,31,244,31,114,31,196,31,196,30,227,31,175,31,247,31,247,30,247,29,25,31,73,31,130,31,14,31,89,31,30,31,124,31,87,31,184,31,96,31,96,30,61,31,61,30,47,31,36,31,227,31,27,31,84,31,84,30,10,31,95,31,90,31,99,31,171,31,9,31,189,31,217,31,28,31,212,31,175,31,207,31,253,31,5,31,188,31,188,30,61,31,21,31,83,31,86,31,188,31,188,30,188,29,188,28,239,31,239,30,229,31,250,31,192,31,48,31,252,31,216,31,216,30,128,31,22,31,21,31,76,31,16,31,112,31,101,31,107,31,107,30,92,31,204,31,63,31,176,31,171,31,171,30,50,31,81,31,118,31,56,31,160,31,248,31,248,30,51,31,51,30,251,31,185,31,185,30,87,31,50,31,235,31,57,31,63,31,140,31,140,30,75,31,75,30,7,31,99,31,218,31,98,31,188,31,36,31,116,31,104,31,77,31,99,31,81,31,81,30,39,31,190,31,203,31,203,30,235,31,133,31,91,31,130,31,130,30,197,31,190,31,190,30,190,29,40,31,33,31,72,31,220,31,23,31,23,30,21,31,161,31,161,30,198,31,198,30,171,31,160,31,160,30,125,31,31,31,59,31,162,31,210,31,170,31,223,31,177,31,93,31,137,31,109,31,109,30,11,31,11,30,49,31,49,30,49,29,209,31,31,31,31,30,109,31,228,31,54,31,165,31,250,31,26,31,26,30,43,31,149,31,35,31,249,31,157,31,253,31,181,31,90,31,75,31,75,30,87,31,42,31,52,31,233,31,107,31,184,31,106,31,150,31,63,31,63,30,222,31,8,31,8,30,181,31,181,30,249,31,183,31,17,31,253,31,104,31,104,30,95,31,183,31,175,31,4,31,206,31,161,31,225,31,233,31,175,31,195,31,195,30,172,31,191,31,191,30,57,31,57,30,71,31,71,30,71,29,71,28,203,31,68,31,95,31,106,31,237,31,237,30,149,31,255,31,255,30,207,31,207,30,125,31,188,31,242,31,242,30,242,29,101,31,240,31,92,31,20,31,222,31,103,31,103,30,72,31,50,31,92,31,113,31,104,31,24,31,40,31,223,31,223,30,223,29,242,31,242,30,200,31,82,31,189,31,164,31,108,31,6,31,255,31,255,30,255,29,155,31,232,31,232,30,232,29,23,31,200,31,200,30,67,31,232,31,161,31,202,31,22,31,207,31,238,31,37,31,37,30,37,29,73,31,158,31,224,31,168,31,144,31,103,31,170,31,217,31,217,30,76,31,176,31,28,31,57,31,117,31,61,31,151,31,177,31,35,31,92,31,92,30,106,31,206,31,113,31,8,31,8,30,149,31,142,31,66,31,66,30,37,31,96,31,97,31,37,31,28,31,230,31,27,31,197,31,196,31,216,31,220,31,64,31,209,31,50,31,33,31,1,31,1,30,218,31,63,31,9,31,150,31,201,31,135,31,63,31,11,31,97,31,219,31,212,31,52,31,85,31,105,31,105,30,217,31,16,31,16,30,16,29,92,31,202,31,202,30,202,29,218,31,143,31,78,31,122,31,122,30,112,31,169,31,169,30,179,31,179,30,120,31,129,31,22,31,22,30,168,31,129,31,189,31,27,31,53,31,118,31,118,30,21,31,21,30,21,29,21,28,48,31,219,31,94,31,94,30,120,31,169,31,168,31,168,30,19,31,19,30,77,31,15,31,15,30,146,31,146,30,7,31,206,31,209,31,11,31,11,30,11,29,225,31,46,31,16,31,11,31,231,31,51,31,62,31,8,31,8,30,135,31,106,31,33,31,33,30,5,31,5,30,144,31,32,31,32,30,124,31,33,31,95,31,10,31,3,31,11,31,11,30,253,31,202,31,139,31,242,31,242,30,242,29,249,31,210,31,25,31,158,31,255,31,84,31,84,30,84,29,78,31,78,30,215,31,189,31,99,31,99,30,108,31,212,31,194,31,195,31,225,31,225,30,62,31,20,31,2,31,2,30,113,31,90,31,90,30,253,31,112,31,154,31,142,31,142,30,142,29,181,31,176,31,134,31,124,31,15,31,15,30,216,31,120,31,120,30,255,31,141,31,141,30,69,31,215,31,221,31,28,31,72,31,169,31,237,31,9,31,38,31,38,30,38,29,57,31,142,31,142,30,99,31,115,31,115,30,3,31,63,31,56,31,61,31,143,31,143,30,110,31,110,30,43,31,208,31,180,31,220,31,99,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
