-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 218;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (123,0,241,0,0,0,0,0,20,0,0,0,0,0,185,0,241,0,0,0,244,0,33,0,108,0,11,0,83,0,70,0,112,0,70,0,140,0,192,0,93,0,116,0,119,0,0,0,93,0,176,0,37,0,49,0,0,0,0,0,3,0,0,0,0,0,206,0,94,0,88,0,106,0,71,0,0,0,0,0,250,0,222,0,20,0,164,0,0,0,211,0,0,0,69,0,246,0,199,0,0,0,87,0,0,0,60,0,191,0,226,0,39,0,10,0,133,0,0,0,156,0,0,0,243,0,166,0,245,0,87,0,183,0,202,0,150,0,43,0,26,0,224,0,207,0,206,0,0,0,0,0,114,0,57,0,65,0,193,0,155,0,57,0,0,0,0,0,148,0,199,0,0,0,33,0,253,0,182,0,47,0,0,0,168,0,76,0,9,0,166,0,222,0,93,0,168,0,167,0,0,0,106,0,0,0,0,0,64,0,71,0,220,0,162,0,225,0,145,0,241,0,230,0,224,0,64,0,221,0,0,0,89,0,122,0,21,0,212,0,0,0,194,0,0,0,101,0,51,0,231,0,167,0,142,0,91,0,176,0,23,0,0,0,45,0,12,0,101,0,222,0,252,0,239,0,0,0,23,0,198,0,100,0,0,0,90,0,254,0,39,0,122,0,224,0,0,0,0,0,247,0,0,0,0,0,242,0,8,0,105,0,112,0,213,0,102,0,8,0,84,0,236,0,46,0,0,0,83,0,8,0,235,0,0,0,41,0,0,0,0,0,0,0,208,0,35,0,0,0,61,0,155,0,41,0,161,0,202,0,254,0,181,0,167,0,0,0,205,0,185,0,152,0,52,0,246,0,32,0,53,0,99,0,221,0,0,0,151,0,228,0,0,0,248,0,0,0,27,0,0,0,144,0,0,0,0,0,106,0,49,0,129,0,36,0,174,0,6,0,20,0,9,0,72,0,228,0,162,0,242,0,170,0,22,0);
signal scenario_full  : scenario_type := (123,31,241,31,241,30,241,29,20,31,20,30,20,29,185,31,241,31,241,30,244,31,33,31,108,31,11,31,83,31,70,31,112,31,70,31,140,31,192,31,93,31,116,31,119,31,119,30,93,31,176,31,37,31,49,31,49,30,49,29,3,31,3,30,3,29,206,31,94,31,88,31,106,31,71,31,71,30,71,29,250,31,222,31,20,31,164,31,164,30,211,31,211,30,69,31,246,31,199,31,199,30,87,31,87,30,60,31,191,31,226,31,39,31,10,31,133,31,133,30,156,31,156,30,243,31,166,31,245,31,87,31,183,31,202,31,150,31,43,31,26,31,224,31,207,31,206,31,206,30,206,29,114,31,57,31,65,31,193,31,155,31,57,31,57,30,57,29,148,31,199,31,199,30,33,31,253,31,182,31,47,31,47,30,168,31,76,31,9,31,166,31,222,31,93,31,168,31,167,31,167,30,106,31,106,30,106,29,64,31,71,31,220,31,162,31,225,31,145,31,241,31,230,31,224,31,64,31,221,31,221,30,89,31,122,31,21,31,212,31,212,30,194,31,194,30,101,31,51,31,231,31,167,31,142,31,91,31,176,31,23,31,23,30,45,31,12,31,101,31,222,31,252,31,239,31,239,30,23,31,198,31,100,31,100,30,90,31,254,31,39,31,122,31,224,31,224,30,224,29,247,31,247,30,247,29,242,31,8,31,105,31,112,31,213,31,102,31,8,31,84,31,236,31,46,31,46,30,83,31,8,31,235,31,235,30,41,31,41,30,41,29,41,28,208,31,35,31,35,30,61,31,155,31,41,31,161,31,202,31,254,31,181,31,167,31,167,30,205,31,185,31,152,31,52,31,246,31,32,31,53,31,99,31,221,31,221,30,151,31,228,31,228,30,248,31,248,30,27,31,27,30,144,31,144,30,144,29,106,31,49,31,129,31,36,31,174,31,6,31,20,31,9,31,72,31,228,31,162,31,242,31,170,31,22,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
