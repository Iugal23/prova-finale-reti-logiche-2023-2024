-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 781;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (248,0,254,0,249,0,0,0,0,0,0,0,145,0,131,0,45,0,144,0,77,0,42,0,172,0,247,0,14,0,135,0,251,0,163,0,171,0,73,0,0,0,152,0,0,0,89,0,31,0,84,0,189,0,0,0,191,0,115,0,142,0,246,0,209,0,224,0,57,0,0,0,135,0,198,0,0,0,0,0,186,0,0,0,170,0,13,0,182,0,24,0,200,0,223,0,109,0,0,0,122,0,192,0,229,0,176,0,129,0,51,0,23,0,111,0,155,0,3,0,224,0,0,0,29,0,76,0,123,0,42,0,101,0,106,0,3,0,153,0,53,0,147,0,255,0,0,0,168,0,0,0,246,0,24,0,52,0,72,0,137,0,194,0,145,0,157,0,95,0,194,0,92,0,142,0,215,0,160,0,207,0,0,0,28,0,81,0,160,0,0,0,13,0,147,0,228,0,61,0,130,0,197,0,82,0,252,0,40,0,14,0,58,0,218,0,15,0,124,0,0,0,0,0,212,0,203,0,0,0,0,0,65,0,226,0,0,0,32,0,242,0,0,0,251,0,1,0,32,0,1,0,151,0,100,0,68,0,218,0,28,0,182,0,237,0,33,0,60,0,193,0,219,0,154,0,138,0,248,0,236,0,138,0,159,0,64,0,8,0,153,0,0,0,18,0,171,0,147,0,0,0,12,0,164,0,12,0,58,0,154,0,103,0,23,0,165,0,5,0,155,0,135,0,0,0,41,0,209,0,21,0,47,0,218,0,74,0,54,0,0,0,181,0,188,0,64,0,0,0,67,0,223,0,48,0,47,0,184,0,202,0,105,0,237,0,34,0,0,0,53,0,0,0,153,0,81,0,181,0,115,0,0,0,200,0,251,0,121,0,0,0,131,0,116,0,242,0,125,0,108,0,249,0,71,0,216,0,65,0,73,0,89,0,43,0,11,0,69,0,202,0,2,0,0,0,149,0,172,0,23,0,0,0,16,0,231,0,60,0,215,0,125,0,118,0,246,0,135,0,0,0,198,0,187,0,0,0,70,0,0,0,119,0,0,0,208,0,222,0,189,0,234,0,0,0,49,0,139,0,231,0,0,0,185,0,218,0,2,0,249,0,142,0,106,0,88,0,33,0,156,0,199,0,253,0,157,0,113,0,49,0,224,0,32,0,222,0,40,0,0,0,152,0,182,0,125,0,170,0,83,0,183,0,137,0,176,0,49,0,110,0,0,0,0,0,198,0,89,0,0,0,91,0,0,0,73,0,15,0,23,0,0,0,0,0,0,0,110,0,249,0,231,0,62,0,211,0,97,0,255,0,34,0,0,0,89,0,65,0,177,0,51,0,5,0,95,0,40,0,0,0,231,0,10,0,42,0,239,0,183,0,125,0,242,0,90,0,60,0,0,0,176,0,201,0,0,0,0,0,25,0,133,0,0,0,0,0,227,0,205,0,174,0,177,0,255,0,85,0,110,0,124,0,251,0,135,0,26,0,0,0,3,0,235,0,198,0,0,0,139,0,96,0,149,0,206,0,18,0,28,0,228,0,192,0,19,0,0,0,70,0,175,0,0,0,0,0,182,0,211,0,27,0,238,0,107,0,0,0,34,0,249,0,24,0,50,0,186,0,178,0,0,0,232,0,0,0,33,0,179,0,167,0,204,0,95,0,242,0,27,0,0,0,127,0,110,0,14,0,0,0,159,0,159,0,133,0,254,0,140,0,152,0,1,0,147,0,205,0,0,0,0,0,65,0,254,0,0,0,116,0,175,0,107,0,150,0,57,0,173,0,149,0,222,0,0,0,179,0,29,0,99,0,21,0,92,0,92,0,129,0,0,0,247,0,220,0,106,0,0,0,226,0,0,0,84,0,136,0,161,0,90,0,194,0,2,0,125,0,50,0,148,0,38,0,76,0,137,0,42,0,0,0,218,0,167,0,194,0,0,0,0,0,0,0,213,0,211,0,37,0,246,0,118,0,179,0,82,0,51,0,86,0,240,0,196,0,0,0,0,0,72,0,118,0,0,0,232,0,0,0,142,0,73,0,175,0,170,0,62,0,130,0,101,0,40,0,179,0,169,0,0,0,144,0,157,0,166,0,103,0,0,0,4,0,121,0,133,0,0,0,131,0,234,0,21,0,0,0,0,0,254,0,149,0,213,0,126,0,85,0,0,0,202,0,252,0,180,0,113,0,48,0,13,0,201,0,253,0,0,0,0,0,0,0,0,0,4,0,0,0,104,0,209,0,0,0,135,0,0,0,193,0,13,0,0,0,166,0,149,0,28,0,18,0,0,0,173,0,0,0,0,0,98,0,0,0,161,0,50,0,22,0,225,0,205,0,12,0,0,0,166,0,176,0,150,0,220,0,170,0,41,0,50,0,56,0,205,0,218,0,46,0,242,0,228,0,246,0,106,0,37,0,0,0,246,0,39,0,169,0,149,0,115,0,48,0,108,0,54,0,79,0,0,0,255,0,30,0,0,0,74,0,122,0,0,0,41,0,205,0,176,0,250,0,157,0,216,0,180,0,98,0,120,0,27,0,143,0,159,0,130,0,7,0,72,0,186,0,33,0,0,0,71,0,0,0,96,0,174,0,195,0,50,0,146,0,178,0,0,0,0,0,0,0,0,0,73,0,107,0,53,0,61,0,129,0,107,0,0,0,239,0,0,0,0,0,188,0,99,0,232,0,0,0,65,0,233,0,0,0,0,0,48,0,0,0,110,0,187,0,78,0,228,0,0,0,210,0,0,0,0,0,0,0,206,0,172,0,90,0,70,0,183,0,0,0,222,0,243,0,0,0,227,0,221,0,29,0,109,0,79,0,0,0,113,0,187,0,143,0,221,0,174,0,0,0,0,0,197,0,219,0,0,0,214,0,0,0,0,0,109,0,55,0,124,0,0,0,169,0,0,0,123,0,0,0,233,0,54,0,163,0,81,0,174,0,231,0,0,0,0,0,51,0,75,0,45,0,132,0,51,0,157,0,109,0,194,0,21,0,0,0,181,0,67,0,81,0,244,0,3,0,118,0,163,0,25,0,76,0,173,0,47,0,31,0,236,0,60,0,244,0,239,0,0,0,57,0,190,0,135,0,0,0,0,0,168,0,106,0,213,0,33,0,0,0,100,0,81,0,254,0,199,0,161,0,208,0,55,0,81,0,241,0,20,0,74,0,176,0,145,0,0,0,226,0,237,0,253,0,0,0,66,0,93,0,217,0,153,0,174,0,155,0,0,0,0,0,18,0,202,0,0,0,199,0,0,0,153,0,163,0,211,0,130,0,184,0,179,0,208,0,141,0,205,0,7,0,28,0,135,0,72,0,144,0,22,0,96,0,229,0,161,0,0,0,50,0,12,0,174,0,43,0,51,0,221,0,187,0,58,0,125,0,190,0,219,0,0,0,154,0,224,0,168,0,142,0,32,0,197,0,99,0,179,0,63,0,245,0,138,0,204,0,247,0,135,0,166,0,12,0,0,0,54,0,132,0,66,0,79,0,134,0,149,0,181,0,201,0);
signal scenario_full  : scenario_type := (248,31,254,31,249,31,249,30,249,29,249,28,145,31,131,31,45,31,144,31,77,31,42,31,172,31,247,31,14,31,135,31,251,31,163,31,171,31,73,31,73,30,152,31,152,30,89,31,31,31,84,31,189,31,189,30,191,31,115,31,142,31,246,31,209,31,224,31,57,31,57,30,135,31,198,31,198,30,198,29,186,31,186,30,170,31,13,31,182,31,24,31,200,31,223,31,109,31,109,30,122,31,192,31,229,31,176,31,129,31,51,31,23,31,111,31,155,31,3,31,224,31,224,30,29,31,76,31,123,31,42,31,101,31,106,31,3,31,153,31,53,31,147,31,255,31,255,30,168,31,168,30,246,31,24,31,52,31,72,31,137,31,194,31,145,31,157,31,95,31,194,31,92,31,142,31,215,31,160,31,207,31,207,30,28,31,81,31,160,31,160,30,13,31,147,31,228,31,61,31,130,31,197,31,82,31,252,31,40,31,14,31,58,31,218,31,15,31,124,31,124,30,124,29,212,31,203,31,203,30,203,29,65,31,226,31,226,30,32,31,242,31,242,30,251,31,1,31,32,31,1,31,151,31,100,31,68,31,218,31,28,31,182,31,237,31,33,31,60,31,193,31,219,31,154,31,138,31,248,31,236,31,138,31,159,31,64,31,8,31,153,31,153,30,18,31,171,31,147,31,147,30,12,31,164,31,12,31,58,31,154,31,103,31,23,31,165,31,5,31,155,31,135,31,135,30,41,31,209,31,21,31,47,31,218,31,74,31,54,31,54,30,181,31,188,31,64,31,64,30,67,31,223,31,48,31,47,31,184,31,202,31,105,31,237,31,34,31,34,30,53,31,53,30,153,31,81,31,181,31,115,31,115,30,200,31,251,31,121,31,121,30,131,31,116,31,242,31,125,31,108,31,249,31,71,31,216,31,65,31,73,31,89,31,43,31,11,31,69,31,202,31,2,31,2,30,149,31,172,31,23,31,23,30,16,31,231,31,60,31,215,31,125,31,118,31,246,31,135,31,135,30,198,31,187,31,187,30,70,31,70,30,119,31,119,30,208,31,222,31,189,31,234,31,234,30,49,31,139,31,231,31,231,30,185,31,218,31,2,31,249,31,142,31,106,31,88,31,33,31,156,31,199,31,253,31,157,31,113,31,49,31,224,31,32,31,222,31,40,31,40,30,152,31,182,31,125,31,170,31,83,31,183,31,137,31,176,31,49,31,110,31,110,30,110,29,198,31,89,31,89,30,91,31,91,30,73,31,15,31,23,31,23,30,23,29,23,28,110,31,249,31,231,31,62,31,211,31,97,31,255,31,34,31,34,30,89,31,65,31,177,31,51,31,5,31,95,31,40,31,40,30,231,31,10,31,42,31,239,31,183,31,125,31,242,31,90,31,60,31,60,30,176,31,201,31,201,30,201,29,25,31,133,31,133,30,133,29,227,31,205,31,174,31,177,31,255,31,85,31,110,31,124,31,251,31,135,31,26,31,26,30,3,31,235,31,198,31,198,30,139,31,96,31,149,31,206,31,18,31,28,31,228,31,192,31,19,31,19,30,70,31,175,31,175,30,175,29,182,31,211,31,27,31,238,31,107,31,107,30,34,31,249,31,24,31,50,31,186,31,178,31,178,30,232,31,232,30,33,31,179,31,167,31,204,31,95,31,242,31,27,31,27,30,127,31,110,31,14,31,14,30,159,31,159,31,133,31,254,31,140,31,152,31,1,31,147,31,205,31,205,30,205,29,65,31,254,31,254,30,116,31,175,31,107,31,150,31,57,31,173,31,149,31,222,31,222,30,179,31,29,31,99,31,21,31,92,31,92,31,129,31,129,30,247,31,220,31,106,31,106,30,226,31,226,30,84,31,136,31,161,31,90,31,194,31,2,31,125,31,50,31,148,31,38,31,76,31,137,31,42,31,42,30,218,31,167,31,194,31,194,30,194,29,194,28,213,31,211,31,37,31,246,31,118,31,179,31,82,31,51,31,86,31,240,31,196,31,196,30,196,29,72,31,118,31,118,30,232,31,232,30,142,31,73,31,175,31,170,31,62,31,130,31,101,31,40,31,179,31,169,31,169,30,144,31,157,31,166,31,103,31,103,30,4,31,121,31,133,31,133,30,131,31,234,31,21,31,21,30,21,29,254,31,149,31,213,31,126,31,85,31,85,30,202,31,252,31,180,31,113,31,48,31,13,31,201,31,253,31,253,30,253,29,253,28,253,27,4,31,4,30,104,31,209,31,209,30,135,31,135,30,193,31,13,31,13,30,166,31,149,31,28,31,18,31,18,30,173,31,173,30,173,29,98,31,98,30,161,31,50,31,22,31,225,31,205,31,12,31,12,30,166,31,176,31,150,31,220,31,170,31,41,31,50,31,56,31,205,31,218,31,46,31,242,31,228,31,246,31,106,31,37,31,37,30,246,31,39,31,169,31,149,31,115,31,48,31,108,31,54,31,79,31,79,30,255,31,30,31,30,30,74,31,122,31,122,30,41,31,205,31,176,31,250,31,157,31,216,31,180,31,98,31,120,31,27,31,143,31,159,31,130,31,7,31,72,31,186,31,33,31,33,30,71,31,71,30,96,31,174,31,195,31,50,31,146,31,178,31,178,30,178,29,178,28,178,27,73,31,107,31,53,31,61,31,129,31,107,31,107,30,239,31,239,30,239,29,188,31,99,31,232,31,232,30,65,31,233,31,233,30,233,29,48,31,48,30,110,31,187,31,78,31,228,31,228,30,210,31,210,30,210,29,210,28,206,31,172,31,90,31,70,31,183,31,183,30,222,31,243,31,243,30,227,31,221,31,29,31,109,31,79,31,79,30,113,31,187,31,143,31,221,31,174,31,174,30,174,29,197,31,219,31,219,30,214,31,214,30,214,29,109,31,55,31,124,31,124,30,169,31,169,30,123,31,123,30,233,31,54,31,163,31,81,31,174,31,231,31,231,30,231,29,51,31,75,31,45,31,132,31,51,31,157,31,109,31,194,31,21,31,21,30,181,31,67,31,81,31,244,31,3,31,118,31,163,31,25,31,76,31,173,31,47,31,31,31,236,31,60,31,244,31,239,31,239,30,57,31,190,31,135,31,135,30,135,29,168,31,106,31,213,31,33,31,33,30,100,31,81,31,254,31,199,31,161,31,208,31,55,31,81,31,241,31,20,31,74,31,176,31,145,31,145,30,226,31,237,31,253,31,253,30,66,31,93,31,217,31,153,31,174,31,155,31,155,30,155,29,18,31,202,31,202,30,199,31,199,30,153,31,163,31,211,31,130,31,184,31,179,31,208,31,141,31,205,31,7,31,28,31,135,31,72,31,144,31,22,31,96,31,229,31,161,31,161,30,50,31,12,31,174,31,43,31,51,31,221,31,187,31,58,31,125,31,190,31,219,31,219,30,154,31,224,31,168,31,142,31,32,31,197,31,99,31,179,31,63,31,245,31,138,31,204,31,247,31,135,31,166,31,12,31,12,30,54,31,132,31,66,31,79,31,134,31,149,31,181,31,201,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
