-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 987;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,231,0,123,0,185,0,52,0,91,0,0,0,7,0,52,0,142,0,0,0,70,0,138,0,212,0,0,0,191,0,157,0,160,0,0,0,82,0,104,0,158,0,126,0,14,0,19,0,54,0,11,0,146,0,243,0,204,0,55,0,82,0,125,0,69,0,0,0,45,0,247,0,84,0,4,0,201,0,219,0,231,0,111,0,175,0,87,0,127,0,0,0,166,0,210,0,0,0,0,0,37,0,126,0,0,0,193,0,66,0,7,0,193,0,93,0,244,0,0,0,147,0,20,0,31,0,129,0,85,0,190,0,2,0,244,0,0,0,95,0,22,0,234,0,85,0,109,0,249,0,189,0,0,0,159,0,62,0,161,0,216,0,135,0,213,0,43,0,175,0,104,0,202,0,206,0,40,0,126,0,230,0,252,0,240,0,0,0,198,0,59,0,59,0,168,0,226,0,32,0,0,0,77,0,255,0,232,0,247,0,32,0,0,0,241,0,90,0,185,0,189,0,202,0,143,0,172,0,167,0,98,0,107,0,221,0,14,0,165,0,139,0,62,0,159,0,0,0,137,0,210,0,72,0,124,0,209,0,91,0,204,0,0,0,110,0,13,0,175,0,0,0,99,0,200,0,201,0,137,0,35,0,128,0,21,0,0,0,243,0,248,0,0,0,143,0,99,0,133,0,0,0,213,0,193,0,90,0,70,0,242,0,0,0,118,0,0,0,150,0,104,0,215,0,234,0,0,0,240,0,129,0,84,0,173,0,0,0,1,0,71,0,206,0,165,0,0,0,203,0,0,0,143,0,128,0,205,0,99,0,0,0,165,0,0,0,165,0,104,0,0,0,42,0,254,0,0,0,177,0,0,0,176,0,110,0,212,0,217,0,0,0,127,0,42,0,98,0,0,0,53,0,74,0,152,0,239,0,0,0,187,0,213,0,148,0,57,0,84,0,199,0,182,0,0,0,142,0,0,0,0,0,218,0,190,0,230,0,132,0,190,0,0,0,116,0,170,0,14,0,68,0,165,0,39,0,137,0,168,0,169,0,192,0,189,0,26,0,220,0,162,0,125,0,72,0,138,0,162,0,74,0,56,0,129,0,37,0,117,0,213,0,36,0,80,0,121,0,0,0,146,0,104,0,170,0,0,0,215,0,229,0,0,0,156,0,45,0,128,0,166,0,0,0,194,0,70,0,234,0,171,0,63,0,117,0,159,0,0,0,55,0,247,0,68,0,0,0,245,0,63,0,120,0,61,0,0,0,42,0,165,0,0,0,207,0,0,0,0,0,0,0,45,0,221,0,52,0,0,0,73,0,45,0,148,0,208,0,0,0,72,0,67,0,0,0,57,0,0,0,168,0,79,0,133,0,60,0,188,0,81,0,248,0,88,0,191,0,147,0,0,0,127,0,96,0,65,0,91,0,58,0,99,0,180,0,0,0,135,0,13,0,90,0,136,0,104,0,18,0,20,0,45,0,223,0,0,0,209,0,66,0,196,0,0,0,39,0,121,0,244,0,46,0,70,0,218,0,0,0,0,0,0,0,144,0,60,0,101,0,43,0,90,0,79,0,0,0,198,0,125,0,0,0,196,0,36,0,38,0,241,0,212,0,71,0,0,0,105,0,28,0,64,0,176,0,15,0,131,0,173,0,246,0,2,0,51,0,0,0,20,0,0,0,183,0,239,0,123,0,0,0,26,0,144,0,166,0,70,0,223,0,110,0,235,0,182,0,78,0,33,0,9,0,74,0,108,0,36,0,247,0,244,0,65,0,101,0,225,0,0,0,40,0,0,0,215,0,147,0,148,0,62,0,159,0,163,0,122,0,166,0,106,0,108,0,112,0,100,0,29,0,35,0,0,0,0,0,197,0,0,0,208,0,244,0,20,0,183,0,102,0,0,0,214,0,253,0,6,0,185,0,231,0,126,0,0,0,220,0,106,0,113,0,8,0,111,0,0,0,0,0,177,0,217,0,91,0,157,0,74,0,236,0,0,0,99,0,147,0,0,0,195,0,0,0,0,0,0,0,244,0,2,0,162,0,140,0,169,0,0,0,223,0,119,0,0,0,75,0,7,0,41,0,65,0,185,0,246,0,0,0,47,0,102,0,0,0,0,0,140,0,217,0,173,0,44,0,254,0,130,0,101,0,5,0,90,0,61,0,147,0,0,0,148,0,142,0,0,0,208,0,3,0,0,0,96,0,237,0,102,0,91,0,4,0,0,0,0,0,0,0,0,0,73,0,87,0,194,0,61,0,0,0,39,0,0,0,56,0,0,0,88,0,59,0,110,0,102,0,142,0,187,0,181,0,34,0,0,0,0,0,210,0,0,0,0,0,0,0,119,0,0,0,252,0,212,0,0,0,0,0,92,0,100,0,255,0,157,0,128,0,0,0,227,0,87,0,42,0,98,0,118,0,153,0,40,0,33,0,249,0,223,0,234,0,244,0,237,0,29,0,67,0,0,0,104,0,26,0,228,0,203,0,192,0,227,0,0,0,101,0,0,0,0,0,157,0,85,0,157,0,158,0,168,0,251,0,47,0,63,0,148,0,104,0,182,0,54,0,0,0,251,0,174,0,177,0,88,0,0,0,214,0,0,0,102,0,47,0,221,0,163,0,133,0,192,0,203,0,118,0,70,0,0,0,143,0,62,0,0,0,207,0,175,0,47,0,126,0,0,0,21,0,150,0,247,0,91,0,109,0,192,0,25,0,0,0,104,0,60,0,136,0,139,0,89,0,105,0,43,0,0,0,137,0,27,0,20,0,0,0,208,0,206,0,228,0,0,0,237,0,55,0,73,0,0,0,68,0,0,0,88,0,197,0,78,0,107,0,211,0,196,0,117,0,231,0,16,0,162,0,139,0,0,0,221,0,0,0,17,0,117,0,80,0,211,0,225,0,162,0,0,0,154,0,0,0,84,0,178,0,72,0,96,0,12,0,144,0,223,0,246,0,157,0,58,0,140,0,218,0,118,0,0,0,0,0,0,0,68,0,90,0,55,0,126,0,117,0,9,0,191,0,250,0,172,0,212,0,0,0,116,0,154,0,38,0,0,0,0,0,107,0,182,0,0,0,201,0,0,0,174,0,0,0,0,0,185,0,166,0,196,0,107,0,220,0,64,0,216,0,10,0,20,0,4,0,0,0,170,0,0,0,36,0,228,0,110,0,234,0,109,0,0,0,211,0,224,0,174,0,228,0,181,0,0,0,126,0,109,0,223,0,0,0,0,0,0,0,60,0,84,0,149,0,2,0,28,0,240,0,0,0,211,0,82,0,41,0,247,0,77,0,101,0,156,0,0,0,196,0,0,0,0,0,0,0,22,0,223,0,13,0,0,0,0,0,14,0,97,0,0,0,239,0,0,0,0,0,25,0,218,0,191,0,0,0,0,0,34,0,27,0,124,0,98,0,206,0,82,0,34,0,182,0,19,0,97,0,199,0,130,0,74,0,199,0,33,0,0,0,16,0,171,0,0,0,0,0,0,0,150,0,0,0,188,0,144,0,0,0,118,0,219,0,126,0,165,0,0,0,180,0,105,0,195,0,196,0,249,0,152,0,124,0,0,0,57,0,0,0,103,0,123,0,0,0,63,0,82,0,0,0,32,0,4,0,0,0,43,0,24,0,71,0,0,0,172,0,107,0,0,0,214,0,18,0,0,0,43,0,74,0,228,0,22,0,208,0,16,0,107,0,9,0,0,0,101,0,114,0,202,0,58,0,0,0,28,0,85,0,115,0,251,0,212,0,194,0,107,0,95,0,0,0,48,0,0,0,15,0,65,0,100,0,0,0,94,0,8,0,198,0,209,0,0,0,49,0,157,0,241,0,0,0,24,0,184,0,191,0,175,0,18,0,0,0,64,0,173,0,236,0,200,0,243,0,41,0,0,0,192,0,168,0,120,0,133,0,0,0,178,0,191,0,105,0,191,0,34,0,223,0,0,0,0,0,47,0,0,0,253,0,8,0,104,0,49,0,110,0,0,0,70,0,104,0,138,0,193,0,196,0,0,0,20,0,109,0,172,0,158,0,8,0,245,0,128,0,227,0,93,0,17,0,83,0,0,0,0,0,240,0,75,0,57,0,95,0,170,0,195,0,79,0,99,0,0,0,193,0,0,0,83,0,179,0,11,0,213,0,103,0,125,0,90,0,2,0,68,0,139,0,127,0,245,0,100,0,0,0,83,0,30,0,157,0,197,0,124,0,194,0,156,0,85,0,152,0,173,0,233,0,0,0,255,0,0,0,91,0,247,0,0,0,240,0,237,0,189,0,37,0,159,0,0,0,241,0,74,0,116,0,96,0,140,0,203,0,19,0,105,0,253,0,153,0,0,0,234,0,231,0,202,0,248,0,111,0,0,0,0,0,0,0,130,0,1,0,104,0,216,0,0,0,183,0,0,0,28,0,119,0,67,0,106,0,75,0,161,0);
signal scenario_full  : scenario_type := (0,0,231,31,123,31,185,31,52,31,91,31,91,30,7,31,52,31,142,31,142,30,70,31,138,31,212,31,212,30,191,31,157,31,160,31,160,30,82,31,104,31,158,31,126,31,14,31,19,31,54,31,11,31,146,31,243,31,204,31,55,31,82,31,125,31,69,31,69,30,45,31,247,31,84,31,4,31,201,31,219,31,231,31,111,31,175,31,87,31,127,31,127,30,166,31,210,31,210,30,210,29,37,31,126,31,126,30,193,31,66,31,7,31,193,31,93,31,244,31,244,30,147,31,20,31,31,31,129,31,85,31,190,31,2,31,244,31,244,30,95,31,22,31,234,31,85,31,109,31,249,31,189,31,189,30,159,31,62,31,161,31,216,31,135,31,213,31,43,31,175,31,104,31,202,31,206,31,40,31,126,31,230,31,252,31,240,31,240,30,198,31,59,31,59,31,168,31,226,31,32,31,32,30,77,31,255,31,232,31,247,31,32,31,32,30,241,31,90,31,185,31,189,31,202,31,143,31,172,31,167,31,98,31,107,31,221,31,14,31,165,31,139,31,62,31,159,31,159,30,137,31,210,31,72,31,124,31,209,31,91,31,204,31,204,30,110,31,13,31,175,31,175,30,99,31,200,31,201,31,137,31,35,31,128,31,21,31,21,30,243,31,248,31,248,30,143,31,99,31,133,31,133,30,213,31,193,31,90,31,70,31,242,31,242,30,118,31,118,30,150,31,104,31,215,31,234,31,234,30,240,31,129,31,84,31,173,31,173,30,1,31,71,31,206,31,165,31,165,30,203,31,203,30,143,31,128,31,205,31,99,31,99,30,165,31,165,30,165,31,104,31,104,30,42,31,254,31,254,30,177,31,177,30,176,31,110,31,212,31,217,31,217,30,127,31,42,31,98,31,98,30,53,31,74,31,152,31,239,31,239,30,187,31,213,31,148,31,57,31,84,31,199,31,182,31,182,30,142,31,142,30,142,29,218,31,190,31,230,31,132,31,190,31,190,30,116,31,170,31,14,31,68,31,165,31,39,31,137,31,168,31,169,31,192,31,189,31,26,31,220,31,162,31,125,31,72,31,138,31,162,31,74,31,56,31,129,31,37,31,117,31,213,31,36,31,80,31,121,31,121,30,146,31,104,31,170,31,170,30,215,31,229,31,229,30,156,31,45,31,128,31,166,31,166,30,194,31,70,31,234,31,171,31,63,31,117,31,159,31,159,30,55,31,247,31,68,31,68,30,245,31,63,31,120,31,61,31,61,30,42,31,165,31,165,30,207,31,207,30,207,29,207,28,45,31,221,31,52,31,52,30,73,31,45,31,148,31,208,31,208,30,72,31,67,31,67,30,57,31,57,30,168,31,79,31,133,31,60,31,188,31,81,31,248,31,88,31,191,31,147,31,147,30,127,31,96,31,65,31,91,31,58,31,99,31,180,31,180,30,135,31,13,31,90,31,136,31,104,31,18,31,20,31,45,31,223,31,223,30,209,31,66,31,196,31,196,30,39,31,121,31,244,31,46,31,70,31,218,31,218,30,218,29,218,28,144,31,60,31,101,31,43,31,90,31,79,31,79,30,198,31,125,31,125,30,196,31,36,31,38,31,241,31,212,31,71,31,71,30,105,31,28,31,64,31,176,31,15,31,131,31,173,31,246,31,2,31,51,31,51,30,20,31,20,30,183,31,239,31,123,31,123,30,26,31,144,31,166,31,70,31,223,31,110,31,235,31,182,31,78,31,33,31,9,31,74,31,108,31,36,31,247,31,244,31,65,31,101,31,225,31,225,30,40,31,40,30,215,31,147,31,148,31,62,31,159,31,163,31,122,31,166,31,106,31,108,31,112,31,100,31,29,31,35,31,35,30,35,29,197,31,197,30,208,31,244,31,20,31,183,31,102,31,102,30,214,31,253,31,6,31,185,31,231,31,126,31,126,30,220,31,106,31,113,31,8,31,111,31,111,30,111,29,177,31,217,31,91,31,157,31,74,31,236,31,236,30,99,31,147,31,147,30,195,31,195,30,195,29,195,28,244,31,2,31,162,31,140,31,169,31,169,30,223,31,119,31,119,30,75,31,7,31,41,31,65,31,185,31,246,31,246,30,47,31,102,31,102,30,102,29,140,31,217,31,173,31,44,31,254,31,130,31,101,31,5,31,90,31,61,31,147,31,147,30,148,31,142,31,142,30,208,31,3,31,3,30,96,31,237,31,102,31,91,31,4,31,4,30,4,29,4,28,4,27,73,31,87,31,194,31,61,31,61,30,39,31,39,30,56,31,56,30,88,31,59,31,110,31,102,31,142,31,187,31,181,31,34,31,34,30,34,29,210,31,210,30,210,29,210,28,119,31,119,30,252,31,212,31,212,30,212,29,92,31,100,31,255,31,157,31,128,31,128,30,227,31,87,31,42,31,98,31,118,31,153,31,40,31,33,31,249,31,223,31,234,31,244,31,237,31,29,31,67,31,67,30,104,31,26,31,228,31,203,31,192,31,227,31,227,30,101,31,101,30,101,29,157,31,85,31,157,31,158,31,168,31,251,31,47,31,63,31,148,31,104,31,182,31,54,31,54,30,251,31,174,31,177,31,88,31,88,30,214,31,214,30,102,31,47,31,221,31,163,31,133,31,192,31,203,31,118,31,70,31,70,30,143,31,62,31,62,30,207,31,175,31,47,31,126,31,126,30,21,31,150,31,247,31,91,31,109,31,192,31,25,31,25,30,104,31,60,31,136,31,139,31,89,31,105,31,43,31,43,30,137,31,27,31,20,31,20,30,208,31,206,31,228,31,228,30,237,31,55,31,73,31,73,30,68,31,68,30,88,31,197,31,78,31,107,31,211,31,196,31,117,31,231,31,16,31,162,31,139,31,139,30,221,31,221,30,17,31,117,31,80,31,211,31,225,31,162,31,162,30,154,31,154,30,84,31,178,31,72,31,96,31,12,31,144,31,223,31,246,31,157,31,58,31,140,31,218,31,118,31,118,30,118,29,118,28,68,31,90,31,55,31,126,31,117,31,9,31,191,31,250,31,172,31,212,31,212,30,116,31,154,31,38,31,38,30,38,29,107,31,182,31,182,30,201,31,201,30,174,31,174,30,174,29,185,31,166,31,196,31,107,31,220,31,64,31,216,31,10,31,20,31,4,31,4,30,170,31,170,30,36,31,228,31,110,31,234,31,109,31,109,30,211,31,224,31,174,31,228,31,181,31,181,30,126,31,109,31,223,31,223,30,223,29,223,28,60,31,84,31,149,31,2,31,28,31,240,31,240,30,211,31,82,31,41,31,247,31,77,31,101,31,156,31,156,30,196,31,196,30,196,29,196,28,22,31,223,31,13,31,13,30,13,29,14,31,97,31,97,30,239,31,239,30,239,29,25,31,218,31,191,31,191,30,191,29,34,31,27,31,124,31,98,31,206,31,82,31,34,31,182,31,19,31,97,31,199,31,130,31,74,31,199,31,33,31,33,30,16,31,171,31,171,30,171,29,171,28,150,31,150,30,188,31,144,31,144,30,118,31,219,31,126,31,165,31,165,30,180,31,105,31,195,31,196,31,249,31,152,31,124,31,124,30,57,31,57,30,103,31,123,31,123,30,63,31,82,31,82,30,32,31,4,31,4,30,43,31,24,31,71,31,71,30,172,31,107,31,107,30,214,31,18,31,18,30,43,31,74,31,228,31,22,31,208,31,16,31,107,31,9,31,9,30,101,31,114,31,202,31,58,31,58,30,28,31,85,31,115,31,251,31,212,31,194,31,107,31,95,31,95,30,48,31,48,30,15,31,65,31,100,31,100,30,94,31,8,31,198,31,209,31,209,30,49,31,157,31,241,31,241,30,24,31,184,31,191,31,175,31,18,31,18,30,64,31,173,31,236,31,200,31,243,31,41,31,41,30,192,31,168,31,120,31,133,31,133,30,178,31,191,31,105,31,191,31,34,31,223,31,223,30,223,29,47,31,47,30,253,31,8,31,104,31,49,31,110,31,110,30,70,31,104,31,138,31,193,31,196,31,196,30,20,31,109,31,172,31,158,31,8,31,245,31,128,31,227,31,93,31,17,31,83,31,83,30,83,29,240,31,75,31,57,31,95,31,170,31,195,31,79,31,99,31,99,30,193,31,193,30,83,31,179,31,11,31,213,31,103,31,125,31,90,31,2,31,68,31,139,31,127,31,245,31,100,31,100,30,83,31,30,31,157,31,197,31,124,31,194,31,156,31,85,31,152,31,173,31,233,31,233,30,255,31,255,30,91,31,247,31,247,30,240,31,237,31,189,31,37,31,159,31,159,30,241,31,74,31,116,31,96,31,140,31,203,31,19,31,105,31,253,31,153,31,153,30,234,31,231,31,202,31,248,31,111,31,111,30,111,29,111,28,130,31,1,31,104,31,216,31,216,30,183,31,183,30,28,31,119,31,67,31,106,31,75,31,161,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
