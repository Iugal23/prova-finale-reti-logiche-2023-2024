-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_458 is
end project_tb_458;

architecture project_tb_arch_458 of project_tb_458 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 968;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (103,0,85,0,0,0,189,0,0,0,74,0,177,0,152,0,224,0,66,0,244,0,41,0,147,0,218,0,96,0,236,0,166,0,51,0,61,0,0,0,0,0,0,0,69,0,25,0,49,0,234,0,108,0,207,0,106,0,129,0,251,0,199,0,0,0,2,0,0,0,190,0,132,0,0,0,182,0,82,0,46,0,83,0,121,0,128,0,131,0,100,0,49,0,21,0,107,0,0,0,186,0,103,0,110,0,35,0,52,0,60,0,177,0,189,0,240,0,249,0,7,0,195,0,0,0,54,0,207,0,0,0,85,0,135,0,184,0,174,0,0,0,5,0,116,0,0,0,0,0,84,0,210,0,164,0,200,0,186,0,15,0,0,0,140,0,154,0,156,0,0,0,247,0,117,0,137,0,179,0,99,0,0,0,59,0,251,0,35,0,44,0,0,0,131,0,0,0,0,0,135,0,20,0,200,0,212,0,111,0,4,0,176,0,56,0,144,0,73,0,0,0,181,0,225,0,239,0,214,0,96,0,73,0,14,0,90,0,132,0,200,0,213,0,0,0,0,0,208,0,30,0,6,0,0,0,120,0,0,0,77,0,251,0,73,0,70,0,74,0,25,0,58,0,47,0,0,0,0,0,41,0,0,0,218,0,59,0,32,0,130,0,0,0,149,0,0,0,56,0,139,0,44,0,14,0,29,0,152,0,91,0,131,0,29,0,0,0,185,0,0,0,7,0,65,0,189,0,153,0,97,0,0,0,70,0,116,0,161,0,0,0,22,0,3,0,255,0,90,0,0,0,160,0,48,0,0,0,124,0,139,0,94,0,159,0,0,0,135,0,243,0,61,0,0,0,93,0,128,0,0,0,0,0,0,0,24,0,181,0,0,0,88,0,225,0,243,0,117,0,154,0,62,0,42,0,196,0,201,0,0,0,0,0,0,0,0,0,7,0,199,0,135,0,185,0,153,0,14,0,235,0,15,0,0,0,112,0,56,0,255,0,76,0,0,0,45,0,54,0,238,0,0,0,75,0,170,0,158,0,217,0,0,0,164,0,0,0,227,0,131,0,82,0,207,0,196,0,228,0,0,0,68,0,252,0,187,0,125,0,125,0,0,0,127,0,34,0,248,0,168,0,86,0,0,0,0,0,0,0,35,0,181,0,95,0,7,0,240,0,134,0,172,0,204,0,0,0,79,0,135,0,169,0,0,0,137,0,52,0,61,0,99,0,215,0,242,0,0,0,197,0,65,0,0,0,66,0,33,0,230,0,41,0,63,0,172,0,0,0,104,0,51,0,227,0,248,0,101,0,196,0,118,0,0,0,93,0,125,0,201,0,57,0,137,0,180,0,124,0,95,0,192,0,200,0,226,0,212,0,61,0,0,0,215,0,176,0,19,0,0,0,0,0,49,0,184,0,245,0,11,0,167,0,187,0,0,0,152,0,86,0,170,0,250,0,226,0,226,0,0,0,115,0,74,0,47,0,0,0,108,0,39,0,226,0,107,0,0,0,171,0,236,0,211,0,0,0,212,0,0,0,161,0,140,0,221,0,245,0,183,0,152,0,101,0,0,0,0,0,251,0,28,0,38,0,182,0,29,0,170,0,0,0,75,0,45,0,183,0,177,0,32,0,114,0,231,0,41,0,83,0,111,0,99,0,250,0,0,0,118,0,128,0,80,0,169,0,231,0,169,0,0,0,120,0,150,0,40,0,215,0,84,0,254,0,0,0,183,0,90,0,236,0,226,0,0,0,11,0,106,0,158,0,43,0,0,0,54,0,32,0,124,0,65,0,78,0,22,0,0,0,210,0,11,0,141,0,35,0,0,0,23,0,150,0,114,0,91,0,17,0,0,0,47,0,153,0,0,0,225,0,193,0,72,0,80,0,22,0,0,0,0,0,255,0,171,0,109,0,252,0,0,0,202,0,71,0,0,0,211,0,37,0,106,0,44,0,0,0,218,0,184,0,49,0,35,0,96,0,72,0,190,0,49,0,0,0,0,0,0,0,186,0,38,0,4,0,23,0,213,0,234,0,0,0,40,0,212,0,91,0,30,0,144,0,33,0,0,0,53,0,104,0,35,0,16,0,162,0,254,0,168,0,0,0,153,0,190,0,97,0,200,0,0,0,233,0,92,0,3,0,0,0,174,0,108,0,66,0,0,0,1,0,20,0,221,0,255,0,0,0,4,0,55,0,139,0,0,0,144,0,14,0,246,0,0,0,186,0,11,0,0,0,207,0,0,0,203,0,79,0,82,0,203,0,134,0,176,0,20,0,229,0,107,0,166,0,32,0,192,0,0,0,51,0,243,0,5,0,156,0,0,0,179,0,92,0,142,0,85,0,2,0,0,0,178,0,137,0,0,0,55,0,210,0,212,0,170,0,102,0,0,0,7,0,121,0,223,0,9,0,212,0,80,0,218,0,19,0,83,0,0,0,58,0,200,0,172,0,169,0,70,0,56,0,85,0,74,0,158,0,72,0,0,0,157,0,85,0,117,0,111,0,0,0,54,0,0,0,80,0,214,0,173,0,0,0,218,0,230,0,184,0,248,0,0,0,149,0,0,0,131,0,64,0,223,0,44,0,50,0,42,0,146,0,0,0,239,0,0,0,76,0,178,0,61,0,243,0,0,0,255,0,0,0,55,0,78,0,0,0,164,0,220,0,144,0,185,0,125,0,0,0,191,0,123,0,239,0,169,0,0,0,69,0,210,0,93,0,117,0,85,0,0,0,173,0,63,0,196,0,26,0,16,0,0,0,134,0,227,0,245,0,215,0,0,0,47,0,217,0,137,0,173,0,0,0,33,0,140,0,164,0,93,0,0,0,192,0,143,0,58,0,77,0,0,0,246,0,154,0,94,0,184,0,146,0,96,0,0,0,13,0,155,0,22,0,44,0,65,0,107,0,218,0,3,0,143,0,80,0,233,0,72,0,243,0,79,0,0,0,111,0,143,0,0,0,30,0,19,0,215,0,228,0,209,0,100,0,217,0,18,0,99,0,116,0,35,0,0,0,0,0,157,0,96,0,171,0,4,0,126,0,123,0,122,0,158,0,255,0,0,0,71,0,24,0,105,0,0,0,101,0,0,0,199,0,130,0,137,0,233,0,225,0,91,0,193,0,0,0,77,0,189,0,0,0,87,0,28,0,150,0,0,0,55,0,132,0,137,0,16,0,0,0,176,0,221,0,50,0,0,0,0,0,152,0,48,0,0,0,187,0,32,0,147,0,182,0,113,0,0,0,133,0,184,0,118,0,243,0,133,0,114,0,83,0,0,0,44,0,0,0,178,0,74,0,149,0,83,0,114,0,164,0,0,0,156,0,84,0,195,0,248,0,62,0,210,0,243,0,37,0,65,0,251,0,0,0,0,0,0,0,147,0,18,0,0,0,136,0,157,0,19,0,57,0,126,0,135,0,175,0,227,0,86,0,165,0,0,0,11,0,0,0,161,0,0,0,165,0,110,0,68,0,52,0,200,0,0,0,205,0,220,0,206,0,0,0,23,0,137,0,117,0,208,0,105,0,128,0,209,0,61,0,214,0,15,0,255,0,245,0,221,0,123,0,80,0,250,0,229,0,19,0,62,0,12,0,203,0,62,0,90,0,170,0,236,0,0,0,0,0,0,0,7,0,206,0,29,0,0,0,157,0,0,0,140,0,161,0,213,0,0,0,241,0,254,0,190,0,56,0,215,0,142,0,206,0,162,0,15,0,100,0,10,0,216,0,1,0,7,0,0,0,76,0,116,0,205,0,48,0,109,0,0,0,0,0,0,0,0,0,232,0,0,0,29,0,161,0,35,0,237,0,108,0,180,0,247,0,0,0,233,0,233,0,195,0,0,0,91,0,53,0,40,0,138,0,239,0,210,0,199,0,224,0,113,0,19,0,0,0,19,0,239,0,130,0,18,0,39,0,101,0,192,0,169,0,145,0,152,0,107,0,10,0,0,0,174,0,54,0,100,0,50,0,113,0,0,0,53,0,40,0,89,0,145,0,242,0,0,0,114,0,0,0,142,0,0,0,0,0,140,0,58,0,232,0,9,0,0,0,0,0,209,0,233,0,179,0,0,0,163,0,18,0,222,0,21,0,214,0,29,0,95,0,24,0,202,0,220,0,156,0,86,0,150,0,92,0,224,0,151,0,0,0,57,0,0,0,220,0,187,0,80,0,108,0,115,0,195,0,25,0,211,0,82,0,221,0,65,0,0,0,0,0,54,0,135,0,31,0,222,0,10,0,152,0,229,0,47,0,104,0,0,0,107,0,215,0,53,0,169,0,233,0,205,0,82,0,254,0,229,0,0,0,142,0,23,0,40,0,125,0,139,0,3,0,0,0,24,0,0,0);
signal scenario_full  : scenario_type := (103,31,85,31,85,30,189,31,189,30,74,31,177,31,152,31,224,31,66,31,244,31,41,31,147,31,218,31,96,31,236,31,166,31,51,31,61,31,61,30,61,29,61,28,69,31,25,31,49,31,234,31,108,31,207,31,106,31,129,31,251,31,199,31,199,30,2,31,2,30,190,31,132,31,132,30,182,31,82,31,46,31,83,31,121,31,128,31,131,31,100,31,49,31,21,31,107,31,107,30,186,31,103,31,110,31,35,31,52,31,60,31,177,31,189,31,240,31,249,31,7,31,195,31,195,30,54,31,207,31,207,30,85,31,135,31,184,31,174,31,174,30,5,31,116,31,116,30,116,29,84,31,210,31,164,31,200,31,186,31,15,31,15,30,140,31,154,31,156,31,156,30,247,31,117,31,137,31,179,31,99,31,99,30,59,31,251,31,35,31,44,31,44,30,131,31,131,30,131,29,135,31,20,31,200,31,212,31,111,31,4,31,176,31,56,31,144,31,73,31,73,30,181,31,225,31,239,31,214,31,96,31,73,31,14,31,90,31,132,31,200,31,213,31,213,30,213,29,208,31,30,31,6,31,6,30,120,31,120,30,77,31,251,31,73,31,70,31,74,31,25,31,58,31,47,31,47,30,47,29,41,31,41,30,218,31,59,31,32,31,130,31,130,30,149,31,149,30,56,31,139,31,44,31,14,31,29,31,152,31,91,31,131,31,29,31,29,30,185,31,185,30,7,31,65,31,189,31,153,31,97,31,97,30,70,31,116,31,161,31,161,30,22,31,3,31,255,31,90,31,90,30,160,31,48,31,48,30,124,31,139,31,94,31,159,31,159,30,135,31,243,31,61,31,61,30,93,31,128,31,128,30,128,29,128,28,24,31,181,31,181,30,88,31,225,31,243,31,117,31,154,31,62,31,42,31,196,31,201,31,201,30,201,29,201,28,201,27,7,31,199,31,135,31,185,31,153,31,14,31,235,31,15,31,15,30,112,31,56,31,255,31,76,31,76,30,45,31,54,31,238,31,238,30,75,31,170,31,158,31,217,31,217,30,164,31,164,30,227,31,131,31,82,31,207,31,196,31,228,31,228,30,68,31,252,31,187,31,125,31,125,31,125,30,127,31,34,31,248,31,168,31,86,31,86,30,86,29,86,28,35,31,181,31,95,31,7,31,240,31,134,31,172,31,204,31,204,30,79,31,135,31,169,31,169,30,137,31,52,31,61,31,99,31,215,31,242,31,242,30,197,31,65,31,65,30,66,31,33,31,230,31,41,31,63,31,172,31,172,30,104,31,51,31,227,31,248,31,101,31,196,31,118,31,118,30,93,31,125,31,201,31,57,31,137,31,180,31,124,31,95,31,192,31,200,31,226,31,212,31,61,31,61,30,215,31,176,31,19,31,19,30,19,29,49,31,184,31,245,31,11,31,167,31,187,31,187,30,152,31,86,31,170,31,250,31,226,31,226,31,226,30,115,31,74,31,47,31,47,30,108,31,39,31,226,31,107,31,107,30,171,31,236,31,211,31,211,30,212,31,212,30,161,31,140,31,221,31,245,31,183,31,152,31,101,31,101,30,101,29,251,31,28,31,38,31,182,31,29,31,170,31,170,30,75,31,45,31,183,31,177,31,32,31,114,31,231,31,41,31,83,31,111,31,99,31,250,31,250,30,118,31,128,31,80,31,169,31,231,31,169,31,169,30,120,31,150,31,40,31,215,31,84,31,254,31,254,30,183,31,90,31,236,31,226,31,226,30,11,31,106,31,158,31,43,31,43,30,54,31,32,31,124,31,65,31,78,31,22,31,22,30,210,31,11,31,141,31,35,31,35,30,23,31,150,31,114,31,91,31,17,31,17,30,47,31,153,31,153,30,225,31,193,31,72,31,80,31,22,31,22,30,22,29,255,31,171,31,109,31,252,31,252,30,202,31,71,31,71,30,211,31,37,31,106,31,44,31,44,30,218,31,184,31,49,31,35,31,96,31,72,31,190,31,49,31,49,30,49,29,49,28,186,31,38,31,4,31,23,31,213,31,234,31,234,30,40,31,212,31,91,31,30,31,144,31,33,31,33,30,53,31,104,31,35,31,16,31,162,31,254,31,168,31,168,30,153,31,190,31,97,31,200,31,200,30,233,31,92,31,3,31,3,30,174,31,108,31,66,31,66,30,1,31,20,31,221,31,255,31,255,30,4,31,55,31,139,31,139,30,144,31,14,31,246,31,246,30,186,31,11,31,11,30,207,31,207,30,203,31,79,31,82,31,203,31,134,31,176,31,20,31,229,31,107,31,166,31,32,31,192,31,192,30,51,31,243,31,5,31,156,31,156,30,179,31,92,31,142,31,85,31,2,31,2,30,178,31,137,31,137,30,55,31,210,31,212,31,170,31,102,31,102,30,7,31,121,31,223,31,9,31,212,31,80,31,218,31,19,31,83,31,83,30,58,31,200,31,172,31,169,31,70,31,56,31,85,31,74,31,158,31,72,31,72,30,157,31,85,31,117,31,111,31,111,30,54,31,54,30,80,31,214,31,173,31,173,30,218,31,230,31,184,31,248,31,248,30,149,31,149,30,131,31,64,31,223,31,44,31,50,31,42,31,146,31,146,30,239,31,239,30,76,31,178,31,61,31,243,31,243,30,255,31,255,30,55,31,78,31,78,30,164,31,220,31,144,31,185,31,125,31,125,30,191,31,123,31,239,31,169,31,169,30,69,31,210,31,93,31,117,31,85,31,85,30,173,31,63,31,196,31,26,31,16,31,16,30,134,31,227,31,245,31,215,31,215,30,47,31,217,31,137,31,173,31,173,30,33,31,140,31,164,31,93,31,93,30,192,31,143,31,58,31,77,31,77,30,246,31,154,31,94,31,184,31,146,31,96,31,96,30,13,31,155,31,22,31,44,31,65,31,107,31,218,31,3,31,143,31,80,31,233,31,72,31,243,31,79,31,79,30,111,31,143,31,143,30,30,31,19,31,215,31,228,31,209,31,100,31,217,31,18,31,99,31,116,31,35,31,35,30,35,29,157,31,96,31,171,31,4,31,126,31,123,31,122,31,158,31,255,31,255,30,71,31,24,31,105,31,105,30,101,31,101,30,199,31,130,31,137,31,233,31,225,31,91,31,193,31,193,30,77,31,189,31,189,30,87,31,28,31,150,31,150,30,55,31,132,31,137,31,16,31,16,30,176,31,221,31,50,31,50,30,50,29,152,31,48,31,48,30,187,31,32,31,147,31,182,31,113,31,113,30,133,31,184,31,118,31,243,31,133,31,114,31,83,31,83,30,44,31,44,30,178,31,74,31,149,31,83,31,114,31,164,31,164,30,156,31,84,31,195,31,248,31,62,31,210,31,243,31,37,31,65,31,251,31,251,30,251,29,251,28,147,31,18,31,18,30,136,31,157,31,19,31,57,31,126,31,135,31,175,31,227,31,86,31,165,31,165,30,11,31,11,30,161,31,161,30,165,31,110,31,68,31,52,31,200,31,200,30,205,31,220,31,206,31,206,30,23,31,137,31,117,31,208,31,105,31,128,31,209,31,61,31,214,31,15,31,255,31,245,31,221,31,123,31,80,31,250,31,229,31,19,31,62,31,12,31,203,31,62,31,90,31,170,31,236,31,236,30,236,29,236,28,7,31,206,31,29,31,29,30,157,31,157,30,140,31,161,31,213,31,213,30,241,31,254,31,190,31,56,31,215,31,142,31,206,31,162,31,15,31,100,31,10,31,216,31,1,31,7,31,7,30,76,31,116,31,205,31,48,31,109,31,109,30,109,29,109,28,109,27,232,31,232,30,29,31,161,31,35,31,237,31,108,31,180,31,247,31,247,30,233,31,233,31,195,31,195,30,91,31,53,31,40,31,138,31,239,31,210,31,199,31,224,31,113,31,19,31,19,30,19,31,239,31,130,31,18,31,39,31,101,31,192,31,169,31,145,31,152,31,107,31,10,31,10,30,174,31,54,31,100,31,50,31,113,31,113,30,53,31,40,31,89,31,145,31,242,31,242,30,114,31,114,30,142,31,142,30,142,29,140,31,58,31,232,31,9,31,9,30,9,29,209,31,233,31,179,31,179,30,163,31,18,31,222,31,21,31,214,31,29,31,95,31,24,31,202,31,220,31,156,31,86,31,150,31,92,31,224,31,151,31,151,30,57,31,57,30,220,31,187,31,80,31,108,31,115,31,195,31,25,31,211,31,82,31,221,31,65,31,65,30,65,29,54,31,135,31,31,31,222,31,10,31,152,31,229,31,47,31,104,31,104,30,107,31,215,31,53,31,169,31,233,31,205,31,82,31,254,31,229,31,229,30,142,31,23,31,40,31,125,31,139,31,3,31,3,30,24,31,24,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
