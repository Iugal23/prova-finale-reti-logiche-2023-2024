-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 675;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (32,0,248,0,1,0,205,0,199,0,246,0,0,0,222,0,74,0,227,0,235,0,29,0,119,0,0,0,82,0,0,0,228,0,0,0,90,0,108,0,242,0,232,0,68,0,0,0,80,0,244,0,16,0,63,0,73,0,138,0,49,0,181,0,81,0,224,0,128,0,107,0,0,0,77,0,128,0,32,0,187,0,240,0,0,0,0,0,22,0,209,0,196,0,12,0,148,0,100,0,251,0,92,0,148,0,254,0,51,0,217,0,0,0,167,0,179,0,68,0,97,0,0,0,0,0,0,0,30,0,22,0,137,0,30,0,100,0,0,0,140,0,0,0,0,0,182,0,183,0,0,0,125,0,0,0,219,0,58,0,0,0,26,0,249,0,237,0,0,0,24,0,195,0,0,0,250,0,137,0,93,0,0,0,72,0,186,0,78,0,166,0,233,0,177,0,127,0,0,0,215,0,102,0,0,0,216,0,0,0,0,0,128,0,0,0,110,0,0,0,167,0,249,0,35,0,183,0,58,0,183,0,0,0,143,0,92,0,0,0,190,0,42,0,124,0,108,0,221,0,0,0,165,0,0,0,181,0,229,0,0,0,0,0,123,0,203,0,163,0,65,0,0,0,0,0,82,0,38,0,251,0,238,0,7,0,86,0,70,0,190,0,19,0,79,0,79,0,0,0,42,0,108,0,234,0,113,0,194,0,97,0,80,0,0,0,7,0,145,0,1,0,58,0,251,0,86,0,175,0,54,0,0,0,253,0,16,0,129,0,0,0,194,0,233,0,99,0,76,0,0,0,0,0,136,0,84,0,59,0,184,0,109,0,40,0,0,0,164,0,30,0,0,0,251,0,0,0,210,0,0,0,0,0,67,0,0,0,121,0,9,0,0,0,0,0,166,0,197,0,60,0,176,0,0,0,0,0,144,0,224,0,0,0,143,0,222,0,14,0,8,0,176,0,162,0,181,0,155,0,40,0,208,0,189,0,67,0,200,0,125,0,65,0,0,0,216,0,214,0,198,0,0,0,138,0,188,0,255,0,240,0,0,0,23,0,30,0,0,0,0,0,0,0,169,0,150,0,187,0,134,0,51,0,55,0,223,0,209,0,81,0,169,0,103,0,146,0,113,0,19,0,202,0,154,0,152,0,0,0,52,0,251,0,247,0,160,0,69,0,20,0,0,0,62,0,117,0,0,0,0,0,87,0,224,0,113,0,0,0,33,0,0,0,0,0,194,0,176,0,13,0,0,0,38,0,85,0,138,0,40,0,199,0,157,0,0,0,99,0,29,0,102,0,0,0,136,0,84,0,138,0,238,0,15,0,0,0,88,0,161,0,14,0,160,0,133,0,154,0,214,0,0,0,126,0,163,0,230,0,72,0,12,0,165,0,0,0,95,0,0,0,26,0,197,0,0,0,159,0,0,0,86,0,108,0,189,0,204,0,145,0,213,0,0,0,40,0,251,0,0,0,220,0,60,0,94,0,122,0,91,0,82,0,97,0,228,0,43,0,197,0,87,0,152,0,13,0,130,0,42,0,48,0,185,0,0,0,0,0,130,0,138,0,141,0,41,0,0,0,57,0,0,0,235,0,126,0,119,0,0,0,115,0,132,0,205,0,67,0,174,0,97,0,34,0,150,0,0,0,38,0,117,0,50,0,65,0,249,0,0,0,0,0,252,0,90,0,126,0,157,0,111,0,231,0,0,0,99,0,100,0,242,0,185,0,46,0,197,0,16,0,74,0,0,0,103,0,249,0,63,0,156,0,173,0,188,0,159,0,248,0,114,0,0,0,94,0,250,0,0,0,9,0,139,0,229,0,34,0,242,0,100,0,184,0,228,0,192,0,138,0,72,0,0,0,26,0,197,0,44,0,228,0,151,0,17,0,22,0,86,0,229,0,21,0,69,0,115,0,114,0,53,0,171,0,95,0,190,0,48,0,41,0,15,0,229,0,17,0,0,0,188,0,165,0,103,0,0,0,73,0,202,0,0,0,71,0,4,0,123,0,242,0,86,0,97,0,80,0,0,0,0,0,0,0,197,0,186,0,164,0,0,0,32,0,204,0,6,0,0,0,116,0,3,0,0,0,65,0,248,0,111,0,127,0,0,0,41,0,71,0,243,0,171,0,135,0,154,0,197,0,0,0,125,0,250,0,27,0,123,0,254,0,155,0,196,0,21,0,169,0,0,0,0,0,167,0,105,0,115,0,169,0,206,0,94,0,58,0,0,0,224,0,156,0,153,0,37,0,249,0,25,0,0,0,224,0,0,0,229,0,13,0,85,0,200,0,125,0,0,0,200,0,176,0,105,0,72,0,79,0,56,0,42,0,25,0,0,0,95,0,5,0,77,0,254,0,199,0,3,0,93,0,0,0,169,0,115,0,0,0,84,0,60,0,5,0,175,0,81,0,170,0,59,0,22,0,80,0,62,0,131,0,146,0,23,0,61,0,0,0,0,0,48,0,174,0,140,0,197,0,63,0,205,0,102,0,0,0,0,0,8,0,249,0,0,0,221,0,112,0,143,0,102,0,221,0,0,0,0,0,166,0,84,0,0,0,96,0,115,0,6,0,155,0,225,0,0,0,60,0,0,0,0,0,98,0,67,0,60,0,120,0,74,0,141,0,228,0,0,0,0,0,211,0,182,0,18,0,130,0,74,0,134,0,0,0,139,0,203,0,209,0,107,0,0,0,0,0,223,0,84,0,175,0,9,0,0,0,63,0,238,0,111,0,0,0,133,0,75,0,188,0,0,0,0,0,92,0,203,0,165,0,0,0,214,0,103,0,207,0,57,0,0,0,0,0,0,0,0,0,143,0,247,0,29,0,0,0,140,0,157,0,0,0,11,0,178,0,156,0,0,0,0,0,40,0,193,0,185,0,143,0,20,0,4,0,1,0,141,0,157,0,0,0,0,0,0,0,63,0,0,0,173,0,209,0,9,0,59,0,15,0,164,0,12,0,0,0,222,0,250,0,225,0,184,0,192,0,0,0,65,0,124,0,113,0,30,0,85,0,207,0,150,0,0,0,223,0);
signal scenario_full  : scenario_type := (32,31,248,31,1,31,205,31,199,31,246,31,246,30,222,31,74,31,227,31,235,31,29,31,119,31,119,30,82,31,82,30,228,31,228,30,90,31,108,31,242,31,232,31,68,31,68,30,80,31,244,31,16,31,63,31,73,31,138,31,49,31,181,31,81,31,224,31,128,31,107,31,107,30,77,31,128,31,32,31,187,31,240,31,240,30,240,29,22,31,209,31,196,31,12,31,148,31,100,31,251,31,92,31,148,31,254,31,51,31,217,31,217,30,167,31,179,31,68,31,97,31,97,30,97,29,97,28,30,31,22,31,137,31,30,31,100,31,100,30,140,31,140,30,140,29,182,31,183,31,183,30,125,31,125,30,219,31,58,31,58,30,26,31,249,31,237,31,237,30,24,31,195,31,195,30,250,31,137,31,93,31,93,30,72,31,186,31,78,31,166,31,233,31,177,31,127,31,127,30,215,31,102,31,102,30,216,31,216,30,216,29,128,31,128,30,110,31,110,30,167,31,249,31,35,31,183,31,58,31,183,31,183,30,143,31,92,31,92,30,190,31,42,31,124,31,108,31,221,31,221,30,165,31,165,30,181,31,229,31,229,30,229,29,123,31,203,31,163,31,65,31,65,30,65,29,82,31,38,31,251,31,238,31,7,31,86,31,70,31,190,31,19,31,79,31,79,31,79,30,42,31,108,31,234,31,113,31,194,31,97,31,80,31,80,30,7,31,145,31,1,31,58,31,251,31,86,31,175,31,54,31,54,30,253,31,16,31,129,31,129,30,194,31,233,31,99,31,76,31,76,30,76,29,136,31,84,31,59,31,184,31,109,31,40,31,40,30,164,31,30,31,30,30,251,31,251,30,210,31,210,30,210,29,67,31,67,30,121,31,9,31,9,30,9,29,166,31,197,31,60,31,176,31,176,30,176,29,144,31,224,31,224,30,143,31,222,31,14,31,8,31,176,31,162,31,181,31,155,31,40,31,208,31,189,31,67,31,200,31,125,31,65,31,65,30,216,31,214,31,198,31,198,30,138,31,188,31,255,31,240,31,240,30,23,31,30,31,30,30,30,29,30,28,169,31,150,31,187,31,134,31,51,31,55,31,223,31,209,31,81,31,169,31,103,31,146,31,113,31,19,31,202,31,154,31,152,31,152,30,52,31,251,31,247,31,160,31,69,31,20,31,20,30,62,31,117,31,117,30,117,29,87,31,224,31,113,31,113,30,33,31,33,30,33,29,194,31,176,31,13,31,13,30,38,31,85,31,138,31,40,31,199,31,157,31,157,30,99,31,29,31,102,31,102,30,136,31,84,31,138,31,238,31,15,31,15,30,88,31,161,31,14,31,160,31,133,31,154,31,214,31,214,30,126,31,163,31,230,31,72,31,12,31,165,31,165,30,95,31,95,30,26,31,197,31,197,30,159,31,159,30,86,31,108,31,189,31,204,31,145,31,213,31,213,30,40,31,251,31,251,30,220,31,60,31,94,31,122,31,91,31,82,31,97,31,228,31,43,31,197,31,87,31,152,31,13,31,130,31,42,31,48,31,185,31,185,30,185,29,130,31,138,31,141,31,41,31,41,30,57,31,57,30,235,31,126,31,119,31,119,30,115,31,132,31,205,31,67,31,174,31,97,31,34,31,150,31,150,30,38,31,117,31,50,31,65,31,249,31,249,30,249,29,252,31,90,31,126,31,157,31,111,31,231,31,231,30,99,31,100,31,242,31,185,31,46,31,197,31,16,31,74,31,74,30,103,31,249,31,63,31,156,31,173,31,188,31,159,31,248,31,114,31,114,30,94,31,250,31,250,30,9,31,139,31,229,31,34,31,242,31,100,31,184,31,228,31,192,31,138,31,72,31,72,30,26,31,197,31,44,31,228,31,151,31,17,31,22,31,86,31,229,31,21,31,69,31,115,31,114,31,53,31,171,31,95,31,190,31,48,31,41,31,15,31,229,31,17,31,17,30,188,31,165,31,103,31,103,30,73,31,202,31,202,30,71,31,4,31,123,31,242,31,86,31,97,31,80,31,80,30,80,29,80,28,197,31,186,31,164,31,164,30,32,31,204,31,6,31,6,30,116,31,3,31,3,30,65,31,248,31,111,31,127,31,127,30,41,31,71,31,243,31,171,31,135,31,154,31,197,31,197,30,125,31,250,31,27,31,123,31,254,31,155,31,196,31,21,31,169,31,169,30,169,29,167,31,105,31,115,31,169,31,206,31,94,31,58,31,58,30,224,31,156,31,153,31,37,31,249,31,25,31,25,30,224,31,224,30,229,31,13,31,85,31,200,31,125,31,125,30,200,31,176,31,105,31,72,31,79,31,56,31,42,31,25,31,25,30,95,31,5,31,77,31,254,31,199,31,3,31,93,31,93,30,169,31,115,31,115,30,84,31,60,31,5,31,175,31,81,31,170,31,59,31,22,31,80,31,62,31,131,31,146,31,23,31,61,31,61,30,61,29,48,31,174,31,140,31,197,31,63,31,205,31,102,31,102,30,102,29,8,31,249,31,249,30,221,31,112,31,143,31,102,31,221,31,221,30,221,29,166,31,84,31,84,30,96,31,115,31,6,31,155,31,225,31,225,30,60,31,60,30,60,29,98,31,67,31,60,31,120,31,74,31,141,31,228,31,228,30,228,29,211,31,182,31,18,31,130,31,74,31,134,31,134,30,139,31,203,31,209,31,107,31,107,30,107,29,223,31,84,31,175,31,9,31,9,30,63,31,238,31,111,31,111,30,133,31,75,31,188,31,188,30,188,29,92,31,203,31,165,31,165,30,214,31,103,31,207,31,57,31,57,30,57,29,57,28,57,27,143,31,247,31,29,31,29,30,140,31,157,31,157,30,11,31,178,31,156,31,156,30,156,29,40,31,193,31,185,31,143,31,20,31,4,31,1,31,141,31,157,31,157,30,157,29,157,28,63,31,63,30,173,31,209,31,9,31,59,31,15,31,164,31,12,31,12,30,222,31,250,31,225,31,184,31,192,31,192,30,65,31,124,31,113,31,30,31,85,31,207,31,150,31,150,30,223,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
