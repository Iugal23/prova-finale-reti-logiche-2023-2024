-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_106 is
end project_tb_106;

architecture project_tb_arch_106 of project_tb_106 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 830;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (121,0,159,0,0,0,239,0,6,0,26,0,48,0,44,0,244,0,214,0,192,0,0,0,11,0,24,0,144,0,28,0,37,0,132,0,183,0,157,0,75,0,217,0,136,0,107,0,102,0,92,0,153,0,0,0,0,0,28,0,83,0,9,0,0,0,127,0,167,0,191,0,19,0,201,0,140,0,0,0,112,0,228,0,159,0,244,0,0,0,0,0,52,0,190,0,161,0,0,0,34,0,0,0,168,0,0,0,181,0,76,0,45,0,169,0,27,0,85,0,229,0,129,0,120,0,0,0,214,0,126,0,106,0,48,0,114,0,206,0,0,0,59,0,148,0,0,0,0,0,93,0,91,0,70,0,54,0,55,0,0,0,28,0,40,0,15,0,0,0,46,0,15,0,99,0,0,0,84,0,0,0,216,0,64,0,142,0,247,0,140,0,169,0,40,0,0,0,16,0,227,0,221,0,226,0,36,0,19,0,88,0,161,0,163,0,0,0,108,0,97,0,0,0,0,0,168,0,175,0,101,0,0,0,17,0,244,0,105,0,20,0,0,0,139,0,172,0,189,0,61,0,100,0,67,0,0,0,0,0,0,0,122,0,233,0,0,0,0,0,16,0,0,0,0,0,22,0,209,0,0,0,17,0,0,0,0,0,203,0,215,0,190,0,153,0,116,0,129,0,0,0,0,0,174,0,181,0,0,0,41,0,163,0,64,0,4,0,229,0,225,0,0,0,155,0,0,0,108,0,36,0,160,0,0,0,199,0,0,0,0,0,0,0,0,0,201,0,12,0,0,0,52,0,150,0,91,0,205,0,166,0,21,0,0,0,59,0,181,0,123,0,20,0,154,0,0,0,133,0,0,0,170,0,38,0,189,0,0,0,0,0,114,0,0,0,9,0,101,0,0,0,254,0,195,0,128,0,217,0,235,0,0,0,98,0,65,0,0,0,20,0,0,0,211,0,236,0,0,0,8,0,0,0,0,0,172,0,0,0,0,0,155,0,143,0,91,0,14,0,0,0,177,0,38,0,196,0,0,0,0,0,0,0,0,0,14,0,94,0,23,0,156,0,167,0,207,0,22,0,27,0,29,0,172,0,113,0,164,0,0,0,168,0,178,0,91,0,224,0,212,0,0,0,41,0,216,0,0,0,159,0,54,0,238,0,50,0,9,0,30,0,113,0,95,0,234,0,133,0,216,0,56,0,0,0,76,0,66,0,212,0,153,0,85,0,64,0,159,0,55,0,163,0,0,0,20,0,168,0,100,0,199,0,185,0,222,0,154,0,247,0,215,0,0,0,95,0,229,0,0,0,151,0,0,0,148,0,53,0,191,0,83,0,155,0,0,0,212,0,154,0,87,0,0,0,0,0,142,0,218,0,203,0,144,0,248,0,7,0,0,0,73,0,210,0,195,0,0,0,119,0,250,0,0,0,0,0,0,0,171,0,16,0,0,0,185,0,47,0,232,0,0,0,15,0,111,0,8,0,48,0,0,0,143,0,231,0,18,0,31,0,0,0,22,0,40,0,89,0,216,0,127,0,0,0,194,0,171,0,67,0,65,0,35,0,115,0,0,0,42,0,5,0,109,0,205,0,133,0,166,0,99,0,17,0,156,0,13,0,205,0,178,0,0,0,0,0,120,0,47,0,0,0,122,0,0,0,234,0,0,0,99,0,0,0,100,0,16,0,106,0,54,0,202,0,111,0,163,0,116,0,73,0,25,0,119,0,140,0,178,0,0,0,100,0,233,0,106,0,120,0,0,0,48,0,115,0,85,0,60,0,193,0,208,0,69,0,123,0,178,0,0,0,84,0,171,0,112,0,0,0,202,0,0,0,52,0,170,0,97,0,36,0,0,0,38,0,34,0,151,0,28,0,0,0,14,0,33,0,49,0,68,0,0,0,0,0,0,0,0,0,0,0,115,0,3,0,71,0,0,0,178,0,84,0,97,0,79,0,241,0,18,0,0,0,79,0,24,0,0,0,113,0,34,0,0,0,144,0,0,0,224,0,11,0,4,0,0,0,0,0,155,0,138,0,185,0,60,0,6,0,177,0,218,0,10,0,98,0,139,0,45,0,34,0,0,0,252,0,157,0,187,0,132,0,25,0,86,0,0,0,189,0,0,0,0,0,136,0,189,0,0,0,111,0,158,0,118,0,11,0,232,0,224,0,66,0,0,0,227,0,211,0,3,0,126,0,195,0,184,0,0,0,81,0,183,0,0,0,206,0,156,0,2,0,206,0,234,0,68,0,105,0,126,0,102,0,183,0,218,0,57,0,209,0,70,0,255,0,54,0,4,0,151,0,8,0,0,0,0,0,23,0,0,0,208,0,172,0,0,0,72,0,53,0,0,0,71,0,97,0,0,0,165,0,128,0,154,0,57,0,38,0,194,0,107,0,0,0,136,0,144,0,95,0,141,0,155,0,30,0,160,0,124,0,0,0,148,0,53,0,70,0,0,0,227,0,28,0,77,0,156,0,217,0,141,0,255,0,0,0,1,0,124,0,220,0,0,0,138,0,239,0,111,0,81,0,150,0,0,0,55,0,229,0,154,0,29,0,29,0,37,0,6,0,71,0,0,0,15,0,105,0,169,0,108,0,245,0,72,0,27,0,82,0,23,0,156,0,0,0,116,0,0,0,247,0,59,0,17,0,211,0,229,0,169,0,184,0,0,0,206,0,85,0,0,0,0,0,0,0,156,0,0,0,185,0,178,0,119,0,0,0,149,0,68,0,102,0,233,0,171,0,169,0,130,0,136,0,85,0,160,0,0,0,42,0,254,0,83,0,174,0,44,0,0,0,116,0,0,0,219,0,63,0,236,0,22,0,0,0,47,0,0,0,0,0,93,0,94,0,201,0,14,0,194,0,161,0,183,0,242,0,43,0,249,0,128,0,238,0,220,0,18,0,7,0,48,0,79,0,0,0,0,0,185,0,166,0,0,0,31,0,154,0,0,0,74,0,211,0,170,0,35,0,0,0,0,0,0,0,37,0,0,0,0,0,120,0,225,0,61,0,174,0,82,0,11,0,149,0,143,0,97,0,146,0,228,0,141,0,146,0,146,0,97,0,0,0,247,0,0,0,0,0,0,0,0,0,182,0,174,0,27,0,65,0,28,0,217,0,247,0,0,0,0,0,228,0,2,0,202,0,199,0,226,0,51,0,64,0,26,0,141,0,12,0,197,0,243,0,81,0,0,0,102,0,21,0,114,0,137,0,18,0,0,0,0,0,150,0,170,0,0,0,165,0,243,0,165,0,79,0,174,0,19,0,129,0,152,0,24,0,75,0,0,0,170,0,0,0,126,0,11,0,101,0,193,0,0,0,61,0,207,0,81,0,192,0,77,0,226,0,0,0,192,0,222,0,52,0,127,0,172,0,243,0,87,0,0,0,63,0,208,0,0,0,13,0,110,0,200,0,188,0,220,0,93,0,139,0,136,0,0,0,87,0,51,0,239,0,90,0,10,0,191,0,192,0,131,0,106,0,223,0,238,0,211,0,61,0,221,0,89,0,208,0,0,0,134,0,11,0,154,0,103,0,13,0,205,0,112,0,163,0,178,0,203,0,0,0,102,0,233,0,22,0,16,0,112,0,87,0,91,0,39,0,72,0,160,0,109,0,0,0,0,0,219,0,217,0,29,0,107,0,128,0,176,0,0,0,255,0,0,0,183,0,239,0,190,0,4,0,163,0,117,0,254,0,211,0,249,0,239,0,0,0,129,0);
signal scenario_full  : scenario_type := (121,31,159,31,159,30,239,31,6,31,26,31,48,31,44,31,244,31,214,31,192,31,192,30,11,31,24,31,144,31,28,31,37,31,132,31,183,31,157,31,75,31,217,31,136,31,107,31,102,31,92,31,153,31,153,30,153,29,28,31,83,31,9,31,9,30,127,31,167,31,191,31,19,31,201,31,140,31,140,30,112,31,228,31,159,31,244,31,244,30,244,29,52,31,190,31,161,31,161,30,34,31,34,30,168,31,168,30,181,31,76,31,45,31,169,31,27,31,85,31,229,31,129,31,120,31,120,30,214,31,126,31,106,31,48,31,114,31,206,31,206,30,59,31,148,31,148,30,148,29,93,31,91,31,70,31,54,31,55,31,55,30,28,31,40,31,15,31,15,30,46,31,15,31,99,31,99,30,84,31,84,30,216,31,64,31,142,31,247,31,140,31,169,31,40,31,40,30,16,31,227,31,221,31,226,31,36,31,19,31,88,31,161,31,163,31,163,30,108,31,97,31,97,30,97,29,168,31,175,31,101,31,101,30,17,31,244,31,105,31,20,31,20,30,139,31,172,31,189,31,61,31,100,31,67,31,67,30,67,29,67,28,122,31,233,31,233,30,233,29,16,31,16,30,16,29,22,31,209,31,209,30,17,31,17,30,17,29,203,31,215,31,190,31,153,31,116,31,129,31,129,30,129,29,174,31,181,31,181,30,41,31,163,31,64,31,4,31,229,31,225,31,225,30,155,31,155,30,108,31,36,31,160,31,160,30,199,31,199,30,199,29,199,28,199,27,201,31,12,31,12,30,52,31,150,31,91,31,205,31,166,31,21,31,21,30,59,31,181,31,123,31,20,31,154,31,154,30,133,31,133,30,170,31,38,31,189,31,189,30,189,29,114,31,114,30,9,31,101,31,101,30,254,31,195,31,128,31,217,31,235,31,235,30,98,31,65,31,65,30,20,31,20,30,211,31,236,31,236,30,8,31,8,30,8,29,172,31,172,30,172,29,155,31,143,31,91,31,14,31,14,30,177,31,38,31,196,31,196,30,196,29,196,28,196,27,14,31,94,31,23,31,156,31,167,31,207,31,22,31,27,31,29,31,172,31,113,31,164,31,164,30,168,31,178,31,91,31,224,31,212,31,212,30,41,31,216,31,216,30,159,31,54,31,238,31,50,31,9,31,30,31,113,31,95,31,234,31,133,31,216,31,56,31,56,30,76,31,66,31,212,31,153,31,85,31,64,31,159,31,55,31,163,31,163,30,20,31,168,31,100,31,199,31,185,31,222,31,154,31,247,31,215,31,215,30,95,31,229,31,229,30,151,31,151,30,148,31,53,31,191,31,83,31,155,31,155,30,212,31,154,31,87,31,87,30,87,29,142,31,218,31,203,31,144,31,248,31,7,31,7,30,73,31,210,31,195,31,195,30,119,31,250,31,250,30,250,29,250,28,171,31,16,31,16,30,185,31,47,31,232,31,232,30,15,31,111,31,8,31,48,31,48,30,143,31,231,31,18,31,31,31,31,30,22,31,40,31,89,31,216,31,127,31,127,30,194,31,171,31,67,31,65,31,35,31,115,31,115,30,42,31,5,31,109,31,205,31,133,31,166,31,99,31,17,31,156,31,13,31,205,31,178,31,178,30,178,29,120,31,47,31,47,30,122,31,122,30,234,31,234,30,99,31,99,30,100,31,16,31,106,31,54,31,202,31,111,31,163,31,116,31,73,31,25,31,119,31,140,31,178,31,178,30,100,31,233,31,106,31,120,31,120,30,48,31,115,31,85,31,60,31,193,31,208,31,69,31,123,31,178,31,178,30,84,31,171,31,112,31,112,30,202,31,202,30,52,31,170,31,97,31,36,31,36,30,38,31,34,31,151,31,28,31,28,30,14,31,33,31,49,31,68,31,68,30,68,29,68,28,68,27,68,26,115,31,3,31,71,31,71,30,178,31,84,31,97,31,79,31,241,31,18,31,18,30,79,31,24,31,24,30,113,31,34,31,34,30,144,31,144,30,224,31,11,31,4,31,4,30,4,29,155,31,138,31,185,31,60,31,6,31,177,31,218,31,10,31,98,31,139,31,45,31,34,31,34,30,252,31,157,31,187,31,132,31,25,31,86,31,86,30,189,31,189,30,189,29,136,31,189,31,189,30,111,31,158,31,118,31,11,31,232,31,224,31,66,31,66,30,227,31,211,31,3,31,126,31,195,31,184,31,184,30,81,31,183,31,183,30,206,31,156,31,2,31,206,31,234,31,68,31,105,31,126,31,102,31,183,31,218,31,57,31,209,31,70,31,255,31,54,31,4,31,151,31,8,31,8,30,8,29,23,31,23,30,208,31,172,31,172,30,72,31,53,31,53,30,71,31,97,31,97,30,165,31,128,31,154,31,57,31,38,31,194,31,107,31,107,30,136,31,144,31,95,31,141,31,155,31,30,31,160,31,124,31,124,30,148,31,53,31,70,31,70,30,227,31,28,31,77,31,156,31,217,31,141,31,255,31,255,30,1,31,124,31,220,31,220,30,138,31,239,31,111,31,81,31,150,31,150,30,55,31,229,31,154,31,29,31,29,31,37,31,6,31,71,31,71,30,15,31,105,31,169,31,108,31,245,31,72,31,27,31,82,31,23,31,156,31,156,30,116,31,116,30,247,31,59,31,17,31,211,31,229,31,169,31,184,31,184,30,206,31,85,31,85,30,85,29,85,28,156,31,156,30,185,31,178,31,119,31,119,30,149,31,68,31,102,31,233,31,171,31,169,31,130,31,136,31,85,31,160,31,160,30,42,31,254,31,83,31,174,31,44,31,44,30,116,31,116,30,219,31,63,31,236,31,22,31,22,30,47,31,47,30,47,29,93,31,94,31,201,31,14,31,194,31,161,31,183,31,242,31,43,31,249,31,128,31,238,31,220,31,18,31,7,31,48,31,79,31,79,30,79,29,185,31,166,31,166,30,31,31,154,31,154,30,74,31,211,31,170,31,35,31,35,30,35,29,35,28,37,31,37,30,37,29,120,31,225,31,61,31,174,31,82,31,11,31,149,31,143,31,97,31,146,31,228,31,141,31,146,31,146,31,97,31,97,30,247,31,247,30,247,29,247,28,247,27,182,31,174,31,27,31,65,31,28,31,217,31,247,31,247,30,247,29,228,31,2,31,202,31,199,31,226,31,51,31,64,31,26,31,141,31,12,31,197,31,243,31,81,31,81,30,102,31,21,31,114,31,137,31,18,31,18,30,18,29,150,31,170,31,170,30,165,31,243,31,165,31,79,31,174,31,19,31,129,31,152,31,24,31,75,31,75,30,170,31,170,30,126,31,11,31,101,31,193,31,193,30,61,31,207,31,81,31,192,31,77,31,226,31,226,30,192,31,222,31,52,31,127,31,172,31,243,31,87,31,87,30,63,31,208,31,208,30,13,31,110,31,200,31,188,31,220,31,93,31,139,31,136,31,136,30,87,31,51,31,239,31,90,31,10,31,191,31,192,31,131,31,106,31,223,31,238,31,211,31,61,31,221,31,89,31,208,31,208,30,134,31,11,31,154,31,103,31,13,31,205,31,112,31,163,31,178,31,203,31,203,30,102,31,233,31,22,31,16,31,112,31,87,31,91,31,39,31,72,31,160,31,109,31,109,30,109,29,219,31,217,31,29,31,107,31,128,31,176,31,176,30,255,31,255,30,183,31,239,31,190,31,4,31,163,31,117,31,254,31,211,31,249,31,239,31,239,30,129,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
