-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_707 is
end project_tb_707;

architecture project_tb_arch_707 of project_tb_707 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 924;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (6,0,2,0,0,0,214,0,203,0,72,0,144,0,140,0,160,0,29,0,51,0,137,0,248,0,231,0,250,0,65,0,0,0,0,0,0,0,212,0,38,0,211,0,162,0,158,0,162,0,88,0,74,0,209,0,43,0,175,0,204,0,158,0,216,0,23,0,26,0,96,0,4,0,222,0,158,0,238,0,0,0,170,0,108,0,15,0,85,0,161,0,159,0,237,0,223,0,239,0,0,0,253,0,50,0,101,0,213,0,0,0,70,0,252,0,240,0,69,0,66,0,245,0,179,0,193,0,228,0,96,0,232,0,0,0,20,0,153,0,176,0,67,0,0,0,166,0,214,0,140,0,157,0,0,0,121,0,0,0,0,0,9,0,115,0,25,0,194,0,84,0,222,0,123,0,0,0,149,0,100,0,0,0,0,0,63,0,30,0,80,0,0,0,166,0,19,0,10,0,132,0,206,0,217,0,0,0,0,0,194,0,145,0,58,0,124,0,178,0,117,0,0,0,249,0,0,0,0,0,150,0,0,0,0,0,79,0,51,0,157,0,0,0,0,0,197,0,0,0,253,0,0,0,184,0,33,0,0,0,0,0,93,0,138,0,232,0,185,0,131,0,243,0,234,0,241,0,38,0,227,0,116,0,227,0,208,0,251,0,80,0,0,0,0,0,44,0,157,0,150,0,2,0,230,0,137,0,92,0,218,0,178,0,227,0,252,0,143,0,186,0,0,0,105,0,188,0,67,0,0,0,164,0,0,0,128,0,223,0,113,0,102,0,115,0,210,0,0,0,224,0,172,0,156,0,38,0,0,0,125,0,100,0,236,0,188,0,149,0,224,0,150,0,194,0,225,0,85,0,48,0,98,0,217,0,0,0,69,0,28,0,219,0,62,0,0,0,25,0,235,0,17,0,210,0,189,0,136,0,198,0,0,0,204,0,140,0,161,0,0,0,201,0,61,0,231,0,90,0,0,0,200,0,2,0,0,0,184,0,0,0,223,0,61,0,232,0,37,0,138,0,12,0,222,0,235,0,161,0,0,0,61,0,75,0,0,0,180,0,0,0,17,0,0,0,0,0,147,0,0,0,134,0,115,0,83,0,133,0,203,0,221,0,96,0,26,0,160,0,46,0,31,0,0,0,1,0,249,0,255,0,16,0,0,0,159,0,114,0,165,0,161,0,208,0,35,0,55,0,165,0,36,0,0,0,173,0,30,0,7,0,0,0,81,0,0,0,154,0,131,0,132,0,101,0,12,0,0,0,104,0,0,0,0,0,0,0,0,0,41,0,213,0,136,0,59,0,246,0,186,0,252,0,228,0,4,0,185,0,169,0,0,0,149,0,24,0,0,0,165,0,52,0,0,0,216,0,45,0,201,0,253,0,2,0,0,0,0,0,98,0,0,0,9,0,0,0,0,0,0,0,149,0,179,0,166,0,173,0,34,0,0,0,0,0,87,0,0,0,45,0,216,0,138,0,114,0,193,0,0,0,197,0,0,0,199,0,82,0,58,0,42,0,69,0,31,0,169,0,179,0,0,0,221,0,166,0,243,0,38,0,0,0,38,0,29,0,79,0,128,0,251,0,149,0,129,0,95,0,247,0,21,0,42,0,74,0,38,0,180,0,245,0,0,0,0,0,108,0,91,0,136,0,21,0,229,0,184,0,167,0,231,0,0,0,163,0,255,0,0,0,0,0,99,0,0,0,60,0,58,0,59,0,222,0,129,0,163,0,0,0,76,0,191,0,226,0,139,0,140,0,0,0,182,0,0,0,0,0,0,0,0,0,6,0,99,0,212,0,255,0,62,0,169,0,140,0,0,0,56,0,0,0,139,0,10,0,118,0,76,0,81,0,15,0,147,0,195,0,71,0,0,0,28,0,218,0,0,0,244,0,68,0,189,0,229,0,0,0,36,0,158,0,39,0,175,0,224,0,57,0,156,0,236,0,234,0,135,0,6,0,0,0,203,0,64,0,230,0,0,0,97,0,217,0,106,0,0,0,85,0,0,0,125,0,118,0,0,0,197,0,125,0,21,0,164,0,133,0,11,0,41,0,90,0,211,0,10,0,0,0,190,0,0,0,0,0,82,0,101,0,5,0,158,0,48,0,218,0,0,0,188,0,49,0,0,0,255,0,54,0,243,0,150,0,16,0,74,0,0,0,247,0,211,0,152,0,0,0,94,0,80,0,0,0,243,0,2,0,0,0,118,0,58,0,242,0,115,0,175,0,9,0,19,0,75,0,176,0,208,0,231,0,0,0,0,0,0,0,220,0,69,0,74,0,230,0,68,0,34,0,0,0,246,0,0,0,185,0,0,0,0,0,228,0,230,0,88,0,93,0,61,0,144,0,0,0,60,0,0,0,239,0,0,0,207,0,0,0,209,0,89,0,210,0,0,0,0,0,0,0,121,0,156,0,0,0,58,0,139,0,202,0,219,0,131,0,17,0,72,0,121,0,0,0,153,0,68,0,105,0,240,0,188,0,224,0,0,0,204,0,224,0,204,0,206,0,143,0,0,0,39,0,86,0,0,0,0,0,0,0,21,0,248,0,246,0,137,0,0,0,58,0,28,0,241,0,40,0,161,0,0,0,4,0,105,0,18,0,48,0,0,0,145,0,76,0,72,0,122,0,35,0,230,0,68,0,130,0,162,0,174,0,240,0,126,0,24,0,36,0,105,0,181,0,145,0,35,0,226,0,37,0,198,0,0,0,42,0,160,0,217,0,9,0,70,0,8,0,44,0,143,0,75,0,0,0,40,0,212,0,65,0,181,0,155,0,149,0,89,0,184,0,1,0,64,0,214,0,0,0,158,0,162,0,0,0,0,0,126,0,70,0,80,0,186,0,92,0,188,0,0,0,232,0,0,0,0,0,69,0,142,0,0,0,0,0,134,0,187,0,0,0,27,0,225,0,7,0,221,0,191,0,35,0,95,0,149,0,72,0,103,0,222,0,134,0,105,0,0,0,0,0,0,0,101,0,68,0,207,0,196,0,181,0,179,0,215,0,68,0,0,0,0,0,187,0,197,0,20,0,0,0,247,0,12,0,187,0,213,0,15,0,89,0,0,0,0,0,0,0,89,0,64,0,0,0,99,0,173,0,93,0,251,0,64,0,6,0,220,0,168,0,0,0,226,0,155,0,233,0,220,0,0,0,91,0,167,0,34,0,0,0,198,0,101,0,0,0,177,0,0,0,117,0,0,0,217,0,139,0,48,0,210,0,158,0,254,0,160,0,0,0,227,0,0,0,220,0,232,0,42,0,70,0,185,0,183,0,0,0,105,0,174,0,0,0,35,0,33,0,125,0,13,0,46,0,178,0,157,0,58,0,128,0,0,0,251,0,26,0,138,0,56,0,12,0,35,0,11,0,204,0,103,0,246,0,58,0,96,0,82,0,17,0,209,0,96,0,0,0,68,0,219,0,232,0,31,0,219,0,80,0,35,0,0,0,253,0,85,0,175,0,230,0,242,0,247,0,182,0,0,0,170,0,127,0,231,0,201,0,193,0,243,0,15,0,191,0,228,0,249,0,105,0,0,0,40,0,190,0,69,0,113,0,0,0,99,0,24,0,66,0,217,0,16,0,19,0,86,0,139,0,247,0,140,0,0,0,130,0,123,0,72,0,236,0,0,0,210,0,156,0,0,0,137,0,136,0,74,0,152,0,77,0,161,0,181,0,106,0,189,0,0,0,82,0,128,0,109,0,226,0,0,0,204,0,43,0,25,0,195,0,167,0,239,0,129,0,107,0,46,0,230,0,132,0,59,0,90,0,217,0,64,0,0,0,153,0,6,0,0,0,35,0,195,0,130,0,38,0,182,0,207,0,232,0,112,0,38,0,48,0,89,0,143,0,0,0,110,0,225,0,217,0,138,0,10,0,191,0,99,0,111,0,8,0,60,0,60,0,92,0,98,0,81,0,175,0,132,0,79,0,58,0,232,0,224,0,27,0,221,0,0,0,32,0,0,0,139,0,70,0,88,0,86,0,140,0,0,0,19,0,39,0,232,0,178,0,236,0,98,0,0,0,212,0,14,0,24,0,25,0,213,0,21,0,63,0,185,0,0,0,169,0,197,0,129,0,159,0,124,0,0,0,0,0,99,0,209,0,250,0,174,0,161,0,150,0,0,0,202,0,0,0,249,0);
signal scenario_full  : scenario_type := (6,31,2,31,2,30,214,31,203,31,72,31,144,31,140,31,160,31,29,31,51,31,137,31,248,31,231,31,250,31,65,31,65,30,65,29,65,28,212,31,38,31,211,31,162,31,158,31,162,31,88,31,74,31,209,31,43,31,175,31,204,31,158,31,216,31,23,31,26,31,96,31,4,31,222,31,158,31,238,31,238,30,170,31,108,31,15,31,85,31,161,31,159,31,237,31,223,31,239,31,239,30,253,31,50,31,101,31,213,31,213,30,70,31,252,31,240,31,69,31,66,31,245,31,179,31,193,31,228,31,96,31,232,31,232,30,20,31,153,31,176,31,67,31,67,30,166,31,214,31,140,31,157,31,157,30,121,31,121,30,121,29,9,31,115,31,25,31,194,31,84,31,222,31,123,31,123,30,149,31,100,31,100,30,100,29,63,31,30,31,80,31,80,30,166,31,19,31,10,31,132,31,206,31,217,31,217,30,217,29,194,31,145,31,58,31,124,31,178,31,117,31,117,30,249,31,249,30,249,29,150,31,150,30,150,29,79,31,51,31,157,31,157,30,157,29,197,31,197,30,253,31,253,30,184,31,33,31,33,30,33,29,93,31,138,31,232,31,185,31,131,31,243,31,234,31,241,31,38,31,227,31,116,31,227,31,208,31,251,31,80,31,80,30,80,29,44,31,157,31,150,31,2,31,230,31,137,31,92,31,218,31,178,31,227,31,252,31,143,31,186,31,186,30,105,31,188,31,67,31,67,30,164,31,164,30,128,31,223,31,113,31,102,31,115,31,210,31,210,30,224,31,172,31,156,31,38,31,38,30,125,31,100,31,236,31,188,31,149,31,224,31,150,31,194,31,225,31,85,31,48,31,98,31,217,31,217,30,69,31,28,31,219,31,62,31,62,30,25,31,235,31,17,31,210,31,189,31,136,31,198,31,198,30,204,31,140,31,161,31,161,30,201,31,61,31,231,31,90,31,90,30,200,31,2,31,2,30,184,31,184,30,223,31,61,31,232,31,37,31,138,31,12,31,222,31,235,31,161,31,161,30,61,31,75,31,75,30,180,31,180,30,17,31,17,30,17,29,147,31,147,30,134,31,115,31,83,31,133,31,203,31,221,31,96,31,26,31,160,31,46,31,31,31,31,30,1,31,249,31,255,31,16,31,16,30,159,31,114,31,165,31,161,31,208,31,35,31,55,31,165,31,36,31,36,30,173,31,30,31,7,31,7,30,81,31,81,30,154,31,131,31,132,31,101,31,12,31,12,30,104,31,104,30,104,29,104,28,104,27,41,31,213,31,136,31,59,31,246,31,186,31,252,31,228,31,4,31,185,31,169,31,169,30,149,31,24,31,24,30,165,31,52,31,52,30,216,31,45,31,201,31,253,31,2,31,2,30,2,29,98,31,98,30,9,31,9,30,9,29,9,28,149,31,179,31,166,31,173,31,34,31,34,30,34,29,87,31,87,30,45,31,216,31,138,31,114,31,193,31,193,30,197,31,197,30,199,31,82,31,58,31,42,31,69,31,31,31,169,31,179,31,179,30,221,31,166,31,243,31,38,31,38,30,38,31,29,31,79,31,128,31,251,31,149,31,129,31,95,31,247,31,21,31,42,31,74,31,38,31,180,31,245,31,245,30,245,29,108,31,91,31,136,31,21,31,229,31,184,31,167,31,231,31,231,30,163,31,255,31,255,30,255,29,99,31,99,30,60,31,58,31,59,31,222,31,129,31,163,31,163,30,76,31,191,31,226,31,139,31,140,31,140,30,182,31,182,30,182,29,182,28,182,27,6,31,99,31,212,31,255,31,62,31,169,31,140,31,140,30,56,31,56,30,139,31,10,31,118,31,76,31,81,31,15,31,147,31,195,31,71,31,71,30,28,31,218,31,218,30,244,31,68,31,189,31,229,31,229,30,36,31,158,31,39,31,175,31,224,31,57,31,156,31,236,31,234,31,135,31,6,31,6,30,203,31,64,31,230,31,230,30,97,31,217,31,106,31,106,30,85,31,85,30,125,31,118,31,118,30,197,31,125,31,21,31,164,31,133,31,11,31,41,31,90,31,211,31,10,31,10,30,190,31,190,30,190,29,82,31,101,31,5,31,158,31,48,31,218,31,218,30,188,31,49,31,49,30,255,31,54,31,243,31,150,31,16,31,74,31,74,30,247,31,211,31,152,31,152,30,94,31,80,31,80,30,243,31,2,31,2,30,118,31,58,31,242,31,115,31,175,31,9,31,19,31,75,31,176,31,208,31,231,31,231,30,231,29,231,28,220,31,69,31,74,31,230,31,68,31,34,31,34,30,246,31,246,30,185,31,185,30,185,29,228,31,230,31,88,31,93,31,61,31,144,31,144,30,60,31,60,30,239,31,239,30,207,31,207,30,209,31,89,31,210,31,210,30,210,29,210,28,121,31,156,31,156,30,58,31,139,31,202,31,219,31,131,31,17,31,72,31,121,31,121,30,153,31,68,31,105,31,240,31,188,31,224,31,224,30,204,31,224,31,204,31,206,31,143,31,143,30,39,31,86,31,86,30,86,29,86,28,21,31,248,31,246,31,137,31,137,30,58,31,28,31,241,31,40,31,161,31,161,30,4,31,105,31,18,31,48,31,48,30,145,31,76,31,72,31,122,31,35,31,230,31,68,31,130,31,162,31,174,31,240,31,126,31,24,31,36,31,105,31,181,31,145,31,35,31,226,31,37,31,198,31,198,30,42,31,160,31,217,31,9,31,70,31,8,31,44,31,143,31,75,31,75,30,40,31,212,31,65,31,181,31,155,31,149,31,89,31,184,31,1,31,64,31,214,31,214,30,158,31,162,31,162,30,162,29,126,31,70,31,80,31,186,31,92,31,188,31,188,30,232,31,232,30,232,29,69,31,142,31,142,30,142,29,134,31,187,31,187,30,27,31,225,31,7,31,221,31,191,31,35,31,95,31,149,31,72,31,103,31,222,31,134,31,105,31,105,30,105,29,105,28,101,31,68,31,207,31,196,31,181,31,179,31,215,31,68,31,68,30,68,29,187,31,197,31,20,31,20,30,247,31,12,31,187,31,213,31,15,31,89,31,89,30,89,29,89,28,89,31,64,31,64,30,99,31,173,31,93,31,251,31,64,31,6,31,220,31,168,31,168,30,226,31,155,31,233,31,220,31,220,30,91,31,167,31,34,31,34,30,198,31,101,31,101,30,177,31,177,30,117,31,117,30,217,31,139,31,48,31,210,31,158,31,254,31,160,31,160,30,227,31,227,30,220,31,232,31,42,31,70,31,185,31,183,31,183,30,105,31,174,31,174,30,35,31,33,31,125,31,13,31,46,31,178,31,157,31,58,31,128,31,128,30,251,31,26,31,138,31,56,31,12,31,35,31,11,31,204,31,103,31,246,31,58,31,96,31,82,31,17,31,209,31,96,31,96,30,68,31,219,31,232,31,31,31,219,31,80,31,35,31,35,30,253,31,85,31,175,31,230,31,242,31,247,31,182,31,182,30,170,31,127,31,231,31,201,31,193,31,243,31,15,31,191,31,228,31,249,31,105,31,105,30,40,31,190,31,69,31,113,31,113,30,99,31,24,31,66,31,217,31,16,31,19,31,86,31,139,31,247,31,140,31,140,30,130,31,123,31,72,31,236,31,236,30,210,31,156,31,156,30,137,31,136,31,74,31,152,31,77,31,161,31,181,31,106,31,189,31,189,30,82,31,128,31,109,31,226,31,226,30,204,31,43,31,25,31,195,31,167,31,239,31,129,31,107,31,46,31,230,31,132,31,59,31,90,31,217,31,64,31,64,30,153,31,6,31,6,30,35,31,195,31,130,31,38,31,182,31,207,31,232,31,112,31,38,31,48,31,89,31,143,31,143,30,110,31,225,31,217,31,138,31,10,31,191,31,99,31,111,31,8,31,60,31,60,31,92,31,98,31,81,31,175,31,132,31,79,31,58,31,232,31,224,31,27,31,221,31,221,30,32,31,32,30,139,31,70,31,88,31,86,31,140,31,140,30,19,31,39,31,232,31,178,31,236,31,98,31,98,30,212,31,14,31,24,31,25,31,213,31,21,31,63,31,185,31,185,30,169,31,197,31,129,31,159,31,124,31,124,30,124,29,99,31,209,31,250,31,174,31,161,31,150,31,150,30,202,31,202,30,249,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
