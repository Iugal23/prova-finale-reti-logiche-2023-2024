-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_464 is
end project_tb_464;

architecture project_tb_arch_464 of project_tb_464 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 329;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (225,0,102,0,180,0,220,0,188,0,196,0,179,0,0,0,87,0,140,0,178,0,0,0,93,0,144,0,0,0,197,0,99,0,226,0,249,0,25,0,60,0,25,0,0,0,166,0,118,0,0,0,0,0,155,0,153,0,41,0,215,0,73,0,222,0,15,0,34,0,92,0,4,0,152,0,1,0,0,0,135,0,223,0,73,0,20,0,101,0,130,0,50,0,114,0,0,0,145,0,146,0,0,0,0,0,169,0,217,0,206,0,99,0,0,0,143,0,43,0,0,0,72,0,80,0,0,0,0,0,72,0,197,0,0,0,22,0,0,0,0,0,219,0,221,0,0,0,122,0,158,0,0,0,127,0,69,0,112,0,163,0,48,0,235,0,212,0,208,0,47,0,127,0,212,0,0,0,221,0,48,0,99,0,56,0,111,0,245,0,37,0,71,0,0,0,0,0,169,0,184,0,0,0,208,0,0,0,0,0,82,0,150,0,169,0,87,0,0,0,51,0,94,0,0,0,0,0,13,0,80,0,141,0,41,0,55,0,0,0,45,0,242,0,66,0,0,0,239,0,23,0,0,0,231,0,71,0,159,0,240,0,0,0,0,0,136,0,196,0,114,0,33,0,80,0,0,0,207,0,17,0,150,0,48,0,60,0,37,0,49,0,192,0,12,0,202,0,58,0,80,0,89,0,146,0,202,0,205,0,210,0,148,0,209,0,220,0,132,0,106,0,0,0,115,0,132,0,4,0,238,0,33,0,107,0,0,0,23,0,166,0,109,0,202,0,165,0,7,0,102,0,0,0,27,0,0,0,190,0,95,0,0,0,175,0,44,0,251,0,0,0,65,0,188,0,37,0,9,0,110,0,0,0,3,0,161,0,226,0,61,0,26,0,129,0,251,0,28,0,32,0,252,0,178,0,165,0,14,0,0,0,0,0,2,0,186,0,53,0,82,0,17,0,0,0,0,0,0,0,0,0,53,0,190,0,52,0,70,0,0,0,206,0,161,0,0,0,228,0,0,0,253,0,0,0,230,0,0,0,237,0,42,0,175,0,239,0,53,0,0,0,159,0,32,0,0,0,163,0,74,0,0,0,228,0,239,0,18,0,19,0,255,0,23,0,103,0,62,0,239,0,178,0,218,0,12,0,206,0,126,0,176,0,0,0,0,0,0,0,231,0,237,0,0,0,213,0,218,0,196,0,27,0,130,0,244,0,126,0,176,0,72,0,45,0,0,0,63,0,20,0,0,0,215,0,136,0,0,0,254,0,94,0,218,0,80,0,37,0,212,0,81,0,9,0,255,0,253,0,0,0,135,0,45,0,37,0,0,0,106,0,0,0,196,0,177,0,102,0,252,0,127,0,95,0,65,0,36,0,168,0,218,0,165,0,0,0,208,0,170,0,87,0,159,0,0,0,66,0,59,0,165,0,106,0,128,0,229,0,0,0,0,0,160,0,91,0,110,0,145,0,208,0,136,0,19,0);
signal scenario_full  : scenario_type := (225,31,102,31,180,31,220,31,188,31,196,31,179,31,179,30,87,31,140,31,178,31,178,30,93,31,144,31,144,30,197,31,99,31,226,31,249,31,25,31,60,31,25,31,25,30,166,31,118,31,118,30,118,29,155,31,153,31,41,31,215,31,73,31,222,31,15,31,34,31,92,31,4,31,152,31,1,31,1,30,135,31,223,31,73,31,20,31,101,31,130,31,50,31,114,31,114,30,145,31,146,31,146,30,146,29,169,31,217,31,206,31,99,31,99,30,143,31,43,31,43,30,72,31,80,31,80,30,80,29,72,31,197,31,197,30,22,31,22,30,22,29,219,31,221,31,221,30,122,31,158,31,158,30,127,31,69,31,112,31,163,31,48,31,235,31,212,31,208,31,47,31,127,31,212,31,212,30,221,31,48,31,99,31,56,31,111,31,245,31,37,31,71,31,71,30,71,29,169,31,184,31,184,30,208,31,208,30,208,29,82,31,150,31,169,31,87,31,87,30,51,31,94,31,94,30,94,29,13,31,80,31,141,31,41,31,55,31,55,30,45,31,242,31,66,31,66,30,239,31,23,31,23,30,231,31,71,31,159,31,240,31,240,30,240,29,136,31,196,31,114,31,33,31,80,31,80,30,207,31,17,31,150,31,48,31,60,31,37,31,49,31,192,31,12,31,202,31,58,31,80,31,89,31,146,31,202,31,205,31,210,31,148,31,209,31,220,31,132,31,106,31,106,30,115,31,132,31,4,31,238,31,33,31,107,31,107,30,23,31,166,31,109,31,202,31,165,31,7,31,102,31,102,30,27,31,27,30,190,31,95,31,95,30,175,31,44,31,251,31,251,30,65,31,188,31,37,31,9,31,110,31,110,30,3,31,161,31,226,31,61,31,26,31,129,31,251,31,28,31,32,31,252,31,178,31,165,31,14,31,14,30,14,29,2,31,186,31,53,31,82,31,17,31,17,30,17,29,17,28,17,27,53,31,190,31,52,31,70,31,70,30,206,31,161,31,161,30,228,31,228,30,253,31,253,30,230,31,230,30,237,31,42,31,175,31,239,31,53,31,53,30,159,31,32,31,32,30,163,31,74,31,74,30,228,31,239,31,18,31,19,31,255,31,23,31,103,31,62,31,239,31,178,31,218,31,12,31,206,31,126,31,176,31,176,30,176,29,176,28,231,31,237,31,237,30,213,31,218,31,196,31,27,31,130,31,244,31,126,31,176,31,72,31,45,31,45,30,63,31,20,31,20,30,215,31,136,31,136,30,254,31,94,31,218,31,80,31,37,31,212,31,81,31,9,31,255,31,253,31,253,30,135,31,45,31,37,31,37,30,106,31,106,30,196,31,177,31,102,31,252,31,127,31,95,31,65,31,36,31,168,31,218,31,165,31,165,30,208,31,170,31,87,31,159,31,159,30,66,31,59,31,165,31,106,31,128,31,229,31,229,30,229,29,160,31,91,31,110,31,145,31,208,31,136,31,19,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
