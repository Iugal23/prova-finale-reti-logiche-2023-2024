-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 764;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (75,0,146,0,158,0,60,0,0,0,0,0,108,0,77,0,34,0,126,0,31,0,14,0,98,0,0,0,225,0,32,0,114,0,0,0,56,0,166,0,0,0,136,0,0,0,0,0,246,0,0,0,160,0,0,0,11,0,36,0,168,0,55,0,131,0,48,0,0,0,180,0,103,0,0,0,0,0,202,0,123,0,28,0,198,0,29,0,0,0,110,0,231,0,43,0,52,0,123,0,0,0,81,0,221,0,32,0,214,0,168,0,220,0,71,0,0,0,52,0,135,0,147,0,130,0,0,0,6,0,19,0,43,0,227,0,146,0,184,0,176,0,0,0,0,0,190,0,89,0,21,0,194,0,50,0,102,0,226,0,146,0,0,0,0,0,142,0,122,0,29,0,50,0,0,0,0,0,141,0,214,0,0,0,0,0,156,0,35,0,0,0,0,0,138,0,109,0,15,0,126,0,9,0,63,0,142,0,0,0,118,0,217,0,0,0,0,0,231,0,53,0,50,0,160,0,4,0,152,0,65,0,190,0,198,0,138,0,34,0,162,0,186,0,83,0,165,0,80,0,0,0,105,0,65,0,33,0,147,0,220,0,126,0,229,0,119,0,0,0,60,0,119,0,129,0,247,0,33,0,140,0,88,0,135,0,56,0,167,0,36,0,0,0,208,0,151,0,251,0,70,0,72,0,146,0,142,0,130,0,0,0,154,0,73,0,0,0,122,0,137,0,62,0,90,0,163,0,0,0,144,0,233,0,123,0,183,0,0,0,119,0,234,0,12,0,0,0,236,0,30,0,209,0,0,0,5,0,50,0,69,0,0,0,55,0,148,0,44,0,220,0,144,0,56,0,239,0,150,0,179,0,0,0,96,0,36,0,0,0,99,0,0,0,141,0,199,0,109,0,183,0,84,0,154,0,187,0,152,0,69,0,176,0,138,0,39,0,196,0,0,0,139,0,160,0,221,0,90,0,0,0,0,0,12,0,0,0,82,0,195,0,82,0,37,0,126,0,112,0,2,0,4,0,80,0,102,0,165,0,32,0,140,0,120,0,165,0,0,0,98,0,0,0,203,0,227,0,217,0,0,0,250,0,41,0,23,0,52,0,3,0,77,0,160,0,115,0,151,0,183,0,44,0,160,0,0,0,233,0,80,0,193,0,235,0,134,0,0,0,182,0,22,0,54,0,0,0,0,0,0,0,0,0,0,0,201,0,190,0,49,0,147,0,159,0,116,0,133,0,106,0,31,0,60,0,98,0,25,0,143,0,161,0,145,0,202,0,0,0,101,0,106,0,168,0,0,0,106,0,26,0,52,0,40,0,239,0,38,0,40,0,132,0,137,0,171,0,175,0,0,0,36,0,95,0,63,0,203,0,0,0,25,0,156,0,21,0,197,0,0,0,0,0,235,0,194,0,70,0,194,0,79,0,0,0,0,0,254,0,207,0,133,0,33,0,0,0,217,0,98,0,158,0,82,0,252,0,245,0,153,0,0,0,140,0,0,0,10,0,25,0,41,0,126,0,184,0,156,0,195,0,14,0,2,0,20,0,108,0,0,0,64,0,6,0,0,0,0,0,0,0,171,0,200,0,0,0,0,0,126,0,239,0,183,0,155,0,229,0,208,0,40,0,200,0,28,0,120,0,195,0,150,0,152,0,164,0,125,0,50,0,238,0,217,0,15,0,145,0,222,0,163,0,103,0,248,0,151,0,35,0,154,0,76,0,143,0,208,0,42,0,144,0,0,0,110,0,251,0,226,0,65,0,174,0,51,0,4,0,58,0,219,0,170,0,200,0,236,0,141,0,163,0,0,0,0,0,0,0,0,0,98,0,0,0,0,0,65,0,170,0,209,0,99,0,62,0,201,0,228,0,15,0,77,0,0,0,196,0,0,0,26,0,71,0,220,0,30,0,67,0,250,0,164,0,219,0,244,0,0,0,0,0,0,0,28,0,0,0,248,0,238,0,22,0,0,0,178,0,0,0,254,0,145,0,53,0,79,0,179,0,0,0,3,0,0,0,155,0,5,0,215,0,223,0,0,0,65,0,55,0,0,0,84,0,171,0,0,0,133,0,90,0,218,0,0,0,186,0,243,0,185,0,46,0,42,0,216,0,219,0,65,0,238,0,7,0,53,0,131,0,60,0,13,0,161,0,49,0,0,0,0,0,112,0,19,0,111,0,51,0,38,0,134,0,102,0,22,0,0,0,84,0,172,0,87,0,52,0,159,0,128,0,123,0,82,0,193,0,31,0,137,0,0,0,28,0,48,0,229,0,111,0,219,0,175,0,66,0,47,0,121,0,0,0,192,0,89,0,35,0,34,0,26,0,140,0,92,0,0,0,0,0,0,0,128,0,106,0,0,0,45,0,192,0,101,0,59,0,143,0,138,0,99,0,195,0,79,0,0,0,0,0,63,0,221,0,123,0,75,0,156,0,0,0,0,0,0,0,175,0,215,0,198,0,240,0,68,0,0,0,224,0,0,0,0,0,156,0,0,0,43,0,3,0,91,0,180,0,127,0,188,0,5,0,0,0,38,0,42,0,163,0,238,0,83,0,2,0,121,0,228,0,182,0,242,0,86,0,236,0,249,0,143,0,176,0,203,0,117,0,11,0,6,0,37,0,102,0,0,0,0,0,0,0,239,0,20,0,73,0,0,0,0,0,164,0,0,0,162,0,254,0,189,0,36,0,210,0,0,0,0,0,0,0,167,0,138,0,0,0,217,0,94,0,24,0,248,0,199,0,142,0,120,0,17,0,95,0,206,0,44,0,158,0,0,0,1,0,0,0,124,0,134,0,180,0,0,0,0,0,176,0,122,0,0,0,36,0,0,0,0,0,79,0,23,0,95,0,37,0,115,0,0,0,30,0,115,0,133,0,0,0,0,0,188,0,73,0,16,0,0,0,98,0,231,0,77,0,0,0,0,0,0,0,219,0,136,0,29,0,248,0,74,0,250,0,64,0,224,0,10,0,0,0,117,0,0,0,222,0,109,0,96,0,0,0,138,0,114,0,217,0,231,0,112,0,150,0,89,0,114,0,0,0,0,0,218,0,0,0,208,0,26,0,0,0,0,0,128,0,134,0,47,0,186,0,15,0,189,0,50,0,0,0,63,0,143,0,227,0,0,0,0,0,0,0,156,0,136,0,0,0,20,0,0,0,200,0,0,0,226,0,15,0,234,0,128,0,57,0,106,0,32,0,145,0,156,0,0,0,0,0,224,0,145,0,248,0,16,0,183,0,35,0,126,0,31,0,200,0,0,0,0,0,68,0,62,0,171,0,110,0,172,0,118,0,235,0,159,0,232,0,134,0,219,0,213,0,0,0,239,0,21,0,87,0,49,0,225,0,118,0,89,0,83,0,0,0,0,0,90,0,0,0,168,0,33,0,40,0,65,0,134,0,126,0,23,0,108,0,0,0,213,0,0,0);
signal scenario_full  : scenario_type := (75,31,146,31,158,31,60,31,60,30,60,29,108,31,77,31,34,31,126,31,31,31,14,31,98,31,98,30,225,31,32,31,114,31,114,30,56,31,166,31,166,30,136,31,136,30,136,29,246,31,246,30,160,31,160,30,11,31,36,31,168,31,55,31,131,31,48,31,48,30,180,31,103,31,103,30,103,29,202,31,123,31,28,31,198,31,29,31,29,30,110,31,231,31,43,31,52,31,123,31,123,30,81,31,221,31,32,31,214,31,168,31,220,31,71,31,71,30,52,31,135,31,147,31,130,31,130,30,6,31,19,31,43,31,227,31,146,31,184,31,176,31,176,30,176,29,190,31,89,31,21,31,194,31,50,31,102,31,226,31,146,31,146,30,146,29,142,31,122,31,29,31,50,31,50,30,50,29,141,31,214,31,214,30,214,29,156,31,35,31,35,30,35,29,138,31,109,31,15,31,126,31,9,31,63,31,142,31,142,30,118,31,217,31,217,30,217,29,231,31,53,31,50,31,160,31,4,31,152,31,65,31,190,31,198,31,138,31,34,31,162,31,186,31,83,31,165,31,80,31,80,30,105,31,65,31,33,31,147,31,220,31,126,31,229,31,119,31,119,30,60,31,119,31,129,31,247,31,33,31,140,31,88,31,135,31,56,31,167,31,36,31,36,30,208,31,151,31,251,31,70,31,72,31,146,31,142,31,130,31,130,30,154,31,73,31,73,30,122,31,137,31,62,31,90,31,163,31,163,30,144,31,233,31,123,31,183,31,183,30,119,31,234,31,12,31,12,30,236,31,30,31,209,31,209,30,5,31,50,31,69,31,69,30,55,31,148,31,44,31,220,31,144,31,56,31,239,31,150,31,179,31,179,30,96,31,36,31,36,30,99,31,99,30,141,31,199,31,109,31,183,31,84,31,154,31,187,31,152,31,69,31,176,31,138,31,39,31,196,31,196,30,139,31,160,31,221,31,90,31,90,30,90,29,12,31,12,30,82,31,195,31,82,31,37,31,126,31,112,31,2,31,4,31,80,31,102,31,165,31,32,31,140,31,120,31,165,31,165,30,98,31,98,30,203,31,227,31,217,31,217,30,250,31,41,31,23,31,52,31,3,31,77,31,160,31,115,31,151,31,183,31,44,31,160,31,160,30,233,31,80,31,193,31,235,31,134,31,134,30,182,31,22,31,54,31,54,30,54,29,54,28,54,27,54,26,201,31,190,31,49,31,147,31,159,31,116,31,133,31,106,31,31,31,60,31,98,31,25,31,143,31,161,31,145,31,202,31,202,30,101,31,106,31,168,31,168,30,106,31,26,31,52,31,40,31,239,31,38,31,40,31,132,31,137,31,171,31,175,31,175,30,36,31,95,31,63,31,203,31,203,30,25,31,156,31,21,31,197,31,197,30,197,29,235,31,194,31,70,31,194,31,79,31,79,30,79,29,254,31,207,31,133,31,33,31,33,30,217,31,98,31,158,31,82,31,252,31,245,31,153,31,153,30,140,31,140,30,10,31,25,31,41,31,126,31,184,31,156,31,195,31,14,31,2,31,20,31,108,31,108,30,64,31,6,31,6,30,6,29,6,28,171,31,200,31,200,30,200,29,126,31,239,31,183,31,155,31,229,31,208,31,40,31,200,31,28,31,120,31,195,31,150,31,152,31,164,31,125,31,50,31,238,31,217,31,15,31,145,31,222,31,163,31,103,31,248,31,151,31,35,31,154,31,76,31,143,31,208,31,42,31,144,31,144,30,110,31,251,31,226,31,65,31,174,31,51,31,4,31,58,31,219,31,170,31,200,31,236,31,141,31,163,31,163,30,163,29,163,28,163,27,98,31,98,30,98,29,65,31,170,31,209,31,99,31,62,31,201,31,228,31,15,31,77,31,77,30,196,31,196,30,26,31,71,31,220,31,30,31,67,31,250,31,164,31,219,31,244,31,244,30,244,29,244,28,28,31,28,30,248,31,238,31,22,31,22,30,178,31,178,30,254,31,145,31,53,31,79,31,179,31,179,30,3,31,3,30,155,31,5,31,215,31,223,31,223,30,65,31,55,31,55,30,84,31,171,31,171,30,133,31,90,31,218,31,218,30,186,31,243,31,185,31,46,31,42,31,216,31,219,31,65,31,238,31,7,31,53,31,131,31,60,31,13,31,161,31,49,31,49,30,49,29,112,31,19,31,111,31,51,31,38,31,134,31,102,31,22,31,22,30,84,31,172,31,87,31,52,31,159,31,128,31,123,31,82,31,193,31,31,31,137,31,137,30,28,31,48,31,229,31,111,31,219,31,175,31,66,31,47,31,121,31,121,30,192,31,89,31,35,31,34,31,26,31,140,31,92,31,92,30,92,29,92,28,128,31,106,31,106,30,45,31,192,31,101,31,59,31,143,31,138,31,99,31,195,31,79,31,79,30,79,29,63,31,221,31,123,31,75,31,156,31,156,30,156,29,156,28,175,31,215,31,198,31,240,31,68,31,68,30,224,31,224,30,224,29,156,31,156,30,43,31,3,31,91,31,180,31,127,31,188,31,5,31,5,30,38,31,42,31,163,31,238,31,83,31,2,31,121,31,228,31,182,31,242,31,86,31,236,31,249,31,143,31,176,31,203,31,117,31,11,31,6,31,37,31,102,31,102,30,102,29,102,28,239,31,20,31,73,31,73,30,73,29,164,31,164,30,162,31,254,31,189,31,36,31,210,31,210,30,210,29,210,28,167,31,138,31,138,30,217,31,94,31,24,31,248,31,199,31,142,31,120,31,17,31,95,31,206,31,44,31,158,31,158,30,1,31,1,30,124,31,134,31,180,31,180,30,180,29,176,31,122,31,122,30,36,31,36,30,36,29,79,31,23,31,95,31,37,31,115,31,115,30,30,31,115,31,133,31,133,30,133,29,188,31,73,31,16,31,16,30,98,31,231,31,77,31,77,30,77,29,77,28,219,31,136,31,29,31,248,31,74,31,250,31,64,31,224,31,10,31,10,30,117,31,117,30,222,31,109,31,96,31,96,30,138,31,114,31,217,31,231,31,112,31,150,31,89,31,114,31,114,30,114,29,218,31,218,30,208,31,26,31,26,30,26,29,128,31,134,31,47,31,186,31,15,31,189,31,50,31,50,30,63,31,143,31,227,31,227,30,227,29,227,28,156,31,136,31,136,30,20,31,20,30,200,31,200,30,226,31,15,31,234,31,128,31,57,31,106,31,32,31,145,31,156,31,156,30,156,29,224,31,145,31,248,31,16,31,183,31,35,31,126,31,31,31,200,31,200,30,200,29,68,31,62,31,171,31,110,31,172,31,118,31,235,31,159,31,232,31,134,31,219,31,213,31,213,30,239,31,21,31,87,31,49,31,225,31,118,31,89,31,83,31,83,30,83,29,90,31,90,30,168,31,33,31,40,31,65,31,134,31,126,31,23,31,108,31,108,30,213,31,213,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
