-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_527 is
end project_tb_527;

architecture project_tb_arch_527 of project_tb_527 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 805;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (245,0,0,0,146,0,125,0,75,0,164,0,103,0,179,0,42,0,110,0,150,0,71,0,126,0,0,0,0,0,37,0,0,0,111,0,160,0,10,0,0,0,27,0,20,0,180,0,165,0,209,0,0,0,180,0,52,0,158,0,22,0,116,0,70,0,64,0,74,0,187,0,2,0,17,0,129,0,63,0,232,0,139,0,156,0,0,0,184,0,189,0,102,0,0,0,164,0,134,0,0,0,189,0,11,0,138,0,213,0,76,0,215,0,219,0,81,0,193,0,238,0,187,0,197,0,218,0,40,0,58,0,0,0,224,0,0,0,0,0,156,0,46,0,158,0,234,0,0,0,52,0,157,0,0,0,58,0,67,0,172,0,109,0,0,0,30,0,115,0,192,0,28,0,0,0,178,0,174,0,164,0,10,0,0,0,51,0,0,0,80,0,127,0,134,0,0,0,100,0,0,0,94,0,246,0,0,0,194,0,97,0,145,0,122,0,24,0,78,0,0,0,170,0,249,0,142,0,40,0,0,0,82,0,150,0,124,0,76,0,0,0,57,0,5,0,238,0,120,0,148,0,133,0,148,0,190,0,0,0,195,0,181,0,20,0,0,0,33,0,167,0,235,0,0,0,158,0,239,0,28,0,241,0,144,0,80,0,87,0,0,0,167,0,83,0,7,0,18,0,71,0,75,0,99,0,223,0,201,0,89,0,193,0,71,0,53,0,184,0,19,0,255,0,110,0,250,0,48,0,4,0,173,0,130,0,69,0,3,0,18,0,128,0,115,0,0,0,162,0,0,0,41,0,102,0,207,0,90,0,211,0,153,0,199,0,99,0,0,0,148,0,61,0,232,0,217,0,0,0,0,0,0,0,250,0,0,0,117,0,67,0,198,0,0,0,0,0,69,0,248,0,139,0,235,0,130,0,222,0,0,0,141,0,0,0,124,0,202,0,7,0,0,0,0,0,106,0,0,0,170,0,0,0,0,0,204,0,0,0,106,0,90,0,67,0,210,0,192,0,0,0,165,0,0,0,115,0,0,0,0,0,36,0,87,0,85,0,79,0,127,0,0,0,120,0,0,0,161,0,127,0,11,0,0,0,215,0,9,0,113,0,84,0,99,0,125,0,184,0,100,0,57,0,0,0,209,0,237,0,137,0,181,0,0,0,149,0,75,0,86,0,67,0,1,0,147,0,0,0,170,0,91,0,191,0,237,0,59,0,195,0,0,0,0,0,12,0,55,0,189,0,58,0,157,0,87,0,100,0,104,0,157,0,83,0,206,0,151,0,137,0,133,0,32,0,37,0,126,0,0,0,19,0,171,0,161,0,165,0,0,0,100,0,0,0,236,0,133,0,186,0,33,0,214,0,43,0,188,0,0,0,167,0,0,0,231,0,0,0,162,0,41,0,160,0,104,0,217,0,141,0,175,0,209,0,221,0,0,0,214,0,174,0,200,0,99,0,43,0,159,0,154,0,108,0,140,0,195,0,119,0,168,0,93,0,13,0,103,0,189,0,60,0,91,0,0,0,0,0,0,0,130,0,242,0,0,0,136,0,0,0,0,0,112,0,247,0,74,0,252,0,188,0,20,0,192,0,136,0,13,0,61,0,65,0,0,0,8,0,249,0,163,0,235,0,234,0,200,0,152,0,202,0,0,0,0,0,182,0,0,0,220,0,0,0,234,0,35,0,0,0,252,0,205,0,141,0,0,0,205,0,0,0,157,0,55,0,205,0,215,0,0,0,75,0,170,0,159,0,0,0,0,0,204,0,0,0,74,0,0,0,90,0,0,0,253,0,108,0,128,0,175,0,0,0,42,0,210,0,0,0,172,0,7,0,56,0,0,0,109,0,212,0,137,0,0,0,115,0,254,0,0,0,239,0,50,0,125,0,27,0,52,0,23,0,119,0,0,0,8,0,15,0,69,0,68,0,9,0,226,0,72,0,0,0,70,0,0,0,126,0,118,0,0,0,79,0,183,0,27,0,174,0,146,0,55,0,89,0,99,0,78,0,133,0,222,0,129,0,0,0,70,0,241,0,200,0,1,0,33,0,185,0,122,0,9,0,0,0,190,0,82,0,12,0,33,0,12,0,224,0,0,0,0,0,0,0,194,0,107,0,130,0,115,0,110,0,192,0,99,0,36,0,71,0,238,0,0,0,172,0,105,0,64,0,21,0,0,0,142,0,0,0,8,0,67,0,151,0,149,0,83,0,222,0,123,0,144,0,190,0,250,0,236,0,0,0,241,0,0,0,72,0,13,0,134,0,206,0,194,0,171,0,91,0,174,0,37,0,0,0,67,0,79,0,251,0,86,0,167,0,191,0,57,0,110,0,203,0,254,0,164,0,79,0,4,0,48,0,139,0,51,0,25,0,136,0,203,0,255,0,108,0,0,0,229,0,100,0,62,0,0,0,195,0,227,0,136,0,154,0,61,0,0,0,0,0,28,0,219,0,222,0,0,0,106,0,188,0,125,0,95,0,225,0,172,0,106,0,116,0,157,0,235,0,0,0,57,0,0,0,216,0,204,0,67,0,97,0,36,0,0,0,170,0,223,0,69,0,118,0,127,0,75,0,0,0,16,0,133,0,255,0,66,0,194,0,0,0,0,0,181,0,230,0,233,0,17,0,151,0,193,0,53,0,144,0,35,0,188,0,18,0,172,0,234,0,176,0,217,0,246,0,0,0,152,0,85,0,68,0,142,0,167,0,181,0,0,0,191,0,41,0,209,0,0,0,41,0,253,0,191,0,59,0,90,0,213,0,29,0,152,0,142,0,158,0,0,0,216,0,106,0,226,0,167,0,4,0,207,0,0,0,35,0,2,0,80,0,0,0,20,0,0,0,245,0,202,0,206,0,252,0,0,0,139,0,215,0,170,0,29,0,27,0,188,0,44,0,28,0,158,0,72,0,11,0,19,0,193,0,0,0,0,0,116,0,0,0,200,0,205,0,11,0,0,0,33,0,206,0,29,0,116,0,108,0,173,0,230,0,140,0,167,0,116,0,208,0,246,0,187,0,78,0,17,0,0,0,0,0,200,0,35,0,237,0,89,0,4,0,63,0,134,0,0,0,123,0,150,0,64,0,8,0,239,0,218,0,0,0,0,0,196,0,73,0,0,0,0,0,0,0,65,0,134,0,91,0,74,0,7,0,0,0,111,0,57,0,189,0,67,0,178,0,196,0,46,0,89,0,216,0,0,0,125,0,0,0,241,0,149,0,136,0,120,0,234,0,151,0,49,0,161,0,133,0,137,0,0,0,85,0,206,0,119,0,0,0,235,0,41,0,12,0,154,0,195,0,9,0,142,0,224,0,76,0,77,0,94,0,175,0,231,0,76,0,119,0,51,0,141,0,245,0,11,0,79,0,0,0,132,0,48,0,0,0,183,0,192,0,135,0,99,0,72,0,145,0,163,0,226,0,112,0,135,0,163,0,233,0,0,0,77,0,138,0,86,0,167,0,54,0,100,0,0,0,228,0,169,0,231,0,38,0,160,0,65,0,0,0,0,0,79,0,0,0,192,0,6,0,112,0,218,0,89,0,214,0,0,0,0,0,0,0,78,0,1,0,42,0,233,0,163,0,187,0,228,0,213,0,40,0,157,0,67,0,234,0);
signal scenario_full  : scenario_type := (245,31,245,30,146,31,125,31,75,31,164,31,103,31,179,31,42,31,110,31,150,31,71,31,126,31,126,30,126,29,37,31,37,30,111,31,160,31,10,31,10,30,27,31,20,31,180,31,165,31,209,31,209,30,180,31,52,31,158,31,22,31,116,31,70,31,64,31,74,31,187,31,2,31,17,31,129,31,63,31,232,31,139,31,156,31,156,30,184,31,189,31,102,31,102,30,164,31,134,31,134,30,189,31,11,31,138,31,213,31,76,31,215,31,219,31,81,31,193,31,238,31,187,31,197,31,218,31,40,31,58,31,58,30,224,31,224,30,224,29,156,31,46,31,158,31,234,31,234,30,52,31,157,31,157,30,58,31,67,31,172,31,109,31,109,30,30,31,115,31,192,31,28,31,28,30,178,31,174,31,164,31,10,31,10,30,51,31,51,30,80,31,127,31,134,31,134,30,100,31,100,30,94,31,246,31,246,30,194,31,97,31,145,31,122,31,24,31,78,31,78,30,170,31,249,31,142,31,40,31,40,30,82,31,150,31,124,31,76,31,76,30,57,31,5,31,238,31,120,31,148,31,133,31,148,31,190,31,190,30,195,31,181,31,20,31,20,30,33,31,167,31,235,31,235,30,158,31,239,31,28,31,241,31,144,31,80,31,87,31,87,30,167,31,83,31,7,31,18,31,71,31,75,31,99,31,223,31,201,31,89,31,193,31,71,31,53,31,184,31,19,31,255,31,110,31,250,31,48,31,4,31,173,31,130,31,69,31,3,31,18,31,128,31,115,31,115,30,162,31,162,30,41,31,102,31,207,31,90,31,211,31,153,31,199,31,99,31,99,30,148,31,61,31,232,31,217,31,217,30,217,29,217,28,250,31,250,30,117,31,67,31,198,31,198,30,198,29,69,31,248,31,139,31,235,31,130,31,222,31,222,30,141,31,141,30,124,31,202,31,7,31,7,30,7,29,106,31,106,30,170,31,170,30,170,29,204,31,204,30,106,31,90,31,67,31,210,31,192,31,192,30,165,31,165,30,115,31,115,30,115,29,36,31,87,31,85,31,79,31,127,31,127,30,120,31,120,30,161,31,127,31,11,31,11,30,215,31,9,31,113,31,84,31,99,31,125,31,184,31,100,31,57,31,57,30,209,31,237,31,137,31,181,31,181,30,149,31,75,31,86,31,67,31,1,31,147,31,147,30,170,31,91,31,191,31,237,31,59,31,195,31,195,30,195,29,12,31,55,31,189,31,58,31,157,31,87,31,100,31,104,31,157,31,83,31,206,31,151,31,137,31,133,31,32,31,37,31,126,31,126,30,19,31,171,31,161,31,165,31,165,30,100,31,100,30,236,31,133,31,186,31,33,31,214,31,43,31,188,31,188,30,167,31,167,30,231,31,231,30,162,31,41,31,160,31,104,31,217,31,141,31,175,31,209,31,221,31,221,30,214,31,174,31,200,31,99,31,43,31,159,31,154,31,108,31,140,31,195,31,119,31,168,31,93,31,13,31,103,31,189,31,60,31,91,31,91,30,91,29,91,28,130,31,242,31,242,30,136,31,136,30,136,29,112,31,247,31,74,31,252,31,188,31,20,31,192,31,136,31,13,31,61,31,65,31,65,30,8,31,249,31,163,31,235,31,234,31,200,31,152,31,202,31,202,30,202,29,182,31,182,30,220,31,220,30,234,31,35,31,35,30,252,31,205,31,141,31,141,30,205,31,205,30,157,31,55,31,205,31,215,31,215,30,75,31,170,31,159,31,159,30,159,29,204,31,204,30,74,31,74,30,90,31,90,30,253,31,108,31,128,31,175,31,175,30,42,31,210,31,210,30,172,31,7,31,56,31,56,30,109,31,212,31,137,31,137,30,115,31,254,31,254,30,239,31,50,31,125,31,27,31,52,31,23,31,119,31,119,30,8,31,15,31,69,31,68,31,9,31,226,31,72,31,72,30,70,31,70,30,126,31,118,31,118,30,79,31,183,31,27,31,174,31,146,31,55,31,89,31,99,31,78,31,133,31,222,31,129,31,129,30,70,31,241,31,200,31,1,31,33,31,185,31,122,31,9,31,9,30,190,31,82,31,12,31,33,31,12,31,224,31,224,30,224,29,224,28,194,31,107,31,130,31,115,31,110,31,192,31,99,31,36,31,71,31,238,31,238,30,172,31,105,31,64,31,21,31,21,30,142,31,142,30,8,31,67,31,151,31,149,31,83,31,222,31,123,31,144,31,190,31,250,31,236,31,236,30,241,31,241,30,72,31,13,31,134,31,206,31,194,31,171,31,91,31,174,31,37,31,37,30,67,31,79,31,251,31,86,31,167,31,191,31,57,31,110,31,203,31,254,31,164,31,79,31,4,31,48,31,139,31,51,31,25,31,136,31,203,31,255,31,108,31,108,30,229,31,100,31,62,31,62,30,195,31,227,31,136,31,154,31,61,31,61,30,61,29,28,31,219,31,222,31,222,30,106,31,188,31,125,31,95,31,225,31,172,31,106,31,116,31,157,31,235,31,235,30,57,31,57,30,216,31,204,31,67,31,97,31,36,31,36,30,170,31,223,31,69,31,118,31,127,31,75,31,75,30,16,31,133,31,255,31,66,31,194,31,194,30,194,29,181,31,230,31,233,31,17,31,151,31,193,31,53,31,144,31,35,31,188,31,18,31,172,31,234,31,176,31,217,31,246,31,246,30,152,31,85,31,68,31,142,31,167,31,181,31,181,30,191,31,41,31,209,31,209,30,41,31,253,31,191,31,59,31,90,31,213,31,29,31,152,31,142,31,158,31,158,30,216,31,106,31,226,31,167,31,4,31,207,31,207,30,35,31,2,31,80,31,80,30,20,31,20,30,245,31,202,31,206,31,252,31,252,30,139,31,215,31,170,31,29,31,27,31,188,31,44,31,28,31,158,31,72,31,11,31,19,31,193,31,193,30,193,29,116,31,116,30,200,31,205,31,11,31,11,30,33,31,206,31,29,31,116,31,108,31,173,31,230,31,140,31,167,31,116,31,208,31,246,31,187,31,78,31,17,31,17,30,17,29,200,31,35,31,237,31,89,31,4,31,63,31,134,31,134,30,123,31,150,31,64,31,8,31,239,31,218,31,218,30,218,29,196,31,73,31,73,30,73,29,73,28,65,31,134,31,91,31,74,31,7,31,7,30,111,31,57,31,189,31,67,31,178,31,196,31,46,31,89,31,216,31,216,30,125,31,125,30,241,31,149,31,136,31,120,31,234,31,151,31,49,31,161,31,133,31,137,31,137,30,85,31,206,31,119,31,119,30,235,31,41,31,12,31,154,31,195,31,9,31,142,31,224,31,76,31,77,31,94,31,175,31,231,31,76,31,119,31,51,31,141,31,245,31,11,31,79,31,79,30,132,31,48,31,48,30,183,31,192,31,135,31,99,31,72,31,145,31,163,31,226,31,112,31,135,31,163,31,233,31,233,30,77,31,138,31,86,31,167,31,54,31,100,31,100,30,228,31,169,31,231,31,38,31,160,31,65,31,65,30,65,29,79,31,79,30,192,31,6,31,112,31,218,31,89,31,214,31,214,30,214,29,214,28,78,31,1,31,42,31,233,31,163,31,187,31,228,31,213,31,40,31,157,31,67,31,234,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
