-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_790 is
end project_tb_790;

architecture project_tb_arch_790 of project_tb_790 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1020;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,22,0,0,0,0,0,62,0,102,0,0,0,133,0,180,0,0,0,45,0,204,0,244,0,155,0,209,0,166,0,0,0,70,0,0,0,0,0,8,0,221,0,19,0,178,0,187,0,8,0,64,0,8,0,42,0,0,0,70,0,180,0,124,0,39,0,0,0,78,0,129,0,179,0,22,0,176,0,0,0,218,0,0,0,121,0,54,0,57,0,35,0,0,0,112,0,56,0,115,0,168,0,44,0,146,0,198,0,52,0,132,0,236,0,21,0,66,0,134,0,23,0,0,0,129,0,160,0,245,0,100,0,0,0,96,0,0,0,189,0,89,0,82,0,153,0,123,0,0,0,162,0,0,0,107,0,206,0,48,0,254,0,221,0,129,0,114,0,9,0,2,0,185,0,162,0,19,0,151,0,0,0,0,0,217,0,80,0,14,0,11,0,232,0,226,0,34,0,63,0,84,0,34,0,135,0,108,0,73,0,0,0,169,0,118,0,0,0,0,0,0,0,0,0,177,0,22,0,14,0,114,0,253,0,223,0,9,0,243,0,14,0,137,0,0,0,211,0,0,0,164,0,93,0,222,0,137,0,142,0,210,0,137,0,240,0,152,0,239,0,235,0,0,0,41,0,89,0,7,0,166,0,194,0,0,0,170,0,64,0,163,0,0,0,136,0,0,0,0,0,181,0,78,0,238,0,0,0,0,0,1,0,12,0,188,0,236,0,129,0,31,0,82,0,0,0,53,0,251,0,0,0,80,0,108,0,183,0,0,0,51,0,94,0,0,0,153,0,136,0,26,0,40,0,93,0,175,0,88,0,105,0,105,0,198,0,170,0,48,0,213,0,52,0,0,0,0,0,122,0,0,0,226,0,0,0,198,0,0,0,161,0,221,0,23,0,240,0,252,0,94,0,116,0,27,0,0,0,247,0,55,0,66,0,23,0,132,0,236,0,249,0,119,0,0,0,229,0,245,0,0,0,238,0,166,0,249,0,62,0,66,0,0,0,0,0,35,0,58,0,0,0,28,0,118,0,222,0,235,0,214,0,91,0,252,0,180,0,13,0,66,0,148,0,13,0,199,0,180,0,33,0,27,0,108,0,140,0,168,0,123,0,0,0,241,0,157,0,25,0,225,0,0,0,11,0,95,0,21,0,119,0,118,0,151,0,42,0,38,0,0,0,0,0,184,0,69,0,0,0,10,0,46,0,166,0,0,0,183,0,28,0,0,0,19,0,33,0,248,0,0,0,21,0,216,0,0,0,199,0,4,0,0,0,84,0,158,0,61,0,127,0,0,0,113,0,86,0,66,0,111,0,33,0,0,0,0,0,132,0,0,0,98,0,35,0,170,0,0,0,209,0,0,0,110,0,0,0,187,0,0,0,92,0,0,0,0,0,77,0,65,0,0,0,18,0,29,0,87,0,210,0,100,0,75,0,65,0,156,0,0,0,192,0,202,0,242,0,0,0,73,0,0,0,226,0,155,0,11,0,198,0,0,0,33,0,221,0,122,0,0,0,0,0,72,0,2,0,0,0,47,0,59,0,43,0,59,0,186,0,47,0,211,0,181,0,0,0,0,0,23,0,128,0,1,0,0,0,0,0,29,0,127,0,0,0,4,0,73,0,168,0,137,0,97,0,81,0,0,0,19,0,0,0,154,0,164,0,121,0,176,0,198,0,69,0,0,0,150,0,239,0,109,0,180,0,53,0,221,0,0,0,19,0,59,0,88,0,215,0,0,0,221,0,87,0,129,0,143,0,242,0,84,0,113,0,212,0,117,0,92,0,183,0,128,0,124,0,130,0,140,0,252,0,47,0,10,0,59,0,101,0,109,0,224,0,0,0,0,0,252,0,225,0,85,0,201,0,75,0,0,0,215,0,188,0,0,0,136,0,97,0,163,0,55,0,212,0,150,0,0,0,215,0,145,0,18,0,148,0,121,0,25,0,53,0,159,0,205,0,58,0,0,0,0,0,0,0,39,0,57,0,0,0,219,0,0,0,94,0,33,0,0,0,194,0,119,0,255,0,194,0,142,0,0,0,77,0,83,0,205,0,0,0,42,0,247,0,179,0,0,0,141,0,192,0,0,0,141,0,132,0,189,0,144,0,115,0,0,0,134,0,94,0,52,0,56,0,12,0,0,0,9,0,0,0,132,0,21,0,89,0,33,0,18,0,183,0,104,0,23,0,214,0,57,0,101,0,64,0,135,0,221,0,64,0,0,0,255,0,29,0,0,0,213,0,141,0,183,0,147,0,111,0,221,0,0,0,187,0,15,0,78,0,188,0,199,0,47,0,224,0,253,0,198,0,49,0,0,0,234,0,176,0,211,0,79,0,131,0,234,0,0,0,253,0,31,0,0,0,0,0,250,0,229,0,200,0,97,0,129,0,21,0,108,0,124,0,69,0,72,0,45,0,66,0,194,0,183,0,0,0,37,0,21,0,0,0,0,0,220,0,225,0,2,0,221,0,42,0,75,0,186,0,13,0,131,0,18,0,84,0,95,0,0,0,218,0,0,0,0,0,230,0,0,0,104,0,211,0,169,0,238,0,63,0,42,0,8,0,26,0,183,0,172,0,0,0,219,0,82,0,45,0,0,0,212,0,206,0,114,0,101,0,0,0,249,0,94,0,0,0,0,0,0,0,0,0,0,0,0,0,221,0,59,0,25,0,199,0,9,0,102,0,175,0,132,0,179,0,128,0,18,0,0,0,49,0,123,0,188,0,0,0,108,0,0,0,249,0,51,0,197,0,65,0,100,0,0,0,86,0,53,0,0,0,218,0,78,0,59,0,30,0,0,0,100,0,231,0,110,0,0,0,0,0,0,0,0,0,0,0,252,0,0,0,212,0,45,0,163,0,149,0,49,0,0,0,128,0,126,0,155,0,41,0,177,0,129,0,0,0,217,0,0,0,135,0,235,0,246,0,8,0,101,0,215,0,0,0,159,0,108,0,99,0,121,0,130,0,233,0,72,0,0,0,113,0,0,0,192,0,42,0,157,0,160,0,191,0,122,0,63,0,0,0,52,0,27,0,110,0,211,0,0,0,11,0,68,0,196,0,210,0,62,0,0,0,168,0,201,0,252,0,174,0,178,0,91,0,244,0,108,0,90,0,0,0,171,0,0,0,33,0,88,0,143,0,66,0,50,0,0,0,217,0,224,0,193,0,23,0,221,0,0,0,0,0,0,0,169,0,168,0,248,0,0,0,167,0,59,0,41,0,225,0,106,0,77,0,159,0,203,0,0,0,252,0,134,0,0,0,243,0,160,0,0,0,0,0,193,0,0,0,6,0,160,0,164,0,147,0,0,0,103,0,140,0,93,0,126,0,0,0,20,0,146,0,254,0,0,0,212,0,176,0,45,0,84,0,222,0,250,0,74,0,222,0,152,0,100,0,6,0,150,0,0,0,0,0,3,0,106,0,114,0,241,0,241,0,35,0,176,0,0,0,70,0,239,0,249,0,160,0,19,0,12,0,68,0,20,0,75,0,0,0,105,0,0,0,63,0,200,0,201,0,0,0,193,0,231,0,138,0,230,0,240,0,15,0,235,0,90,0,183,0,166,0,216,0,228,0,255,0,200,0,156,0,201,0,0,0,249,0,38,0,108,0,82,0,113,0,96,0,35,0,123,0,1,0,0,0,32,0,208,0,0,0,28,0,167,0,11,0,148,0,161,0,8,0,0,0,12,0,225,0,1,0,139,0,94,0,79,0,177,0,38,0,0,0,128,0,56,0,91,0,0,0,100,0,89,0,194,0,194,0,13,0,161,0,219,0,81,0,106,0,84,0,69,0,0,0,26,0,96,0,138,0,52,0,0,0,26,0,211,0,133,0,44,0,114,0,209,0,244,0,69,0,134,0,68,0,197,0,114,0,187,0,92,0,239,0,130,0,0,0,171,0,250,0,61,0,118,0,233,0,78,0,84,0,0,0,0,0,4,0,9,0,81,0,43,0,87,0,243,0,0,0,233,0,101,0,212,0,0,0,230,0,188,0,63,0,0,0,58,0,0,0,195,0,199,0,10,0,105,0,0,0,14,0,123,0,254,0,0,0,237,0,89,0,246,0,16,0,0,0,67,0,73,0,0,0,70,0,245,0,69,0,96,0,221,0,241,0,0,0,13,0,31,0,194,0,50,0,141,0,244,0,103,0,204,0,0,0,0,0,0,0,0,0,172,0,241,0,0,0,0,0,219,0,225,0,103,0,254,0,103,0,197,0,232,0,138,0,181,0,119,0,38,0,141,0,65,0,0,0,12,0,34,0,22,0,175,0,73,0,8,0,58,0,155,0,171,0,250,0,90,0,35,0,154,0,0,0,90,0,41,0,0,0,126,0,178,0,181,0,25,0,232,0,0,0,181,0,78,0,241,0,32,0,105,0,221,0,49,0,28,0,143,0,95,0,110,0,250,0,45,0,250,0,47,0,0,0,204,0,127,0,169,0,191,0,35,0,51,0,176,0,0,0,78,0,153,0,207,0,199,0,130,0,148,0,255,0,8,0,200,0,190,0,190,0,77,0,144,0,87,0,65,0,210,0,70,0,52,0,95,0,185,0,203,0,126,0,136,0,45,0);
signal scenario_full  : scenario_type := (0,0,22,31,22,30,22,29,62,31,102,31,102,30,133,31,180,31,180,30,45,31,204,31,244,31,155,31,209,31,166,31,166,30,70,31,70,30,70,29,8,31,221,31,19,31,178,31,187,31,8,31,64,31,8,31,42,31,42,30,70,31,180,31,124,31,39,31,39,30,78,31,129,31,179,31,22,31,176,31,176,30,218,31,218,30,121,31,54,31,57,31,35,31,35,30,112,31,56,31,115,31,168,31,44,31,146,31,198,31,52,31,132,31,236,31,21,31,66,31,134,31,23,31,23,30,129,31,160,31,245,31,100,31,100,30,96,31,96,30,189,31,89,31,82,31,153,31,123,31,123,30,162,31,162,30,107,31,206,31,48,31,254,31,221,31,129,31,114,31,9,31,2,31,185,31,162,31,19,31,151,31,151,30,151,29,217,31,80,31,14,31,11,31,232,31,226,31,34,31,63,31,84,31,34,31,135,31,108,31,73,31,73,30,169,31,118,31,118,30,118,29,118,28,118,27,177,31,22,31,14,31,114,31,253,31,223,31,9,31,243,31,14,31,137,31,137,30,211,31,211,30,164,31,93,31,222,31,137,31,142,31,210,31,137,31,240,31,152,31,239,31,235,31,235,30,41,31,89,31,7,31,166,31,194,31,194,30,170,31,64,31,163,31,163,30,136,31,136,30,136,29,181,31,78,31,238,31,238,30,238,29,1,31,12,31,188,31,236,31,129,31,31,31,82,31,82,30,53,31,251,31,251,30,80,31,108,31,183,31,183,30,51,31,94,31,94,30,153,31,136,31,26,31,40,31,93,31,175,31,88,31,105,31,105,31,198,31,170,31,48,31,213,31,52,31,52,30,52,29,122,31,122,30,226,31,226,30,198,31,198,30,161,31,221,31,23,31,240,31,252,31,94,31,116,31,27,31,27,30,247,31,55,31,66,31,23,31,132,31,236,31,249,31,119,31,119,30,229,31,245,31,245,30,238,31,166,31,249,31,62,31,66,31,66,30,66,29,35,31,58,31,58,30,28,31,118,31,222,31,235,31,214,31,91,31,252,31,180,31,13,31,66,31,148,31,13,31,199,31,180,31,33,31,27,31,108,31,140,31,168,31,123,31,123,30,241,31,157,31,25,31,225,31,225,30,11,31,95,31,21,31,119,31,118,31,151,31,42,31,38,31,38,30,38,29,184,31,69,31,69,30,10,31,46,31,166,31,166,30,183,31,28,31,28,30,19,31,33,31,248,31,248,30,21,31,216,31,216,30,199,31,4,31,4,30,84,31,158,31,61,31,127,31,127,30,113,31,86,31,66,31,111,31,33,31,33,30,33,29,132,31,132,30,98,31,35,31,170,31,170,30,209,31,209,30,110,31,110,30,187,31,187,30,92,31,92,30,92,29,77,31,65,31,65,30,18,31,29,31,87,31,210,31,100,31,75,31,65,31,156,31,156,30,192,31,202,31,242,31,242,30,73,31,73,30,226,31,155,31,11,31,198,31,198,30,33,31,221,31,122,31,122,30,122,29,72,31,2,31,2,30,47,31,59,31,43,31,59,31,186,31,47,31,211,31,181,31,181,30,181,29,23,31,128,31,1,31,1,30,1,29,29,31,127,31,127,30,4,31,73,31,168,31,137,31,97,31,81,31,81,30,19,31,19,30,154,31,164,31,121,31,176,31,198,31,69,31,69,30,150,31,239,31,109,31,180,31,53,31,221,31,221,30,19,31,59,31,88,31,215,31,215,30,221,31,87,31,129,31,143,31,242,31,84,31,113,31,212,31,117,31,92,31,183,31,128,31,124,31,130,31,140,31,252,31,47,31,10,31,59,31,101,31,109,31,224,31,224,30,224,29,252,31,225,31,85,31,201,31,75,31,75,30,215,31,188,31,188,30,136,31,97,31,163,31,55,31,212,31,150,31,150,30,215,31,145,31,18,31,148,31,121,31,25,31,53,31,159,31,205,31,58,31,58,30,58,29,58,28,39,31,57,31,57,30,219,31,219,30,94,31,33,31,33,30,194,31,119,31,255,31,194,31,142,31,142,30,77,31,83,31,205,31,205,30,42,31,247,31,179,31,179,30,141,31,192,31,192,30,141,31,132,31,189,31,144,31,115,31,115,30,134,31,94,31,52,31,56,31,12,31,12,30,9,31,9,30,132,31,21,31,89,31,33,31,18,31,183,31,104,31,23,31,214,31,57,31,101,31,64,31,135,31,221,31,64,31,64,30,255,31,29,31,29,30,213,31,141,31,183,31,147,31,111,31,221,31,221,30,187,31,15,31,78,31,188,31,199,31,47,31,224,31,253,31,198,31,49,31,49,30,234,31,176,31,211,31,79,31,131,31,234,31,234,30,253,31,31,31,31,30,31,29,250,31,229,31,200,31,97,31,129,31,21,31,108,31,124,31,69,31,72,31,45,31,66,31,194,31,183,31,183,30,37,31,21,31,21,30,21,29,220,31,225,31,2,31,221,31,42,31,75,31,186,31,13,31,131,31,18,31,84,31,95,31,95,30,218,31,218,30,218,29,230,31,230,30,104,31,211,31,169,31,238,31,63,31,42,31,8,31,26,31,183,31,172,31,172,30,219,31,82,31,45,31,45,30,212,31,206,31,114,31,101,31,101,30,249,31,94,31,94,30,94,29,94,28,94,27,94,26,94,25,221,31,59,31,25,31,199,31,9,31,102,31,175,31,132,31,179,31,128,31,18,31,18,30,49,31,123,31,188,31,188,30,108,31,108,30,249,31,51,31,197,31,65,31,100,31,100,30,86,31,53,31,53,30,218,31,78,31,59,31,30,31,30,30,100,31,231,31,110,31,110,30,110,29,110,28,110,27,110,26,252,31,252,30,212,31,45,31,163,31,149,31,49,31,49,30,128,31,126,31,155,31,41,31,177,31,129,31,129,30,217,31,217,30,135,31,235,31,246,31,8,31,101,31,215,31,215,30,159,31,108,31,99,31,121,31,130,31,233,31,72,31,72,30,113,31,113,30,192,31,42,31,157,31,160,31,191,31,122,31,63,31,63,30,52,31,27,31,110,31,211,31,211,30,11,31,68,31,196,31,210,31,62,31,62,30,168,31,201,31,252,31,174,31,178,31,91,31,244,31,108,31,90,31,90,30,171,31,171,30,33,31,88,31,143,31,66,31,50,31,50,30,217,31,224,31,193,31,23,31,221,31,221,30,221,29,221,28,169,31,168,31,248,31,248,30,167,31,59,31,41,31,225,31,106,31,77,31,159,31,203,31,203,30,252,31,134,31,134,30,243,31,160,31,160,30,160,29,193,31,193,30,6,31,160,31,164,31,147,31,147,30,103,31,140,31,93,31,126,31,126,30,20,31,146,31,254,31,254,30,212,31,176,31,45,31,84,31,222,31,250,31,74,31,222,31,152,31,100,31,6,31,150,31,150,30,150,29,3,31,106,31,114,31,241,31,241,31,35,31,176,31,176,30,70,31,239,31,249,31,160,31,19,31,12,31,68,31,20,31,75,31,75,30,105,31,105,30,63,31,200,31,201,31,201,30,193,31,231,31,138,31,230,31,240,31,15,31,235,31,90,31,183,31,166,31,216,31,228,31,255,31,200,31,156,31,201,31,201,30,249,31,38,31,108,31,82,31,113,31,96,31,35,31,123,31,1,31,1,30,32,31,208,31,208,30,28,31,167,31,11,31,148,31,161,31,8,31,8,30,12,31,225,31,1,31,139,31,94,31,79,31,177,31,38,31,38,30,128,31,56,31,91,31,91,30,100,31,89,31,194,31,194,31,13,31,161,31,219,31,81,31,106,31,84,31,69,31,69,30,26,31,96,31,138,31,52,31,52,30,26,31,211,31,133,31,44,31,114,31,209,31,244,31,69,31,134,31,68,31,197,31,114,31,187,31,92,31,239,31,130,31,130,30,171,31,250,31,61,31,118,31,233,31,78,31,84,31,84,30,84,29,4,31,9,31,81,31,43,31,87,31,243,31,243,30,233,31,101,31,212,31,212,30,230,31,188,31,63,31,63,30,58,31,58,30,195,31,199,31,10,31,105,31,105,30,14,31,123,31,254,31,254,30,237,31,89,31,246,31,16,31,16,30,67,31,73,31,73,30,70,31,245,31,69,31,96,31,221,31,241,31,241,30,13,31,31,31,194,31,50,31,141,31,244,31,103,31,204,31,204,30,204,29,204,28,204,27,172,31,241,31,241,30,241,29,219,31,225,31,103,31,254,31,103,31,197,31,232,31,138,31,181,31,119,31,38,31,141,31,65,31,65,30,12,31,34,31,22,31,175,31,73,31,8,31,58,31,155,31,171,31,250,31,90,31,35,31,154,31,154,30,90,31,41,31,41,30,126,31,178,31,181,31,25,31,232,31,232,30,181,31,78,31,241,31,32,31,105,31,221,31,49,31,28,31,143,31,95,31,110,31,250,31,45,31,250,31,47,31,47,30,204,31,127,31,169,31,191,31,35,31,51,31,176,31,176,30,78,31,153,31,207,31,199,31,130,31,148,31,255,31,8,31,200,31,190,31,190,31,77,31,144,31,87,31,65,31,210,31,70,31,52,31,95,31,185,31,203,31,126,31,136,31,45,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
