-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 632;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (253,0,64,0,50,0,132,0,78,0,123,0,210,0,179,0,208,0,201,0,82,0,117,0,200,0,0,0,228,0,72,0,32,0,141,0,120,0,0,0,137,0,63,0,0,0,223,0,195,0,0,0,25,0,135,0,50,0,94,0,0,0,153,0,0,0,150,0,169,0,231,0,56,0,33,0,113,0,0,0,0,0,127,0,0,0,119,0,187,0,106,0,201,0,106,0,217,0,43,0,125,0,157,0,192,0,47,0,65,0,83,0,106,0,27,0,238,0,244,0,222,0,49,0,86,0,184,0,120,0,211,0,59,0,16,0,55,0,232,0,0,0,240,0,209,0,216,0,0,0,136,0,189,0,0,0,0,0,0,0,63,0,142,0,100,0,70,0,251,0,0,0,147,0,174,0,0,0,230,0,27,0,124,0,19,0,188,0,112,0,45,0,53,0,0,0,203,0,17,0,10,0,81,0,51,0,24,0,130,0,240,0,190,0,0,0,134,0,190,0,247,0,24,0,239,0,171,0,184,0,153,0,73,0,82,0,26,0,94,0,0,0,0,0,250,0,100,0,45,0,219,0,56,0,59,0,0,0,136,0,43,0,65,0,0,0,0,0,133,0,0,0,65,0,88,0,13,0,83,0,1,0,166,0,0,0,116,0,0,0,126,0,44,0,108,0,0,0,66,0,239,0,100,0,0,0,29,0,69,0,0,0,83,0,0,0,47,0,0,0,245,0,241,0,41,0,64,0,212,0,102,0,42,0,174,0,39,0,50,0,235,0,0,0,78,0,179,0,77,0,6,0,0,0,154,0,86,0,0,0,0,0,249,0,135,0,82,0,0,0,9,0,32,0,253,0,200,0,117,0,65,0,139,0,0,0,0,0,0,0,243,0,63,0,64,0,0,0,242,0,124,0,208,0,89,0,141,0,0,0,148,0,0,0,241,0,58,0,23,0,15,0,37,0,113,0,243,0,112,0,246,0,59,0,247,0,107,0,79,0,25,0,7,0,169,0,206,0,234,0,252,0,97,0,0,0,103,0,197,0,255,0,153,0,0,0,187,0,53,0,233,0,227,0,0,0,255,0,110,0,120,0,58,0,141,0,137,0,251,0,155,0,0,0,173,0,141,0,221,0,165,0,105,0,0,0,54,0,238,0,16,0,128,0,242,0,96,0,0,0,57,0,0,0,0,0,0,0,0,0,205,0,244,0,212,0,218,0,0,0,218,0,53,0,164,0,0,0,12,0,145,0,100,0,71,0,158,0,0,0,169,0,26,0,226,0,80,0,88,0,63,0,232,0,69,0,98,0,97,0,219,0,255,0,0,0,0,0,56,0,226,0,237,0,56,0,87,0,101,0,222,0,112,0,225,0,168,0,102,0,102,0,64,0,169,0,226,0,232,0,45,0,69,0,0,0,150,0,241,0,235,0,85,0,125,0,129,0,0,0,0,0,0,0,217,0,24,0,156,0,0,0,51,0,13,0,28,0,49,0,246,0,153,0,0,0,146,0,0,0,0,0,151,0,210,0,147,0,190,0,58,0,215,0,0,0,252,0,201,0,61,0,19,0,115,0,115,0,0,0,0,0,91,0,197,0,188,0,94,0,35,0,165,0,136,0,2,0,0,0,94,0,0,0,0,0,246,0,171,0,70,0,128,0,28,0,0,0,124,0,45,0,97,0,152,0,116,0,216,0,159,0,206,0,0,0,107,0,63,0,177,0,116,0,95,0,209,0,149,0,0,0,59,0,41,0,116,0,3,0,72,0,2,0,194,0,200,0,148,0,208,0,0,0,43,0,9,0,0,0,127,0,78,0,16,0,121,0,57,0,194,0,0,0,206,0,28,0,197,0,51,0,100,0,70,0,178,0,193,0,73,0,0,0,0,0,42,0,92,0,104,0,125,0,0,0,51,0,0,0,0,0,195,0,148,0,182,0,0,0,65,0,0,0,28,0,139,0,0,0,41,0,0,0,169,0,147,0,197,0,0,0,208,0,0,0,213,0,44,0,140,0,34,0,0,0,0,0,31,0,248,0,172,0,143,0,128,0,81,0,153,0,71,0,116,0,0,0,0,0,247,0,130,0,207,0,0,0,0,0,253,0,135,0,181,0,201,0,26,0,107,0,173,0,177,0,142,0,102,0,0,0,14,0,40,0,246,0,211,0,115,0,167,0,0,0,29,0,19,0,94,0,25,0,182,0,125,0,150,0,0,0,108,0,189,0,226,0,230,0,0,0,168,0,0,0,0,0,49,0,108,0,224,0,85,0,240,0,145,0,0,0,31,0,131,0,86,0,0,0,16,0,9,0,234,0,245,0,202,0,246,0,140,0,47,0,227,0,41,0,144,0,248,0,72,0,68,0,200,0,0,0,15,0,193,0,0,0,149,0,158,0,77,0,0,0,0,0,131,0,86,0,199,0,238,0,78,0,11,0,249,0,197,0,37,0,171,0,59,0,45,0,244,0,103,0,101,0,0,0,0,0,22,0,201,0,0,0,149,0,0,0,122,0,246,0,160,0,224,0,15,0,133,0,0,0,2,0,0,0,0,0,238,0,121,0,0,0,11,0,190,0,236,0,131,0,192,0,239,0,188,0,50,0,14,0,197,0,234,0,0,0,198,0,195,0,16,0,140,0,44,0,96,0,82,0,220,0,56,0,112,0,30,0,0,0,92,0,0,0,0,0,12,0,0,0,0,0,62,0,201,0,13,0,153,0,10,0,31,0,90,0,78,0,0,0,88,0,68,0,46,0,83,0,220,0,66,0,24,0,245,0,175,0,0,0,0,0,254,0,249,0,21,0,206,0,253,0,54,0,0,0,157,0,78,0,0,0,98,0,12,0,87,0);
signal scenario_full  : scenario_type := (253,31,64,31,50,31,132,31,78,31,123,31,210,31,179,31,208,31,201,31,82,31,117,31,200,31,200,30,228,31,72,31,32,31,141,31,120,31,120,30,137,31,63,31,63,30,223,31,195,31,195,30,25,31,135,31,50,31,94,31,94,30,153,31,153,30,150,31,169,31,231,31,56,31,33,31,113,31,113,30,113,29,127,31,127,30,119,31,187,31,106,31,201,31,106,31,217,31,43,31,125,31,157,31,192,31,47,31,65,31,83,31,106,31,27,31,238,31,244,31,222,31,49,31,86,31,184,31,120,31,211,31,59,31,16,31,55,31,232,31,232,30,240,31,209,31,216,31,216,30,136,31,189,31,189,30,189,29,189,28,63,31,142,31,100,31,70,31,251,31,251,30,147,31,174,31,174,30,230,31,27,31,124,31,19,31,188,31,112,31,45,31,53,31,53,30,203,31,17,31,10,31,81,31,51,31,24,31,130,31,240,31,190,31,190,30,134,31,190,31,247,31,24,31,239,31,171,31,184,31,153,31,73,31,82,31,26,31,94,31,94,30,94,29,250,31,100,31,45,31,219,31,56,31,59,31,59,30,136,31,43,31,65,31,65,30,65,29,133,31,133,30,65,31,88,31,13,31,83,31,1,31,166,31,166,30,116,31,116,30,126,31,44,31,108,31,108,30,66,31,239,31,100,31,100,30,29,31,69,31,69,30,83,31,83,30,47,31,47,30,245,31,241,31,41,31,64,31,212,31,102,31,42,31,174,31,39,31,50,31,235,31,235,30,78,31,179,31,77,31,6,31,6,30,154,31,86,31,86,30,86,29,249,31,135,31,82,31,82,30,9,31,32,31,253,31,200,31,117,31,65,31,139,31,139,30,139,29,139,28,243,31,63,31,64,31,64,30,242,31,124,31,208,31,89,31,141,31,141,30,148,31,148,30,241,31,58,31,23,31,15,31,37,31,113,31,243,31,112,31,246,31,59,31,247,31,107,31,79,31,25,31,7,31,169,31,206,31,234,31,252,31,97,31,97,30,103,31,197,31,255,31,153,31,153,30,187,31,53,31,233,31,227,31,227,30,255,31,110,31,120,31,58,31,141,31,137,31,251,31,155,31,155,30,173,31,141,31,221,31,165,31,105,31,105,30,54,31,238,31,16,31,128,31,242,31,96,31,96,30,57,31,57,30,57,29,57,28,57,27,205,31,244,31,212,31,218,31,218,30,218,31,53,31,164,31,164,30,12,31,145,31,100,31,71,31,158,31,158,30,169,31,26,31,226,31,80,31,88,31,63,31,232,31,69,31,98,31,97,31,219,31,255,31,255,30,255,29,56,31,226,31,237,31,56,31,87,31,101,31,222,31,112,31,225,31,168,31,102,31,102,31,64,31,169,31,226,31,232,31,45,31,69,31,69,30,150,31,241,31,235,31,85,31,125,31,129,31,129,30,129,29,129,28,217,31,24,31,156,31,156,30,51,31,13,31,28,31,49,31,246,31,153,31,153,30,146,31,146,30,146,29,151,31,210,31,147,31,190,31,58,31,215,31,215,30,252,31,201,31,61,31,19,31,115,31,115,31,115,30,115,29,91,31,197,31,188,31,94,31,35,31,165,31,136,31,2,31,2,30,94,31,94,30,94,29,246,31,171,31,70,31,128,31,28,31,28,30,124,31,45,31,97,31,152,31,116,31,216,31,159,31,206,31,206,30,107,31,63,31,177,31,116,31,95,31,209,31,149,31,149,30,59,31,41,31,116,31,3,31,72,31,2,31,194,31,200,31,148,31,208,31,208,30,43,31,9,31,9,30,127,31,78,31,16,31,121,31,57,31,194,31,194,30,206,31,28,31,197,31,51,31,100,31,70,31,178,31,193,31,73,31,73,30,73,29,42,31,92,31,104,31,125,31,125,30,51,31,51,30,51,29,195,31,148,31,182,31,182,30,65,31,65,30,28,31,139,31,139,30,41,31,41,30,169,31,147,31,197,31,197,30,208,31,208,30,213,31,44,31,140,31,34,31,34,30,34,29,31,31,248,31,172,31,143,31,128,31,81,31,153,31,71,31,116,31,116,30,116,29,247,31,130,31,207,31,207,30,207,29,253,31,135,31,181,31,201,31,26,31,107,31,173,31,177,31,142,31,102,31,102,30,14,31,40,31,246,31,211,31,115,31,167,31,167,30,29,31,19,31,94,31,25,31,182,31,125,31,150,31,150,30,108,31,189,31,226,31,230,31,230,30,168,31,168,30,168,29,49,31,108,31,224,31,85,31,240,31,145,31,145,30,31,31,131,31,86,31,86,30,16,31,9,31,234,31,245,31,202,31,246,31,140,31,47,31,227,31,41,31,144,31,248,31,72,31,68,31,200,31,200,30,15,31,193,31,193,30,149,31,158,31,77,31,77,30,77,29,131,31,86,31,199,31,238,31,78,31,11,31,249,31,197,31,37,31,171,31,59,31,45,31,244,31,103,31,101,31,101,30,101,29,22,31,201,31,201,30,149,31,149,30,122,31,246,31,160,31,224,31,15,31,133,31,133,30,2,31,2,30,2,29,238,31,121,31,121,30,11,31,190,31,236,31,131,31,192,31,239,31,188,31,50,31,14,31,197,31,234,31,234,30,198,31,195,31,16,31,140,31,44,31,96,31,82,31,220,31,56,31,112,31,30,31,30,30,92,31,92,30,92,29,12,31,12,30,12,29,62,31,201,31,13,31,153,31,10,31,31,31,90,31,78,31,78,30,88,31,68,31,46,31,83,31,220,31,66,31,24,31,245,31,175,31,175,30,175,29,254,31,249,31,21,31,206,31,253,31,54,31,54,30,157,31,78,31,78,30,98,31,12,31,87,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
