-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 689;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (212,0,102,0,121,0,75,0,69,0,61,0,238,0,22,0,82,0,0,0,164,0,0,0,59,0,151,0,221,0,198,0,183,0,44,0,165,0,193,0,99,0,64,0,0,0,172,0,0,0,0,0,247,0,154,0,237,0,156,0,0,0,14,0,157,0,139,0,226,0,0,0,18,0,0,0,224,0,49,0,0,0,0,0,45,0,153,0,0,0,222,0,91,0,0,0,220,0,116,0,34,0,180,0,151,0,22,0,195,0,53,0,179,0,90,0,50,0,0,0,109,0,189,0,238,0,112,0,23,0,253,0,0,0,224,0,121,0,161,0,149,0,0,0,244,0,0,0,169,0,0,0,48,0,29,0,10,0,110,0,60,0,0,0,0,0,152,0,155,0,191,0,203,0,245,0,0,0,61,0,0,0,126,0,202,0,115,0,164,0,224,0,73,0,252,0,232,0,117,0,50,0,195,0,160,0,97,0,97,0,0,0,248,0,14,0,0,0,243,0,160,0,144,0,145,0,161,0,0,0,0,0,142,0,31,0,141,0,238,0,3,0,177,0,133,0,36,0,80,0,0,0,214,0,30,0,136,0,247,0,191,0,0,0,86,0,241,0,18,0,196,0,57,0,0,0,138,0,52,0,0,0,86,0,68,0,84,0,0,0,55,0,231,0,0,0,0,0,143,0,0,0,187,0,195,0,150,0,0,0,167,0,253,0,0,0,65,0,101,0,0,0,52,0,80,0,213,0,0,0,0,0,0,0,109,0,96,0,13,0,135,0,63,0,228,0,5,0,229,0,0,0,16,0,103,0,196,0,206,0,208,0,231,0,209,0,123,0,0,0,0,0,0,0,0,0,168,0,83,0,71,0,69,0,1,0,11,0,137,0,0,0,77,0,236,0,33,0,247,0,11,0,37,0,202,0,0,0,77,0,198,0,185,0,186,0,254,0,144,0,45,0,0,0,0,0,62,0,0,0,220,0,206,0,207,0,214,0,92,0,171,0,43,0,173,0,150,0,229,0,65,0,0,0,238,0,158,0,160,0,50,0,149,0,120,0,65,0,189,0,0,0,0,0,179,0,192,0,138,0,135,0,34,0,78,0,93,0,136,0,134,0,45,0,228,0,38,0,185,0,128,0,122,0,233,0,21,0,0,0,119,0,0,0,0,0,163,0,79,0,212,0,2,0,0,0,84,0,200,0,153,0,125,0,191,0,0,0,0,0,95,0,189,0,30,0,202,0,67,0,214,0,0,0,28,0,44,0,218,0,41,0,0,0,119,0,154,0,30,0,98,0,0,0,0,0,134,0,88,0,117,0,68,0,104,0,192,0,0,0,0,0,50,0,0,0,234,0,0,0,79,0,0,0,0,0,0,0,86,0,226,0,0,0,129,0,0,0,112,0,253,0,0,0,237,0,127,0,150,0,0,0,46,0,82,0,147,0,79,0,175,0,200,0,30,0,0,0,133,0,209,0,51,0,249,0,62,0,250,0,221,0,104,0,132,0,242,0,61,0,126,0,45,0,0,0,211,0,0,0,52,0,0,0,14,0,11,0,143,0,38,0,68,0,59,0,217,0,0,0,0,0,136,0,149,0,137,0,0,0,166,0,103,0,48,0,1,0,12,0,129,0,0,0,253,0,250,0,150,0,227,0,0,0,0,0,252,0,200,0,203,0,183,0,0,0,180,0,0,0,247,0,0,0,121,0,84,0,3,0,142,0,53,0,228,0,15,0,176,0,98,0,175,0,71,0,109,0,111,0,0,0,177,0,237,0,106,0,228,0,92,0,127,0,0,0,37,0,45,0,69,0,196,0,21,0,237,0,0,0,186,0,64,0,76,0,250,0,78,0,25,0,218,0,123,0,89,0,209,0,206,0,89,0,5,0,94,0,142,0,42,0,177,0,42,0,176,0,202,0,156,0,27,0,64,0,0,0,17,0,0,0,195,0,228,0,0,0,32,0,187,0,232,0,37,0,0,0,132,0,25,0,158,0,83,0,143,0,175,0,0,0,194,0,142,0,94,0,0,0,0,0,200,0,0,0,78,0,73,0,18,0,22,0,0,0,97,0,0,0,113,0,253,0,151,0,83,0,0,0,114,0,254,0,127,0,89,0,135,0,0,0,247,0,0,0,0,0,170,0,27,0,108,0,103,0,34,0,156,0,225,0,166,0,205,0,20,0,168,0,215,0,85,0,213,0,237,0,0,0,34,0,0,0,0,0,126,0,175,0,0,0,69,0,157,0,243,0,5,0,59,0,110,0,61,0,42,0,198,0,67,0,0,0,24,0,46,0,51,0,0,0,93,0,86,0,233,0,209,0,127,0,47,0,148,0,116,0,192,0,225,0,0,0,56,0,0,0,164,0,222,0,87,0,128,0,27,0,0,0,24,0,193,0,214,0,222,0,44,0,180,0,0,0,246,0,0,0,98,0,0,0,58,0,65,0,16,0,0,0,0,0,233,0,253,0,110,0,92,0,128,0,58,0,42,0,165,0,0,0,0,0,8,0,56,0,201,0,222,0,146,0,239,0,242,0,43,0,121,0,30,0,0,0,47,0,0,0,130,0,64,0,112,0,168,0,244,0,143,0,124,0,153,0,200,0,0,0,186,0,79,0,77,0,225,0,216,0,218,0,39,0,84,0,202,0,0,0,151,0,184,0,90,0,210,0,0,0,126,0,242,0,88,0,0,0,103,0,30,0,113,0,0,0,0,0,25,0,0,0,250,0,20,0,130,0,0,0,197,0,167,0,94,0,58,0,156,0,6,0,0,0,209,0,81,0,224,0,39,0,241,0,90,0,0,0,212,0,165,0,18,0,195,0,0,0,0,0,148,0,69,0,57,0,202,0,143,0,175,0,30,0,24,0,105,0,0,0,218,0,179,0,20,0,104,0,83,0,205,0,63,0,104,0,106,0,139,0,0,0,200,0,0,0,243,0,117,0,0,0,10,0,255,0,202,0,148,0,219,0,110,0,230,0,123,0,149,0,252,0,180,0,57,0,40,0,43,0,111,0,0,0,218,0,9,0,74,0,75,0,0,0,0,0,172,0,53,0,225,0,253,0,184,0,141,0,249,0,0,0,16,0,0,0,245,0,159,0);
signal scenario_full  : scenario_type := (212,31,102,31,121,31,75,31,69,31,61,31,238,31,22,31,82,31,82,30,164,31,164,30,59,31,151,31,221,31,198,31,183,31,44,31,165,31,193,31,99,31,64,31,64,30,172,31,172,30,172,29,247,31,154,31,237,31,156,31,156,30,14,31,157,31,139,31,226,31,226,30,18,31,18,30,224,31,49,31,49,30,49,29,45,31,153,31,153,30,222,31,91,31,91,30,220,31,116,31,34,31,180,31,151,31,22,31,195,31,53,31,179,31,90,31,50,31,50,30,109,31,189,31,238,31,112,31,23,31,253,31,253,30,224,31,121,31,161,31,149,31,149,30,244,31,244,30,169,31,169,30,48,31,29,31,10,31,110,31,60,31,60,30,60,29,152,31,155,31,191,31,203,31,245,31,245,30,61,31,61,30,126,31,202,31,115,31,164,31,224,31,73,31,252,31,232,31,117,31,50,31,195,31,160,31,97,31,97,31,97,30,248,31,14,31,14,30,243,31,160,31,144,31,145,31,161,31,161,30,161,29,142,31,31,31,141,31,238,31,3,31,177,31,133,31,36,31,80,31,80,30,214,31,30,31,136,31,247,31,191,31,191,30,86,31,241,31,18,31,196,31,57,31,57,30,138,31,52,31,52,30,86,31,68,31,84,31,84,30,55,31,231,31,231,30,231,29,143,31,143,30,187,31,195,31,150,31,150,30,167,31,253,31,253,30,65,31,101,31,101,30,52,31,80,31,213,31,213,30,213,29,213,28,109,31,96,31,13,31,135,31,63,31,228,31,5,31,229,31,229,30,16,31,103,31,196,31,206,31,208,31,231,31,209,31,123,31,123,30,123,29,123,28,123,27,168,31,83,31,71,31,69,31,1,31,11,31,137,31,137,30,77,31,236,31,33,31,247,31,11,31,37,31,202,31,202,30,77,31,198,31,185,31,186,31,254,31,144,31,45,31,45,30,45,29,62,31,62,30,220,31,206,31,207,31,214,31,92,31,171,31,43,31,173,31,150,31,229,31,65,31,65,30,238,31,158,31,160,31,50,31,149,31,120,31,65,31,189,31,189,30,189,29,179,31,192,31,138,31,135,31,34,31,78,31,93,31,136,31,134,31,45,31,228,31,38,31,185,31,128,31,122,31,233,31,21,31,21,30,119,31,119,30,119,29,163,31,79,31,212,31,2,31,2,30,84,31,200,31,153,31,125,31,191,31,191,30,191,29,95,31,189,31,30,31,202,31,67,31,214,31,214,30,28,31,44,31,218,31,41,31,41,30,119,31,154,31,30,31,98,31,98,30,98,29,134,31,88,31,117,31,68,31,104,31,192,31,192,30,192,29,50,31,50,30,234,31,234,30,79,31,79,30,79,29,79,28,86,31,226,31,226,30,129,31,129,30,112,31,253,31,253,30,237,31,127,31,150,31,150,30,46,31,82,31,147,31,79,31,175,31,200,31,30,31,30,30,133,31,209,31,51,31,249,31,62,31,250,31,221,31,104,31,132,31,242,31,61,31,126,31,45,31,45,30,211,31,211,30,52,31,52,30,14,31,11,31,143,31,38,31,68,31,59,31,217,31,217,30,217,29,136,31,149,31,137,31,137,30,166,31,103,31,48,31,1,31,12,31,129,31,129,30,253,31,250,31,150,31,227,31,227,30,227,29,252,31,200,31,203,31,183,31,183,30,180,31,180,30,247,31,247,30,121,31,84,31,3,31,142,31,53,31,228,31,15,31,176,31,98,31,175,31,71,31,109,31,111,31,111,30,177,31,237,31,106,31,228,31,92,31,127,31,127,30,37,31,45,31,69,31,196,31,21,31,237,31,237,30,186,31,64,31,76,31,250,31,78,31,25,31,218,31,123,31,89,31,209,31,206,31,89,31,5,31,94,31,142,31,42,31,177,31,42,31,176,31,202,31,156,31,27,31,64,31,64,30,17,31,17,30,195,31,228,31,228,30,32,31,187,31,232,31,37,31,37,30,132,31,25,31,158,31,83,31,143,31,175,31,175,30,194,31,142,31,94,31,94,30,94,29,200,31,200,30,78,31,73,31,18,31,22,31,22,30,97,31,97,30,113,31,253,31,151,31,83,31,83,30,114,31,254,31,127,31,89,31,135,31,135,30,247,31,247,30,247,29,170,31,27,31,108,31,103,31,34,31,156,31,225,31,166,31,205,31,20,31,168,31,215,31,85,31,213,31,237,31,237,30,34,31,34,30,34,29,126,31,175,31,175,30,69,31,157,31,243,31,5,31,59,31,110,31,61,31,42,31,198,31,67,31,67,30,24,31,46,31,51,31,51,30,93,31,86,31,233,31,209,31,127,31,47,31,148,31,116,31,192,31,225,31,225,30,56,31,56,30,164,31,222,31,87,31,128,31,27,31,27,30,24,31,193,31,214,31,222,31,44,31,180,31,180,30,246,31,246,30,98,31,98,30,58,31,65,31,16,31,16,30,16,29,233,31,253,31,110,31,92,31,128,31,58,31,42,31,165,31,165,30,165,29,8,31,56,31,201,31,222,31,146,31,239,31,242,31,43,31,121,31,30,31,30,30,47,31,47,30,130,31,64,31,112,31,168,31,244,31,143,31,124,31,153,31,200,31,200,30,186,31,79,31,77,31,225,31,216,31,218,31,39,31,84,31,202,31,202,30,151,31,184,31,90,31,210,31,210,30,126,31,242,31,88,31,88,30,103,31,30,31,113,31,113,30,113,29,25,31,25,30,250,31,20,31,130,31,130,30,197,31,167,31,94,31,58,31,156,31,6,31,6,30,209,31,81,31,224,31,39,31,241,31,90,31,90,30,212,31,165,31,18,31,195,31,195,30,195,29,148,31,69,31,57,31,202,31,143,31,175,31,30,31,24,31,105,31,105,30,218,31,179,31,20,31,104,31,83,31,205,31,63,31,104,31,106,31,139,31,139,30,200,31,200,30,243,31,117,31,117,30,10,31,255,31,202,31,148,31,219,31,110,31,230,31,123,31,149,31,252,31,180,31,57,31,40,31,43,31,111,31,111,30,218,31,9,31,74,31,75,31,75,30,75,29,172,31,53,31,225,31,253,31,184,31,141,31,249,31,249,30,16,31,16,30,245,31,159,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
