-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 646;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (175,0,230,0,202,0,4,0,0,0,0,0,105,0,201,0,2,0,228,0,107,0,104,0,252,0,89,0,0,0,172,0,65,0,243,0,62,0,57,0,49,0,248,0,82,0,220,0,13,0,0,0,55,0,126,0,31,0,169,0,99,0,96,0,251,0,194,0,0,0,114,0,0,0,65,0,203,0,18,0,31,0,164,0,108,0,0,0,185,0,55,0,0,0,34,0,107,0,60,0,114,0,226,0,0,0,183,0,239,0,122,0,225,0,253,0,189,0,250,0,0,0,196,0,160,0,20,0,116,0,2,0,95,0,40,0,203,0,198,0,68,0,104,0,53,0,85,0,150,0,0,0,165,0,134,0,78,0,203,0,0,0,88,0,250,0,177,0,211,0,214,0,232,0,166,0,54,0,130,0,0,0,0,0,0,0,124,0,135,0,108,0,116,0,0,0,196,0,159,0,37,0,212,0,95,0,22,0,157,0,0,0,0,0,180,0,59,0,135,0,197,0,163,0,238,0,59,0,178,0,18,0,128,0,65,0,175,0,225,0,0,0,0,0,231,0,254,0,23,0,130,0,75,0,173,0,100,0,154,0,9,0,12,0,0,0,43,0,181,0,156,0,0,0,0,0,1,0,53,0,74,0,0,0,176,0,145,0,160,0,129,0,251,0,99,0,146,0,158,0,105,0,0,0,240,0,0,0,126,0,0,0,206,0,222,0,248,0,113,0,0,0,206,0,0,0,42,0,75,0,47,0,76,0,78,0,50,0,60,0,162,0,0,0,202,0,186,0,0,0,0,0,81,0,0,0,27,0,31,0,91,0,201,0,204,0,220,0,0,0,130,0,49,0,38,0,133,0,135,0,146,0,77,0,0,0,0,0,191,0,40,0,55,0,66,0,102,0,21,0,0,0,227,0,0,0,187,0,0,0,84,0,46,0,225,0,0,0,81,0,118,0,211,0,89,0,84,0,241,0,138,0,0,0,7,0,52,0,237,0,4,0,0,0,0,0,59,0,50,0,149,0,0,0,251,0,175,0,77,0,215,0,200,0,184,0,214,0,0,0,60,0,0,0,84,0,139,0,168,0,161,0,167,0,6,0,227,0,0,0,171,0,98,0,20,0,229,0,240,0,0,0,31,0,24,0,32,0,222,0,135,0,153,0,48,0,0,0,135,0,123,0,177,0,173,0,7,0,58,0,1,0,214,0,0,0,0,0,111,0,22,0,0,0,25,0,43,0,254,0,20,0,24,0,0,0,254,0,173,0,238,0,53,0,12,0,231,0,25,0,51,0,221,0,0,0,234,0,84,0,35,0,160,0,144,0,246,0,108,0,84,0,99,0,63,0,65,0,62,0,86,0,39,0,250,0,154,0,250,0,208,0,118,0,0,0,156,0,188,0,207,0,207,0,0,0,128,0,212,0,40,0,141,0,0,0,0,0,196,0,101,0,246,0,5,0,15,0,81,0,151,0,167,0,93,0,88,0,0,0,28,0,70,0,42,0,63,0,123,0,34,0,176,0,151,0,48,0,23,0,204,0,93,0,97,0,177,0,126,0,191,0,223,0,173,0,0,0,202,0,0,0,58,0,47,0,231,0,198,0,3,0,142,0,81,0,0,0,182,0,97,0,183,0,152,0,54,0,163,0,235,0,0,0,24,0,0,0,0,0,208,0,0,0,110,0,0,0,99,0,114,0,233,0,92,0,68,0,99,0,191,0,164,0,129,0,118,0,56,0,64,0,221,0,2,0,99,0,0,0,88,0,50,0,85,0,235,0,0,0,0,0,0,0,119,0,243,0,120,0,236,0,116,0,0,0,118,0,0,0,94,0,0,0,126,0,205,0,218,0,21,0,197,0,151,0,35,0,197,0,168,0,0,0,164,0,50,0,0,0,207,0,71,0,18,0,220,0,95,0,0,0,58,0,0,0,252,0,67,0,0,0,0,0,0,0,12,0,58,0,117,0,12,0,176,0,103,0,17,0,91,0,31,0,127,0,3,0,0,0,0,0,108,0,160,0,196,0,155,0,79,0,88,0,219,0,71,0,122,0,253,0,166,0,0,0,226,0,253,0,138,0,0,0,22,0,159,0,38,0,0,0,243,0,0,0,36,0,243,0,222,0,0,0,0,0,25,0,175,0,0,0,198,0,0,0,27,0,128,0,3,0,27,0,136,0,177,0,0,0,75,0,41,0,12,0,0,0,91,0,221,0,37,0,133,0,60,0,53,0,0,0,0,0,216,0,0,0,123,0,231,0,240,0,60,0,52,0,36,0,197,0,0,0,89,0,71,0,68,0,242,0,253,0,81,0,0,0,44,0,21,0,207,0,182,0,69,0,17,0,235,0,159,0,237,0,27,0,0,0,0,0,185,0,0,0,0,0,122,0,131,0,158,0,119,0,141,0,131,0,200,0,239,0,95,0,92,0,22,0,16,0,95,0,77,0,211,0,106,0,164,0,119,0,101,0,0,0,0,0,178,0,70,0,53,0,205,0,222,0,223,0,206,0,0,0,69,0,86,0,0,0,152,0,123,0,20,0,73,0,37,0,252,0,0,0,0,0,0,0,251,0,201,0,0,0,69,0,48,0,195,0,56,0,73,0,15,0,123,0,96,0,179,0,101,0,104,0,211,0,219,0,142,0,211,0,217,0,162,0,226,0,0,0,16,0,219,0,17,0,0,0,70,0,0,0,37,0,112,0,1,0,247,0,0,0,44,0,31,0,44,0,154,0,15,0,83,0,134,0,84,0,0,0,181,0,245,0,0,0,126,0,0,0,192,0,0,0,217,0,130,0,207,0,222,0,0,0,219,0,240,0,253,0,169,0,107,0,6,0,228,0,0,0,138,0,15,0,21,0,109,0,149,0,0,0,174,0,86,0,57,0,0,0,0,0,0,0,17,0,0,0);
signal scenario_full  : scenario_type := (175,31,230,31,202,31,4,31,4,30,4,29,105,31,201,31,2,31,228,31,107,31,104,31,252,31,89,31,89,30,172,31,65,31,243,31,62,31,57,31,49,31,248,31,82,31,220,31,13,31,13,30,55,31,126,31,31,31,169,31,99,31,96,31,251,31,194,31,194,30,114,31,114,30,65,31,203,31,18,31,31,31,164,31,108,31,108,30,185,31,55,31,55,30,34,31,107,31,60,31,114,31,226,31,226,30,183,31,239,31,122,31,225,31,253,31,189,31,250,31,250,30,196,31,160,31,20,31,116,31,2,31,95,31,40,31,203,31,198,31,68,31,104,31,53,31,85,31,150,31,150,30,165,31,134,31,78,31,203,31,203,30,88,31,250,31,177,31,211,31,214,31,232,31,166,31,54,31,130,31,130,30,130,29,130,28,124,31,135,31,108,31,116,31,116,30,196,31,159,31,37,31,212,31,95,31,22,31,157,31,157,30,157,29,180,31,59,31,135,31,197,31,163,31,238,31,59,31,178,31,18,31,128,31,65,31,175,31,225,31,225,30,225,29,231,31,254,31,23,31,130,31,75,31,173,31,100,31,154,31,9,31,12,31,12,30,43,31,181,31,156,31,156,30,156,29,1,31,53,31,74,31,74,30,176,31,145,31,160,31,129,31,251,31,99,31,146,31,158,31,105,31,105,30,240,31,240,30,126,31,126,30,206,31,222,31,248,31,113,31,113,30,206,31,206,30,42,31,75,31,47,31,76,31,78,31,50,31,60,31,162,31,162,30,202,31,186,31,186,30,186,29,81,31,81,30,27,31,31,31,91,31,201,31,204,31,220,31,220,30,130,31,49,31,38,31,133,31,135,31,146,31,77,31,77,30,77,29,191,31,40,31,55,31,66,31,102,31,21,31,21,30,227,31,227,30,187,31,187,30,84,31,46,31,225,31,225,30,81,31,118,31,211,31,89,31,84,31,241,31,138,31,138,30,7,31,52,31,237,31,4,31,4,30,4,29,59,31,50,31,149,31,149,30,251,31,175,31,77,31,215,31,200,31,184,31,214,31,214,30,60,31,60,30,84,31,139,31,168,31,161,31,167,31,6,31,227,31,227,30,171,31,98,31,20,31,229,31,240,31,240,30,31,31,24,31,32,31,222,31,135,31,153,31,48,31,48,30,135,31,123,31,177,31,173,31,7,31,58,31,1,31,214,31,214,30,214,29,111,31,22,31,22,30,25,31,43,31,254,31,20,31,24,31,24,30,254,31,173,31,238,31,53,31,12,31,231,31,25,31,51,31,221,31,221,30,234,31,84,31,35,31,160,31,144,31,246,31,108,31,84,31,99,31,63,31,65,31,62,31,86,31,39,31,250,31,154,31,250,31,208,31,118,31,118,30,156,31,188,31,207,31,207,31,207,30,128,31,212,31,40,31,141,31,141,30,141,29,196,31,101,31,246,31,5,31,15,31,81,31,151,31,167,31,93,31,88,31,88,30,28,31,70,31,42,31,63,31,123,31,34,31,176,31,151,31,48,31,23,31,204,31,93,31,97,31,177,31,126,31,191,31,223,31,173,31,173,30,202,31,202,30,58,31,47,31,231,31,198,31,3,31,142,31,81,31,81,30,182,31,97,31,183,31,152,31,54,31,163,31,235,31,235,30,24,31,24,30,24,29,208,31,208,30,110,31,110,30,99,31,114,31,233,31,92,31,68,31,99,31,191,31,164,31,129,31,118,31,56,31,64,31,221,31,2,31,99,31,99,30,88,31,50,31,85,31,235,31,235,30,235,29,235,28,119,31,243,31,120,31,236,31,116,31,116,30,118,31,118,30,94,31,94,30,126,31,205,31,218,31,21,31,197,31,151,31,35,31,197,31,168,31,168,30,164,31,50,31,50,30,207,31,71,31,18,31,220,31,95,31,95,30,58,31,58,30,252,31,67,31,67,30,67,29,67,28,12,31,58,31,117,31,12,31,176,31,103,31,17,31,91,31,31,31,127,31,3,31,3,30,3,29,108,31,160,31,196,31,155,31,79,31,88,31,219,31,71,31,122,31,253,31,166,31,166,30,226,31,253,31,138,31,138,30,22,31,159,31,38,31,38,30,243,31,243,30,36,31,243,31,222,31,222,30,222,29,25,31,175,31,175,30,198,31,198,30,27,31,128,31,3,31,27,31,136,31,177,31,177,30,75,31,41,31,12,31,12,30,91,31,221,31,37,31,133,31,60,31,53,31,53,30,53,29,216,31,216,30,123,31,231,31,240,31,60,31,52,31,36,31,197,31,197,30,89,31,71,31,68,31,242,31,253,31,81,31,81,30,44,31,21,31,207,31,182,31,69,31,17,31,235,31,159,31,237,31,27,31,27,30,27,29,185,31,185,30,185,29,122,31,131,31,158,31,119,31,141,31,131,31,200,31,239,31,95,31,92,31,22,31,16,31,95,31,77,31,211,31,106,31,164,31,119,31,101,31,101,30,101,29,178,31,70,31,53,31,205,31,222,31,223,31,206,31,206,30,69,31,86,31,86,30,152,31,123,31,20,31,73,31,37,31,252,31,252,30,252,29,252,28,251,31,201,31,201,30,69,31,48,31,195,31,56,31,73,31,15,31,123,31,96,31,179,31,101,31,104,31,211,31,219,31,142,31,211,31,217,31,162,31,226,31,226,30,16,31,219,31,17,31,17,30,70,31,70,30,37,31,112,31,1,31,247,31,247,30,44,31,31,31,44,31,154,31,15,31,83,31,134,31,84,31,84,30,181,31,245,31,245,30,126,31,126,30,192,31,192,30,217,31,130,31,207,31,222,31,222,30,219,31,240,31,253,31,169,31,107,31,6,31,228,31,228,30,138,31,15,31,21,31,109,31,149,31,149,30,174,31,86,31,57,31,57,30,57,29,57,28,17,31,17,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
