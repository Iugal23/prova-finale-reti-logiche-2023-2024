-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 585;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (233,0,0,0,0,0,176,0,111,0,159,0,119,0,185,0,150,0,14,0,240,0,205,0,75,0,0,0,75,0,154,0,158,0,15,0,0,0,32,0,212,0,53,0,0,0,132,0,0,0,132,0,126,0,152,0,88,0,0,0,0,0,166,0,5,0,144,0,69,0,0,0,194,0,235,0,208,0,36,0,54,0,18,0,9,0,52,0,60,0,196,0,252,0,111,0,9,0,158,0,48,0,169,0,31,0,143,0,165,0,0,0,199,0,185,0,238,0,101,0,195,0,0,0,213,0,203,0,0,0,28,0,80,0,161,0,0,0,10,0,22,0,190,0,187,0,12,0,100,0,0,0,75,0,0,0,0,0,82,0,59,0,14,0,0,0,102,0,90,0,105,0,0,0,156,0,245,0,0,0,0,0,120,0,0,0,96,0,61,0,193,0,119,0,90,0,0,0,127,0,42,0,110,0,0,0,98,0,0,0,32,0,0,0,157,0,0,0,0,0,0,0,185,0,11,0,164,0,255,0,206,0,63,0,214,0,231,0,0,0,0,0,67,0,0,0,161,0,42,0,125,0,131,0,221,0,117,0,225,0,23,0,0,0,211,0,203,0,0,0,89,0,254,0,0,0,0,0,125,0,104,0,72,0,241,0,67,0,142,0,13,0,0,0,0,0,234,0,201,0,192,0,194,0,0,0,0,0,243,0,58,0,135,0,4,0,248,0,0,0,0,0,43,0,0,0,94,0,170,0,0,0,108,0,0,0,0,0,161,0,86,0,0,0,137,0,0,0,0,0,85,0,246,0,0,0,139,0,206,0,186,0,117,0,199,0,0,0,102,0,175,0,13,0,123,0,124,0,231,0,91,0,67,0,167,0,122,0,0,0,240,0,0,0,0,0,33,0,12,0,86,0,110,0,178,0,38,0,161,0,0,0,40,0,19,0,0,0,213,0,0,0,0,0,44,0,133,0,114,0,62,0,0,0,73,0,86,0,39,0,84,0,25,0,214,0,142,0,0,0,144,0,208,0,37,0,144,0,0,0,138,0,0,0,131,0,97,0,246,0,128,0,124,0,79,0,209,0,121,0,39,0,234,0,121,0,0,0,158,0,109,0,222,0,26,0,0,0,110,0,36,0,0,0,154,0,195,0,55,0,61,0,32,0,164,0,120,0,69,0,61,0,19,0,121,0,220,0,0,0,232,0,247,0,53,0,0,0,0,0,7,0,226,0,72,0,159,0,0,0,0,0,76,0,236,0,7,0,186,0,7,0,174,0,126,0,0,0,206,0,129,0,139,0,37,0,145,0,0,0,96,0,229,0,201,0,0,0,0,0,54,0,79,0,56,0,0,0,88,0,237,0,91,0,35,0,219,0,0,0,210,0,1,0,234,0,148,0,37,0,0,0,106,0,174,0,49,0,217,0,155,0,192,0,19,0,60,0,47,0,39,0,217,0,0,0,180,0,76,0,124,0,0,0,195,0,34,0,197,0,165,0,138,0,167,0,28,0,218,0,189,0,229,0,208,0,4,0,50,0,14,0,199,0,0,0,197,0,68,0,103,0,207,0,194,0,0,0,129,0,26,0,6,0,19,0,184,0,47,0,48,0,98,0,115,0,0,0,0,0,0,0,31,0,231,0,160,0,0,0,239,0,106,0,67,0,39,0,0,0,151,0,107,0,81,0,50,0,0,0,6,0,97,0,158,0,0,0,122,0,17,0,194,0,0,0,254,0,218,0,0,0,33,0,0,0,192,0,246,0,0,0,184,0,126,0,36,0,228,0,134,0,250,0,55,0,0,0,165,0,234,0,194,0,202,0,98,0,141,0,47,0,211,0,0,0,60,0,34,0,0,0,0,0,157,0,226,0,244,0,0,0,229,0,148,0,133,0,124,0,186,0,31,0,192,0,0,0,235,0,24,0,219,0,0,0,77,0,191,0,79,0,113,0,15,0,239,0,3,0,58,0,229,0,220,0,204,0,59,0,254,0,71,0,7,0,0,0,231,0,75,0,139,0,76,0,0,0,152,0,0,0,117,0,0,0,221,0,56,0,0,0,0,0,83,0,234,0,219,0,50,0,0,0,207,0,77,0,0,0,208,0,159,0,11,0,0,0,93,0,48,0,144,0,147,0,61,0,150,0,29,0,0,0,60,0,246,0,177,0,220,0,189,0,103,0,0,0,179,0,250,0,100,0,232,0,88,0,90,0,7,0,0,0,74,0,243,0,133,0,250,0,175,0,0,0,183,0,182,0,41,0,31,0,169,0,53,0,68,0,239,0,0,0,215,0,108,0,220,0,253,0,81,0,153,0,253,0,71,0,120,0,235,0,4,0,232,0,174,0,0,0,242,0,91,0,86,0,81,0,137,0,163,0,207,0,147,0,0,0,151,0,165,0,232,0,63,0,51,0,146,0,0,0,0,0,150,0,69,0,248,0,166,0,0,0,36,0,26,0,2,0,85,0,70,0,0,0,164,0,178,0,99,0,198,0,55,0,194,0,79,0,58,0,184,0,121,0,49,0,21,0,95,0,69,0,81,0,141,0,218,0,240,0,22,0,29,0,248,0,25,0,232,0,212,0,167,0,168,0,96,0,43,0,0,0,0,0,0,0,62,0,118,0,241,0,44,0,166,0);
signal scenario_full  : scenario_type := (233,31,233,30,233,29,176,31,111,31,159,31,119,31,185,31,150,31,14,31,240,31,205,31,75,31,75,30,75,31,154,31,158,31,15,31,15,30,32,31,212,31,53,31,53,30,132,31,132,30,132,31,126,31,152,31,88,31,88,30,88,29,166,31,5,31,144,31,69,31,69,30,194,31,235,31,208,31,36,31,54,31,18,31,9,31,52,31,60,31,196,31,252,31,111,31,9,31,158,31,48,31,169,31,31,31,143,31,165,31,165,30,199,31,185,31,238,31,101,31,195,31,195,30,213,31,203,31,203,30,28,31,80,31,161,31,161,30,10,31,22,31,190,31,187,31,12,31,100,31,100,30,75,31,75,30,75,29,82,31,59,31,14,31,14,30,102,31,90,31,105,31,105,30,156,31,245,31,245,30,245,29,120,31,120,30,96,31,61,31,193,31,119,31,90,31,90,30,127,31,42,31,110,31,110,30,98,31,98,30,32,31,32,30,157,31,157,30,157,29,157,28,185,31,11,31,164,31,255,31,206,31,63,31,214,31,231,31,231,30,231,29,67,31,67,30,161,31,42,31,125,31,131,31,221,31,117,31,225,31,23,31,23,30,211,31,203,31,203,30,89,31,254,31,254,30,254,29,125,31,104,31,72,31,241,31,67,31,142,31,13,31,13,30,13,29,234,31,201,31,192,31,194,31,194,30,194,29,243,31,58,31,135,31,4,31,248,31,248,30,248,29,43,31,43,30,94,31,170,31,170,30,108,31,108,30,108,29,161,31,86,31,86,30,137,31,137,30,137,29,85,31,246,31,246,30,139,31,206,31,186,31,117,31,199,31,199,30,102,31,175,31,13,31,123,31,124,31,231,31,91,31,67,31,167,31,122,31,122,30,240,31,240,30,240,29,33,31,12,31,86,31,110,31,178,31,38,31,161,31,161,30,40,31,19,31,19,30,213,31,213,30,213,29,44,31,133,31,114,31,62,31,62,30,73,31,86,31,39,31,84,31,25,31,214,31,142,31,142,30,144,31,208,31,37,31,144,31,144,30,138,31,138,30,131,31,97,31,246,31,128,31,124,31,79,31,209,31,121,31,39,31,234,31,121,31,121,30,158,31,109,31,222,31,26,31,26,30,110,31,36,31,36,30,154,31,195,31,55,31,61,31,32,31,164,31,120,31,69,31,61,31,19,31,121,31,220,31,220,30,232,31,247,31,53,31,53,30,53,29,7,31,226,31,72,31,159,31,159,30,159,29,76,31,236,31,7,31,186,31,7,31,174,31,126,31,126,30,206,31,129,31,139,31,37,31,145,31,145,30,96,31,229,31,201,31,201,30,201,29,54,31,79,31,56,31,56,30,88,31,237,31,91,31,35,31,219,31,219,30,210,31,1,31,234,31,148,31,37,31,37,30,106,31,174,31,49,31,217,31,155,31,192,31,19,31,60,31,47,31,39,31,217,31,217,30,180,31,76,31,124,31,124,30,195,31,34,31,197,31,165,31,138,31,167,31,28,31,218,31,189,31,229,31,208,31,4,31,50,31,14,31,199,31,199,30,197,31,68,31,103,31,207,31,194,31,194,30,129,31,26,31,6,31,19,31,184,31,47,31,48,31,98,31,115,31,115,30,115,29,115,28,31,31,231,31,160,31,160,30,239,31,106,31,67,31,39,31,39,30,151,31,107,31,81,31,50,31,50,30,6,31,97,31,158,31,158,30,122,31,17,31,194,31,194,30,254,31,218,31,218,30,33,31,33,30,192,31,246,31,246,30,184,31,126,31,36,31,228,31,134,31,250,31,55,31,55,30,165,31,234,31,194,31,202,31,98,31,141,31,47,31,211,31,211,30,60,31,34,31,34,30,34,29,157,31,226,31,244,31,244,30,229,31,148,31,133,31,124,31,186,31,31,31,192,31,192,30,235,31,24,31,219,31,219,30,77,31,191,31,79,31,113,31,15,31,239,31,3,31,58,31,229,31,220,31,204,31,59,31,254,31,71,31,7,31,7,30,231,31,75,31,139,31,76,31,76,30,152,31,152,30,117,31,117,30,221,31,56,31,56,30,56,29,83,31,234,31,219,31,50,31,50,30,207,31,77,31,77,30,208,31,159,31,11,31,11,30,93,31,48,31,144,31,147,31,61,31,150,31,29,31,29,30,60,31,246,31,177,31,220,31,189,31,103,31,103,30,179,31,250,31,100,31,232,31,88,31,90,31,7,31,7,30,74,31,243,31,133,31,250,31,175,31,175,30,183,31,182,31,41,31,31,31,169,31,53,31,68,31,239,31,239,30,215,31,108,31,220,31,253,31,81,31,153,31,253,31,71,31,120,31,235,31,4,31,232,31,174,31,174,30,242,31,91,31,86,31,81,31,137,31,163,31,207,31,147,31,147,30,151,31,165,31,232,31,63,31,51,31,146,31,146,30,146,29,150,31,69,31,248,31,166,31,166,30,36,31,26,31,2,31,85,31,70,31,70,30,164,31,178,31,99,31,198,31,55,31,194,31,79,31,58,31,184,31,121,31,49,31,21,31,95,31,69,31,81,31,141,31,218,31,240,31,22,31,29,31,248,31,25,31,232,31,212,31,167,31,168,31,96,31,43,31,43,30,43,29,43,28,62,31,118,31,241,31,44,31,166,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
