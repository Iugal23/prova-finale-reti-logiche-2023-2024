-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 626;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (217,0,220,0,19,0,216,0,96,0,159,0,156,0,174,0,77,0,138,0,94,0,98,0,222,0,218,0,37,0,0,0,248,0,16,0,0,0,176,0,252,0,107,0,145,0,94,0,118,0,1,0,157,0,189,0,0,0,170,0,184,0,25,0,211,0,62,0,242,0,0,0,212,0,111,0,0,0,124,0,0,0,0,0,216,0,0,0,176,0,99,0,74,0,18,0,150,0,110,0,0,0,0,0,123,0,183,0,0,0,166,0,116,0,0,0,107,0,60,0,0,0,0,0,173,0,217,0,0,0,2,0,244,0,0,0,20,0,160,0,45,0,224,0,196,0,203,0,61,0,14,0,201,0,194,0,141,0,171,0,0,0,47,0,0,0,62,0,99,0,1,0,0,0,0,0,0,0,0,0,54,0,15,0,68,0,124,0,68,0,233,0,73,0,144,0,242,0,247,0,149,0,228,0,6,0,232,0,30,0,192,0,0,0,82,0,116,0,194,0,0,0,0,0,71,0,15,0,31,0,27,0,84,0,52,0,55,0,245,0,177,0,0,0,62,0,7,0,88,0,24,0,6,0,115,0,45,0,0,0,122,0,241,0,9,0,43,0,1,0,140,0,32,0,55,0,56,0,158,0,237,0,125,0,151,0,37,0,120,0,47,0,29,0,0,0,221,0,71,0,0,0,0,0,147,0,94,0,113,0,9,0,252,0,106,0,40,0,154,0,0,0,136,0,6,0,228,0,27,0,10,0,239,0,66,0,161,0,113,0,0,0,83,0,215,0,243,0,21,0,220,0,102,0,180,0,19,0,12,0,0,0,84,0,133,0,0,0,169,0,44,0,134,0,153,0,152,0,192,0,241,0,214,0,109,0,192,0,98,0,78,0,238,0,182,0,65,0,238,0,4,0,20,0,0,0,150,0,86,0,74,0,0,0,156,0,76,0,10,0,34,0,8,0,140,0,253,0,0,0,0,0,0,0,214,0,0,0,142,0,137,0,178,0,20,0,31,0,75,0,149,0,2,0,197,0,118,0,157,0,234,0,0,0,110,0,240,0,41,0,234,0,149,0,0,0,49,0,137,0,0,0,0,0,119,0,210,0,243,0,166,0,0,0,182,0,18,0,195,0,0,0,0,0,131,0,29,0,62,0,137,0,217,0,250,0,0,0,0,0,0,0,195,0,28,0,62,0,20,0,0,0,127,0,127,0,243,0,45,0,233,0,0,0,0,0,252,0,70,0,90,0,216,0,142,0,71,0,90,0,154,0,40,0,219,0,0,0,118,0,216,0,210,0,151,0,30,0,85,0,232,0,131,0,0,0,73,0,160,0,161,0,0,0,227,0,196,0,98,0,153,0,188,0,162,0,0,0,137,0,124,0,213,0,55,0,18,0,0,0,56,0,89,0,248,0,65,0,113,0,99,0,0,0,0,0,0,0,0,0,227,0,36,0,0,0,44,0,0,0,221,0,187,0,0,0,0,0,142,0,38,0,18,0,65,0,31,0,27,0,40,0,135,0,52,0,0,0,0,0,239,0,249,0,202,0,82,0,0,0,26,0,139,0,110,0,207,0,6,0,0,0,162,0,108,0,0,0,80,0,0,0,111,0,0,0,0,0,235,0,56,0,210,0,228,0,113,0,79,0,17,0,192,0,141,0,142,0,34,0,0,0,32,0,0,0,82,0,233,0,106,0,82,0,175,0,24,0,189,0,0,0,97,0,177,0,200,0,0,0,0,0,0,0,234,0,255,0,17,0,97,0,187,0,222,0,71,0,135,0,103,0,0,0,72,0,168,0,246,0,64,0,219,0,240,0,0,0,65,0,223,0,200,0,6,0,17,0,19,0,7,0,97,0,0,0,4,0,11,0,135,0,121,0,176,0,75,0,0,0,3,0,101,0,163,0,132,0,8,0,0,0,0,0,0,0,9,0,177,0,247,0,0,0,55,0,0,0,91,0,83,0,0,0,131,0,201,0,0,0,242,0,205,0,47,0,136,0,0,0,214,0,0,0,143,0,38,0,0,0,0,0,0,0,0,0,29,0,0,0,131,0,188,0,0,0,158,0,0,0,0,0,71,0,77,0,228,0,112,0,248,0,105,0,9,0,78,0,138,0,0,0,0,0,0,0,210,0,157,0,87,0,107,0,0,0,227,0,100,0,221,0,2,0,200,0,75,0,243,0,0,0,0,0,150,0,0,0,195,0,39,0,143,0,87,0,250,0,0,0,19,0,202,0,30,0,241,0,13,0,0,0,200,0,78,0,59,0,174,0,228,0,0,0,0,0,132,0,0,0,145,0,35,0,113,0,0,0,63,0,148,0,103,0,118,0,0,0,162,0,0,0,0,0,180,0,180,0,158,0,228,0,231,0,203,0,0,0,82,0,27,0,150,0,0,0,223,0,63,0,131,0,88,0,54,0,8,0,144,0,0,0,0,0,44,0,47,0,66,0,24,0,5,0,0,0,219,0,128,0,202,0,71,0,33,0,83,0,25,0,136,0,91,0,16,0,0,0,53,0,86,0,12,0,73,0,154,0,119,0,0,0,158,0,97,0,31,0,163,0,47,0,115,0,46,0,0,0,30,0,0,0,0,0,116,0,244,0,116,0,36,0,0,0,192,0,101,0,155,0,4,0,106,0,0,0,105,0,74,0,21,0,0,0,93,0,84,0,234,0,79,0,87,0,0,0,101,0,221,0,0,0,21,0,235,0,85,0,0,0,0,0,157,0,0,0,0,0,214,0,20,0,64,0,82,0,0,0,82,0,176,0,93,0,169,0,0,0,89,0,119,0,0,0,90,0,166,0,246,0,0,0);
signal scenario_full  : scenario_type := (217,31,220,31,19,31,216,31,96,31,159,31,156,31,174,31,77,31,138,31,94,31,98,31,222,31,218,31,37,31,37,30,248,31,16,31,16,30,176,31,252,31,107,31,145,31,94,31,118,31,1,31,157,31,189,31,189,30,170,31,184,31,25,31,211,31,62,31,242,31,242,30,212,31,111,31,111,30,124,31,124,30,124,29,216,31,216,30,176,31,99,31,74,31,18,31,150,31,110,31,110,30,110,29,123,31,183,31,183,30,166,31,116,31,116,30,107,31,60,31,60,30,60,29,173,31,217,31,217,30,2,31,244,31,244,30,20,31,160,31,45,31,224,31,196,31,203,31,61,31,14,31,201,31,194,31,141,31,171,31,171,30,47,31,47,30,62,31,99,31,1,31,1,30,1,29,1,28,1,27,54,31,15,31,68,31,124,31,68,31,233,31,73,31,144,31,242,31,247,31,149,31,228,31,6,31,232,31,30,31,192,31,192,30,82,31,116,31,194,31,194,30,194,29,71,31,15,31,31,31,27,31,84,31,52,31,55,31,245,31,177,31,177,30,62,31,7,31,88,31,24,31,6,31,115,31,45,31,45,30,122,31,241,31,9,31,43,31,1,31,140,31,32,31,55,31,56,31,158,31,237,31,125,31,151,31,37,31,120,31,47,31,29,31,29,30,221,31,71,31,71,30,71,29,147,31,94,31,113,31,9,31,252,31,106,31,40,31,154,31,154,30,136,31,6,31,228,31,27,31,10,31,239,31,66,31,161,31,113,31,113,30,83,31,215,31,243,31,21,31,220,31,102,31,180,31,19,31,12,31,12,30,84,31,133,31,133,30,169,31,44,31,134,31,153,31,152,31,192,31,241,31,214,31,109,31,192,31,98,31,78,31,238,31,182,31,65,31,238,31,4,31,20,31,20,30,150,31,86,31,74,31,74,30,156,31,76,31,10,31,34,31,8,31,140,31,253,31,253,30,253,29,253,28,214,31,214,30,142,31,137,31,178,31,20,31,31,31,75,31,149,31,2,31,197,31,118,31,157,31,234,31,234,30,110,31,240,31,41,31,234,31,149,31,149,30,49,31,137,31,137,30,137,29,119,31,210,31,243,31,166,31,166,30,182,31,18,31,195,31,195,30,195,29,131,31,29,31,62,31,137,31,217,31,250,31,250,30,250,29,250,28,195,31,28,31,62,31,20,31,20,30,127,31,127,31,243,31,45,31,233,31,233,30,233,29,252,31,70,31,90,31,216,31,142,31,71,31,90,31,154,31,40,31,219,31,219,30,118,31,216,31,210,31,151,31,30,31,85,31,232,31,131,31,131,30,73,31,160,31,161,31,161,30,227,31,196,31,98,31,153,31,188,31,162,31,162,30,137,31,124,31,213,31,55,31,18,31,18,30,56,31,89,31,248,31,65,31,113,31,99,31,99,30,99,29,99,28,99,27,227,31,36,31,36,30,44,31,44,30,221,31,187,31,187,30,187,29,142,31,38,31,18,31,65,31,31,31,27,31,40,31,135,31,52,31,52,30,52,29,239,31,249,31,202,31,82,31,82,30,26,31,139,31,110,31,207,31,6,31,6,30,162,31,108,31,108,30,80,31,80,30,111,31,111,30,111,29,235,31,56,31,210,31,228,31,113,31,79,31,17,31,192,31,141,31,142,31,34,31,34,30,32,31,32,30,82,31,233,31,106,31,82,31,175,31,24,31,189,31,189,30,97,31,177,31,200,31,200,30,200,29,200,28,234,31,255,31,17,31,97,31,187,31,222,31,71,31,135,31,103,31,103,30,72,31,168,31,246,31,64,31,219,31,240,31,240,30,65,31,223,31,200,31,6,31,17,31,19,31,7,31,97,31,97,30,4,31,11,31,135,31,121,31,176,31,75,31,75,30,3,31,101,31,163,31,132,31,8,31,8,30,8,29,8,28,9,31,177,31,247,31,247,30,55,31,55,30,91,31,83,31,83,30,131,31,201,31,201,30,242,31,205,31,47,31,136,31,136,30,214,31,214,30,143,31,38,31,38,30,38,29,38,28,38,27,29,31,29,30,131,31,188,31,188,30,158,31,158,30,158,29,71,31,77,31,228,31,112,31,248,31,105,31,9,31,78,31,138,31,138,30,138,29,138,28,210,31,157,31,87,31,107,31,107,30,227,31,100,31,221,31,2,31,200,31,75,31,243,31,243,30,243,29,150,31,150,30,195,31,39,31,143,31,87,31,250,31,250,30,19,31,202,31,30,31,241,31,13,31,13,30,200,31,78,31,59,31,174,31,228,31,228,30,228,29,132,31,132,30,145,31,35,31,113,31,113,30,63,31,148,31,103,31,118,31,118,30,162,31,162,30,162,29,180,31,180,31,158,31,228,31,231,31,203,31,203,30,82,31,27,31,150,31,150,30,223,31,63,31,131,31,88,31,54,31,8,31,144,31,144,30,144,29,44,31,47,31,66,31,24,31,5,31,5,30,219,31,128,31,202,31,71,31,33,31,83,31,25,31,136,31,91,31,16,31,16,30,53,31,86,31,12,31,73,31,154,31,119,31,119,30,158,31,97,31,31,31,163,31,47,31,115,31,46,31,46,30,30,31,30,30,30,29,116,31,244,31,116,31,36,31,36,30,192,31,101,31,155,31,4,31,106,31,106,30,105,31,74,31,21,31,21,30,93,31,84,31,234,31,79,31,87,31,87,30,101,31,221,31,221,30,21,31,235,31,85,31,85,30,85,29,157,31,157,30,157,29,214,31,20,31,64,31,82,31,82,30,82,31,176,31,93,31,169,31,169,30,89,31,119,31,119,30,90,31,166,31,246,31,246,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
