-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 169;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (156,0,0,0,13,0,86,0,131,0,185,0,0,0,0,0,181,0,216,0,191,0,106,0,0,0,71,0,49,0,0,0,19,0,0,0,162,0,0,0,100,0,43,0,0,0,110,0,199,0,79,0,151,0,0,0,18,0,245,0,0,0,101,0,0,0,177,0,163,0,127,0,0,0,219,0,85,0,82,0,11,0,197,0,44,0,140,0,146,0,85,0,253,0,223,0,173,0,12,0,46,0,209,0,178,0,126,0,25,0,214,0,85,0,230,0,175,0,113,0,120,0,0,0,57,0,247,0,90,0,174,0,57,0,112,0,164,0,130,0,224,0,212,0,126,0,86,0,0,0,133,0,34,0,98,0,93,0,0,0,91,0,177,0,112,0,8,0,24,0,238,0,173,0,64,0,142,0,87,0,194,0,128,0,154,0,70,0,37,0,39,0,208,0,25,0,0,0,41,0,202,0,231,0,253,0,62,0,58,0,5,0,0,0,133,0,208,0,91,0,90,0,49,0,17,0,161,0,0,0,206,0,152,0,10,0,144,0,87,0,229,0,49,0,84,0,185,0,170,0,43,0,49,0,132,0,162,0,23,0,0,0,77,0,120,0,86,0,0,0,98,0,10,0,4,0,165,0,19,0,168,0,137,0,77,0,148,0,234,0,125,0,229,0,179,0,142,0,94,0,223,0,0,0,249,0,155,0,236,0,91,0,110,0,29,0,0,0,122,0,11,0,35,0,223,0,91,0,125,0,107,0,87,0,248,0,130,0);
signal scenario_full  : scenario_type := (156,31,156,30,13,31,86,31,131,31,185,31,185,30,185,29,181,31,216,31,191,31,106,31,106,30,71,31,49,31,49,30,19,31,19,30,162,31,162,30,100,31,43,31,43,30,110,31,199,31,79,31,151,31,151,30,18,31,245,31,245,30,101,31,101,30,177,31,163,31,127,31,127,30,219,31,85,31,82,31,11,31,197,31,44,31,140,31,146,31,85,31,253,31,223,31,173,31,12,31,46,31,209,31,178,31,126,31,25,31,214,31,85,31,230,31,175,31,113,31,120,31,120,30,57,31,247,31,90,31,174,31,57,31,112,31,164,31,130,31,224,31,212,31,126,31,86,31,86,30,133,31,34,31,98,31,93,31,93,30,91,31,177,31,112,31,8,31,24,31,238,31,173,31,64,31,142,31,87,31,194,31,128,31,154,31,70,31,37,31,39,31,208,31,25,31,25,30,41,31,202,31,231,31,253,31,62,31,58,31,5,31,5,30,133,31,208,31,91,31,90,31,49,31,17,31,161,31,161,30,206,31,152,31,10,31,144,31,87,31,229,31,49,31,84,31,185,31,170,31,43,31,49,31,132,31,162,31,23,31,23,30,77,31,120,31,86,31,86,30,98,31,10,31,4,31,165,31,19,31,168,31,137,31,77,31,148,31,234,31,125,31,229,31,179,31,142,31,94,31,223,31,223,30,249,31,155,31,236,31,91,31,110,31,29,31,29,30,122,31,11,31,35,31,223,31,91,31,125,31,107,31,87,31,248,31,130,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
