-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 335;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (175,0,185,0,0,0,18,0,0,0,3,0,216,0,70,0,223,0,200,0,1,0,111,0,205,0,0,0,85,0,173,0,58,0,196,0,0,0,159,0,200,0,102,0,198,0,126,0,0,0,148,0,0,0,103,0,198,0,42,0,131,0,147,0,244,0,161,0,179,0,0,0,205,0,186,0,0,0,190,0,233,0,243,0,0,0,69,0,249,0,252,0,151,0,85,0,13,0,179,0,218,0,164,0,34,0,190,0,0,0,0,0,0,0,228,0,0,0,51,0,241,0,252,0,0,0,151,0,224,0,8,0,78,0,105,0,0,0,21,0,71,0,0,0,33,0,40,0,188,0,246,0,198,0,0,0,127,0,216,0,41,0,0,0,69,0,143,0,0,0,68,0,229,0,180,0,0,0,161,0,9,0,93,0,140,0,253,0,124,0,12,0,39,0,2,0,15,0,40,0,75,0,0,0,101,0,178,0,0,0,128,0,11,0,32,0,73,0,91,0,0,0,255,0,213,0,52,0,178,0,0,0,73,0,110,0,0,0,11,0,87,0,198,0,29,0,247,0,43,0,233,0,200,0,231,0,172,0,30,0,131,0,137,0,0,0,11,0,49,0,143,0,0,0,71,0,10,0,207,0,98,0,217,0,201,0,0,0,9,0,166,0,204,0,23,0,27,0,51,0,194,0,134,0,119,0,192,0,110,0,46,0,50,0,21,0,225,0,193,0,192,0,207,0,28,0,150,0,96,0,155,0,164,0,7,0,221,0,80,0,150,0,150,0,4,0,127,0,227,0,0,0,0,0,180,0,84,0,96,0,80,0,37,0,74,0,47,0,25,0,114,0,207,0,179,0,97,0,157,0,81,0,0,0,241,0,219,0,68,0,38,0,108,0,186,0,140,0,0,0,82,0,0,0,86,0,0,0,191,0,39,0,97,0,0,0,221,0,91,0,69,0,8,0,52,0,0,0,73,0,0,0,213,0,138,0,119,0,208,0,0,0,59,0,110,0,169,0,65,0,13,0,247,0,0,0,0,0,240,0,169,0,79,0,83,0,151,0,178,0,93,0,217,0,1,0,0,0,0,0,182,0,14,0,179,0,0,0,153,0,0,0,77,0,174,0,103,0,0,0,0,0,2,0,0,0,245,0,0,0,0,0,0,0,27,0,12,0,185,0,0,0,217,0,221,0,145,0,153,0,68,0,0,0,172,0,0,0,0,0,0,0,119,0,175,0,106,0,119,0,178,0,169,0,199,0,0,0,89,0,156,0,111,0,51,0,237,0,69,0,118,0,239,0,81,0,32,0,37,0,0,0,24,0,159,0,0,0,83,0,76,0,252,0,127,0,0,0,120,0,194,0,229,0,178,0,235,0,0,0,142,0,185,0,245,0,185,0,2,0,0,0,124,0,248,0,224,0,204,0,204,0,74,0,88,0,186,0,149,0,252,0,222,0,0,0,15,0,208,0,171,0,113,0,0,0,0,0,144,0,86,0,120,0,160,0,0,0,247,0);
signal scenario_full  : scenario_type := (175,31,185,31,185,30,18,31,18,30,3,31,216,31,70,31,223,31,200,31,1,31,111,31,205,31,205,30,85,31,173,31,58,31,196,31,196,30,159,31,200,31,102,31,198,31,126,31,126,30,148,31,148,30,103,31,198,31,42,31,131,31,147,31,244,31,161,31,179,31,179,30,205,31,186,31,186,30,190,31,233,31,243,31,243,30,69,31,249,31,252,31,151,31,85,31,13,31,179,31,218,31,164,31,34,31,190,31,190,30,190,29,190,28,228,31,228,30,51,31,241,31,252,31,252,30,151,31,224,31,8,31,78,31,105,31,105,30,21,31,71,31,71,30,33,31,40,31,188,31,246,31,198,31,198,30,127,31,216,31,41,31,41,30,69,31,143,31,143,30,68,31,229,31,180,31,180,30,161,31,9,31,93,31,140,31,253,31,124,31,12,31,39,31,2,31,15,31,40,31,75,31,75,30,101,31,178,31,178,30,128,31,11,31,32,31,73,31,91,31,91,30,255,31,213,31,52,31,178,31,178,30,73,31,110,31,110,30,11,31,87,31,198,31,29,31,247,31,43,31,233,31,200,31,231,31,172,31,30,31,131,31,137,31,137,30,11,31,49,31,143,31,143,30,71,31,10,31,207,31,98,31,217,31,201,31,201,30,9,31,166,31,204,31,23,31,27,31,51,31,194,31,134,31,119,31,192,31,110,31,46,31,50,31,21,31,225,31,193,31,192,31,207,31,28,31,150,31,96,31,155,31,164,31,7,31,221,31,80,31,150,31,150,31,4,31,127,31,227,31,227,30,227,29,180,31,84,31,96,31,80,31,37,31,74,31,47,31,25,31,114,31,207,31,179,31,97,31,157,31,81,31,81,30,241,31,219,31,68,31,38,31,108,31,186,31,140,31,140,30,82,31,82,30,86,31,86,30,191,31,39,31,97,31,97,30,221,31,91,31,69,31,8,31,52,31,52,30,73,31,73,30,213,31,138,31,119,31,208,31,208,30,59,31,110,31,169,31,65,31,13,31,247,31,247,30,247,29,240,31,169,31,79,31,83,31,151,31,178,31,93,31,217,31,1,31,1,30,1,29,182,31,14,31,179,31,179,30,153,31,153,30,77,31,174,31,103,31,103,30,103,29,2,31,2,30,245,31,245,30,245,29,245,28,27,31,12,31,185,31,185,30,217,31,221,31,145,31,153,31,68,31,68,30,172,31,172,30,172,29,172,28,119,31,175,31,106,31,119,31,178,31,169,31,199,31,199,30,89,31,156,31,111,31,51,31,237,31,69,31,118,31,239,31,81,31,32,31,37,31,37,30,24,31,159,31,159,30,83,31,76,31,252,31,127,31,127,30,120,31,194,31,229,31,178,31,235,31,235,30,142,31,185,31,245,31,185,31,2,31,2,30,124,31,248,31,224,31,204,31,204,31,74,31,88,31,186,31,149,31,252,31,222,31,222,30,15,31,208,31,171,31,113,31,113,30,113,29,144,31,86,31,120,31,160,31,160,30,247,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
