-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_320 is
end project_tb_320;

architecture project_tb_arch_320 of project_tb_320 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 729;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,192,0,184,0,9,0,33,0,102,0,151,0,166,0,59,0,72,0,87,0,175,0,0,0,51,0,246,0,0,0,234,0,30,0,0,0,0,0,117,0,0,0,209,0,0,0,158,0,223,0,0,0,224,0,166,0,119,0,125,0,10,0,45,0,0,0,0,0,230,0,251,0,232,0,215,0,45,0,153,0,162,0,0,0,0,0,126,0,21,0,0,0,0,0,79,0,0,0,0,0,16,0,183,0,177,0,84,0,0,0,192,0,28,0,107,0,174,0,48,0,0,0,149,0,200,0,31,0,21,0,222,0,136,0,33,0,0,0,0,0,69,0,0,0,59,0,204,0,0,0,147,0,0,0,0,0,107,0,0,0,108,0,48,0,236,0,206,0,5,0,87,0,251,0,148,0,34,0,121,0,157,0,0,0,64,0,51,0,139,0,16,0,0,0,182,0,197,0,211,0,202,0,29,0,203,0,119,0,246,0,120,0,231,0,0,0,92,0,86,0,52,0,176,0,135,0,51,0,200,0,230,0,54,0,35,0,23,0,232,0,41,0,0,0,142,0,136,0,109,0,18,0,160,0,189,0,0,0,98,0,0,0,91,0,0,0,238,0,159,0,219,0,104,0,78,0,208,0,178,0,35,0,241,0,0,0,194,0,0,0,80,0,134,0,0,0,244,0,3,0,189,0,241,0,245,0,34,0,0,0,190,0,11,0,30,0,110,0,195,0,112,0,103,0,17,0,74,0,235,0,0,0,0,0,170,0,68,0,178,0,133,0,86,0,0,0,0,0,37,0,9,0,171,0,82,0,137,0,183,0,214,0,39,0,12,0,17,0,177,0,92,0,0,0,118,0,0,0,171,0,44,0,0,0,0,0,114,0,148,0,58,0,77,0,227,0,9,0,232,0,67,0,38,0,0,0,230,0,0,0,185,0,108,0,120,0,203,0,232,0,0,0,0,0,245,0,0,0,87,0,127,0,0,0,23,0,0,0,176,0,170,0,204,0,57,0,248,0,67,0,142,0,0,0,242,0,0,0,33,0,174,0,64,0,133,0,47,0,169,0,64,0,126,0,0,0,0,0,108,0,233,0,162,0,45,0,14,0,52,0,0,0,153,0,93,0,74,0,169,0,0,0,161,0,22,0,51,0,255,0,152,0,79,0,0,0,197,0,181,0,71,0,28,0,122,0,209,0,0,0,94,0,223,0,224,0,116,0,143,0,196,0,0,0,109,0,0,0,156,0,237,0,0,0,133,0,0,0,45,0,158,0,0,0,0,0,193,0,93,0,31,0,104,0,11,0,230,0,229,0,0,0,43,0,154,0,201,0,0,0,162,0,93,0,37,0,237,0,0,0,241,0,245,0,6,0,228,0,144,0,48,0,198,0,0,0,182,0,64,0,0,0,6,0,6,0,207,0,213,0,160,0,88,0,198,0,83,0,76,0,104,0,111,0,44,0,241,0,93,0,244,0,7,0,173,0,51,0,86,0,137,0,0,0,0,0,169,0,165,0,16,0,0,0,13,0,178,0,0,0,168,0,145,0,0,0,117,0,241,0,223,0,254,0,0,0,186,0,142,0,238,0,0,0,0,0,228,0,44,0,9,0,243,0,216,0,33,0,251,0,187,0,187,0,29,0,38,0,115,0,216,0,118,0,246,0,34,0,93,0,186,0,214,0,216,0,21,0,59,0,64,0,64,0,31,0,252,0,123,0,207,0,164,0,0,0,0,0,162,0,111,0,27,0,12,0,17,0,59,0,135,0,15,0,121,0,156,0,147,0,164,0,175,0,0,0,0,0,226,0,33,0,0,0,138,0,6,0,174,0,102,0,82,0,0,0,43,0,162,0,0,0,123,0,116,0,151,0,194,0,0,0,214,0,186,0,16,0,100,0,42,0,189,0,19,0,0,0,138,0,215,0,254,0,238,0,155,0,230,0,109,0,5,0,112,0,176,0,169,0,233,0,0,0,1,0,232,0,14,0,128,0,0,0,200,0,219,0,0,0,58,0,221,0,198,0,0,0,0,0,137,0,176,0,0,0,199,0,176,0,207,0,155,0,219,0,209,0,19,0,0,0,0,0,84,0,16,0,95,0,240,0,200,0,0,0,55,0,175,0,180,0,211,0,207,0,116,0,1,0,193,0,66,0,7,0,78,0,0,0,0,0,38,0,165,0,183,0,0,0,140,0,179,0,108,0,156,0,46,0,100,0,237,0,146,0,0,0,45,0,7,0,124,0,0,0,97,0,0,0,176,0,136,0,247,0,139,0,245,0,37,0,167,0,22,0,76,0,0,0,235,0,22,0,17,0,122,0,29,0,148,0,113,0,31,0,66,0,204,0,0,0,177,0,81,0,156,0,100,0,116,0,178,0,147,0,5,0,200,0,73,0,42,0,107,0,138,0,0,0,172,0,51,0,0,0,68,0,241,0,196,0,236,0,119,0,207,0,0,0,177,0,150,0,0,0,213,0,191,0,185,0,166,0,15,0,134,0,126,0,136,0,237,0,59,0,52,0,13,0,196,0,0,0,108,0,0,0,2,0,19,0,235,0,60,0,0,0,185,0,0,0,80,0,160,0,144,0,182,0,180,0,140,0,10,0,226,0,53,0,173,0,0,0,209,0,167,0,43,0,240,0,0,0,255,0,186,0,0,0,143,0,33,0,61,0,0,0,3,0,207,0,134,0,176,0,120,0,22,0,139,0,251,0,105,0,142,0,99,0,140,0,230,0,72,0,0,0,161,0,133,0,231,0,0,0,8,0,149,0,91,0,177,0,73,0,0,0,83,0,238,0,0,0,220,0,80,0,67,0,33,0,83,0,188,0,52,0,0,0,58,0,184,0,0,0,133,0,224,0,36,0,90,0,234,0,0,0,108,0,0,0,132,0,156,0,158,0,0,0,0,0,169,0,0,0,138,0,0,0,0,0,50,0,106,0,15,0,185,0,171,0,0,0,0,0,0,0,240,0,177,0,0,0,112,0,0,0,0,0,113,0,139,0,16,0,47,0,0,0,47,0,0,0,112,0,149,0,183,0,143,0,97,0,46,0,123,0,233,0,66,0,0,0,29,0,203,0,243,0,246,0,225,0,155,0,197,0,0,0,41,0,71,0,58,0,0,0,210,0,26,0,105,0,91,0,45,0,97,0,0,0,29,0,94,0,178,0,226,0,0,0,212,0,221,0,35,0,227,0,222,0,195,0,187,0,97,0,253,0,224,0,0,0,0,0,248,0,184,0,0,0,41,0,218,0,85,0,14,0,199,0,96,0);
signal scenario_full  : scenario_type := (0,0,0,0,192,31,184,31,9,31,33,31,102,31,151,31,166,31,59,31,72,31,87,31,175,31,175,30,51,31,246,31,246,30,234,31,30,31,30,30,30,29,117,31,117,30,209,31,209,30,158,31,223,31,223,30,224,31,166,31,119,31,125,31,10,31,45,31,45,30,45,29,230,31,251,31,232,31,215,31,45,31,153,31,162,31,162,30,162,29,126,31,21,31,21,30,21,29,79,31,79,30,79,29,16,31,183,31,177,31,84,31,84,30,192,31,28,31,107,31,174,31,48,31,48,30,149,31,200,31,31,31,21,31,222,31,136,31,33,31,33,30,33,29,69,31,69,30,59,31,204,31,204,30,147,31,147,30,147,29,107,31,107,30,108,31,48,31,236,31,206,31,5,31,87,31,251,31,148,31,34,31,121,31,157,31,157,30,64,31,51,31,139,31,16,31,16,30,182,31,197,31,211,31,202,31,29,31,203,31,119,31,246,31,120,31,231,31,231,30,92,31,86,31,52,31,176,31,135,31,51,31,200,31,230,31,54,31,35,31,23,31,232,31,41,31,41,30,142,31,136,31,109,31,18,31,160,31,189,31,189,30,98,31,98,30,91,31,91,30,238,31,159,31,219,31,104,31,78,31,208,31,178,31,35,31,241,31,241,30,194,31,194,30,80,31,134,31,134,30,244,31,3,31,189,31,241,31,245,31,34,31,34,30,190,31,11,31,30,31,110,31,195,31,112,31,103,31,17,31,74,31,235,31,235,30,235,29,170,31,68,31,178,31,133,31,86,31,86,30,86,29,37,31,9,31,171,31,82,31,137,31,183,31,214,31,39,31,12,31,17,31,177,31,92,31,92,30,118,31,118,30,171,31,44,31,44,30,44,29,114,31,148,31,58,31,77,31,227,31,9,31,232,31,67,31,38,31,38,30,230,31,230,30,185,31,108,31,120,31,203,31,232,31,232,30,232,29,245,31,245,30,87,31,127,31,127,30,23,31,23,30,176,31,170,31,204,31,57,31,248,31,67,31,142,31,142,30,242,31,242,30,33,31,174,31,64,31,133,31,47,31,169,31,64,31,126,31,126,30,126,29,108,31,233,31,162,31,45,31,14,31,52,31,52,30,153,31,93,31,74,31,169,31,169,30,161,31,22,31,51,31,255,31,152,31,79,31,79,30,197,31,181,31,71,31,28,31,122,31,209,31,209,30,94,31,223,31,224,31,116,31,143,31,196,31,196,30,109,31,109,30,156,31,237,31,237,30,133,31,133,30,45,31,158,31,158,30,158,29,193,31,93,31,31,31,104,31,11,31,230,31,229,31,229,30,43,31,154,31,201,31,201,30,162,31,93,31,37,31,237,31,237,30,241,31,245,31,6,31,228,31,144,31,48,31,198,31,198,30,182,31,64,31,64,30,6,31,6,31,207,31,213,31,160,31,88,31,198,31,83,31,76,31,104,31,111,31,44,31,241,31,93,31,244,31,7,31,173,31,51,31,86,31,137,31,137,30,137,29,169,31,165,31,16,31,16,30,13,31,178,31,178,30,168,31,145,31,145,30,117,31,241,31,223,31,254,31,254,30,186,31,142,31,238,31,238,30,238,29,228,31,44,31,9,31,243,31,216,31,33,31,251,31,187,31,187,31,29,31,38,31,115,31,216,31,118,31,246,31,34,31,93,31,186,31,214,31,216,31,21,31,59,31,64,31,64,31,31,31,252,31,123,31,207,31,164,31,164,30,164,29,162,31,111,31,27,31,12,31,17,31,59,31,135,31,15,31,121,31,156,31,147,31,164,31,175,31,175,30,175,29,226,31,33,31,33,30,138,31,6,31,174,31,102,31,82,31,82,30,43,31,162,31,162,30,123,31,116,31,151,31,194,31,194,30,214,31,186,31,16,31,100,31,42,31,189,31,19,31,19,30,138,31,215,31,254,31,238,31,155,31,230,31,109,31,5,31,112,31,176,31,169,31,233,31,233,30,1,31,232,31,14,31,128,31,128,30,200,31,219,31,219,30,58,31,221,31,198,31,198,30,198,29,137,31,176,31,176,30,199,31,176,31,207,31,155,31,219,31,209,31,19,31,19,30,19,29,84,31,16,31,95,31,240,31,200,31,200,30,55,31,175,31,180,31,211,31,207,31,116,31,1,31,193,31,66,31,7,31,78,31,78,30,78,29,38,31,165,31,183,31,183,30,140,31,179,31,108,31,156,31,46,31,100,31,237,31,146,31,146,30,45,31,7,31,124,31,124,30,97,31,97,30,176,31,136,31,247,31,139,31,245,31,37,31,167,31,22,31,76,31,76,30,235,31,22,31,17,31,122,31,29,31,148,31,113,31,31,31,66,31,204,31,204,30,177,31,81,31,156,31,100,31,116,31,178,31,147,31,5,31,200,31,73,31,42,31,107,31,138,31,138,30,172,31,51,31,51,30,68,31,241,31,196,31,236,31,119,31,207,31,207,30,177,31,150,31,150,30,213,31,191,31,185,31,166,31,15,31,134,31,126,31,136,31,237,31,59,31,52,31,13,31,196,31,196,30,108,31,108,30,2,31,19,31,235,31,60,31,60,30,185,31,185,30,80,31,160,31,144,31,182,31,180,31,140,31,10,31,226,31,53,31,173,31,173,30,209,31,167,31,43,31,240,31,240,30,255,31,186,31,186,30,143,31,33,31,61,31,61,30,3,31,207,31,134,31,176,31,120,31,22,31,139,31,251,31,105,31,142,31,99,31,140,31,230,31,72,31,72,30,161,31,133,31,231,31,231,30,8,31,149,31,91,31,177,31,73,31,73,30,83,31,238,31,238,30,220,31,80,31,67,31,33,31,83,31,188,31,52,31,52,30,58,31,184,31,184,30,133,31,224,31,36,31,90,31,234,31,234,30,108,31,108,30,132,31,156,31,158,31,158,30,158,29,169,31,169,30,138,31,138,30,138,29,50,31,106,31,15,31,185,31,171,31,171,30,171,29,171,28,240,31,177,31,177,30,112,31,112,30,112,29,113,31,139,31,16,31,47,31,47,30,47,31,47,30,112,31,149,31,183,31,143,31,97,31,46,31,123,31,233,31,66,31,66,30,29,31,203,31,243,31,246,31,225,31,155,31,197,31,197,30,41,31,71,31,58,31,58,30,210,31,26,31,105,31,91,31,45,31,97,31,97,30,29,31,94,31,178,31,226,31,226,30,212,31,221,31,35,31,227,31,222,31,195,31,187,31,97,31,253,31,224,31,224,30,224,29,248,31,184,31,184,30,41,31,218,31,85,31,14,31,199,31,96,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
