-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_23 is
end project_tb_23;

architecture project_tb_arch_23 of project_tb_23 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 323;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (105,0,147,0,86,0,193,0,122,0,236,0,189,0,177,0,253,0,159,0,32,0,0,0,37,0,0,0,133,0,245,0,103,0,54,0,209,0,146,0,142,0,46,0,105,0,0,0,209,0,101,0,0,0,196,0,32,0,34,0,241,0,199,0,0,0,0,0,251,0,105,0,239,0,119,0,92,0,29,0,0,0,31,0,0,0,236,0,0,0,244,0,29,0,68,0,83,0,0,0,247,0,60,0,215,0,151,0,183,0,17,0,178,0,183,0,35,0,124,0,88,0,77,0,140,0,0,0,161,0,58,0,88,0,61,0,0,0,193,0,241,0,231,0,205,0,129,0,56,0,42,0,205,0,180,0,96,0,173,0,0,0,140,0,0,0,37,0,0,0,18,0,0,0,32,0,11,0,0,0,10,0,137,0,62,0,78,0,0,0,124,0,223,0,129,0,0,0,230,0,74,0,0,0,240,0,201,0,73,0,8,0,251,0,35,0,197,0,168,0,223,0,173,0,6,0,204,0,114,0,47,0,241,0,101,0,192,0,51,0,59,0,0,0,88,0,0,0,3,0,94,0,208,0,0,0,235,0,94,0,0,0,62,0,112,0,0,0,131,0,229,0,163,0,22,0,250,0,0,0,62,0,193,0,175,0,128,0,42,0,254,0,0,0,115,0,93,0,14,0,240,0,223,0,162,0,253,0,29,0,61,0,243,0,169,0,235,0,40,0,244,0,142,0,222,0,213,0,107,0,3,0,121,0,56,0,161,0,145,0,0,0,46,0,0,0,54,0,49,0,0,0,176,0,76,0,192,0,169,0,195,0,75,0,0,0,234,0,0,0,53,0,0,0,233,0,74,0,99,0,175,0,0,0,48,0,0,0,216,0,58,0,0,0,84,0,0,0,180,0,207,0,27,0,26,0,0,0,128,0,144,0,164,0,223,0,77,0,197,0,164,0,230,0,146,0,252,0,227,0,154,0,15,0,80,0,247,0,0,0,42,0,0,0,154,0,0,0,47,0,105,0,3,0,20,0,67,0,186,0,0,0,210,0,212,0,214,0,140,0,238,0,129,0,0,0,217,0,185,0,129,0,59,0,30,0,13,0,54,0,166,0,82,0,47,0,0,0,199,0,0,0,0,0,4,0,28,0,247,0,0,0,92,0,106,0,173,0,79,0,51,0,4,0,0,0,86,0,0,0,0,0,0,0,0,0,245,0,6,0,100,0,77,0,136,0,0,0,91,0,61,0,0,0,206,0,153,0,40,0,0,0,219,0,53,0,75,0,0,0,67,0,70,0,160,0,0,0,0,0,34,0,0,0,224,0,135,0,69,0,0,0,96,0,0,0,0,0,90,0,13,0,41,0,225,0,170,0,197,0,0,0,217,0,0,0,64,0,224,0,19,0,93,0,46,0,111,0,50,0,103,0,25,0,209,0,58,0,0,0,54,0,0,0,157,0);
signal scenario_full  : scenario_type := (105,31,147,31,86,31,193,31,122,31,236,31,189,31,177,31,253,31,159,31,32,31,32,30,37,31,37,30,133,31,245,31,103,31,54,31,209,31,146,31,142,31,46,31,105,31,105,30,209,31,101,31,101,30,196,31,32,31,34,31,241,31,199,31,199,30,199,29,251,31,105,31,239,31,119,31,92,31,29,31,29,30,31,31,31,30,236,31,236,30,244,31,29,31,68,31,83,31,83,30,247,31,60,31,215,31,151,31,183,31,17,31,178,31,183,31,35,31,124,31,88,31,77,31,140,31,140,30,161,31,58,31,88,31,61,31,61,30,193,31,241,31,231,31,205,31,129,31,56,31,42,31,205,31,180,31,96,31,173,31,173,30,140,31,140,30,37,31,37,30,18,31,18,30,32,31,11,31,11,30,10,31,137,31,62,31,78,31,78,30,124,31,223,31,129,31,129,30,230,31,74,31,74,30,240,31,201,31,73,31,8,31,251,31,35,31,197,31,168,31,223,31,173,31,6,31,204,31,114,31,47,31,241,31,101,31,192,31,51,31,59,31,59,30,88,31,88,30,3,31,94,31,208,31,208,30,235,31,94,31,94,30,62,31,112,31,112,30,131,31,229,31,163,31,22,31,250,31,250,30,62,31,193,31,175,31,128,31,42,31,254,31,254,30,115,31,93,31,14,31,240,31,223,31,162,31,253,31,29,31,61,31,243,31,169,31,235,31,40,31,244,31,142,31,222,31,213,31,107,31,3,31,121,31,56,31,161,31,145,31,145,30,46,31,46,30,54,31,49,31,49,30,176,31,76,31,192,31,169,31,195,31,75,31,75,30,234,31,234,30,53,31,53,30,233,31,74,31,99,31,175,31,175,30,48,31,48,30,216,31,58,31,58,30,84,31,84,30,180,31,207,31,27,31,26,31,26,30,128,31,144,31,164,31,223,31,77,31,197,31,164,31,230,31,146,31,252,31,227,31,154,31,15,31,80,31,247,31,247,30,42,31,42,30,154,31,154,30,47,31,105,31,3,31,20,31,67,31,186,31,186,30,210,31,212,31,214,31,140,31,238,31,129,31,129,30,217,31,185,31,129,31,59,31,30,31,13,31,54,31,166,31,82,31,47,31,47,30,199,31,199,30,199,29,4,31,28,31,247,31,247,30,92,31,106,31,173,31,79,31,51,31,4,31,4,30,86,31,86,30,86,29,86,28,86,27,245,31,6,31,100,31,77,31,136,31,136,30,91,31,61,31,61,30,206,31,153,31,40,31,40,30,219,31,53,31,75,31,75,30,67,31,70,31,160,31,160,30,160,29,34,31,34,30,224,31,135,31,69,31,69,30,96,31,96,30,96,29,90,31,13,31,41,31,225,31,170,31,197,31,197,30,217,31,217,30,64,31,224,31,19,31,93,31,46,31,111,31,50,31,103,31,25,31,209,31,58,31,58,30,54,31,54,30,157,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
