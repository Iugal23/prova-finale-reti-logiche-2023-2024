-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 678;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (11,0,223,0,129,0,0,0,30,0,190,0,90,0,39,0,62,0,83,0,172,0,0,0,108,0,0,0,186,0,0,0,0,0,110,0,113,0,6,0,159,0,211,0,78,0,29,0,224,0,0,0,107,0,116,0,238,0,246,0,0,0,0,0,224,0,79,0,195,0,0,0,82,0,0,0,224,0,0,0,241,0,53,0,67,0,79,0,0,0,139,0,91,0,0,0,0,0,17,0,219,0,243,0,131,0,0,0,0,0,86,0,0,0,190,0,112,0,171,0,95,0,233,0,133,0,169,0,101,0,3,0,0,0,0,0,177,0,244,0,119,0,0,0,100,0,8,0,54,0,244,0,138,0,162,0,0,0,0,0,193,0,208,0,196,0,0,0,96,0,0,0,0,0,0,0,99,0,114,0,37,0,114,0,171,0,74,0,182,0,0,0,41,0,142,0,1,0,45,0,181,0,162,0,0,0,0,0,169,0,70,0,119,0,190,0,0,0,246,0,41,0,195,0,123,0,57,0,153,0,0,0,141,0,104,0,177,0,131,0,104,0,206,0,226,0,147,0,38,0,39,0,184,0,108,0,136,0,0,0,234,0,54,0,206,0,163,0,0,0,8,0,78,0,0,0,0,0,38,0,152,0,150,0,89,0,133,0,127,0,0,0,195,0,18,0,218,0,60,0,195,0,165,0,0,0,75,0,232,0,236,0,144,0,98,0,0,0,84,0,167,0,0,0,26,0,82,0,172,0,31,0,197,0,0,0,0,0,0,0,123,0,58,0,0,0,249,0,0,0,138,0,86,0,0,0,126,0,249,0,192,0,107,0,40,0,79,0,58,0,155,0,0,0,46,0,0,0,229,0,0,0,248,0,232,0,66,0,19,0,248,0,119,0,0,0,176,0,129,0,34,0,205,0,0,0,0,0,179,0,42,0,194,0,174,0,181,0,107,0,232,0,0,0,223,0,148,0,101,0,178,0,46,0,228,0,211,0,0,0,196,0,19,0,192,0,30,0,183,0,94,0,0,0,93,0,0,0,24,0,13,0,116,0,136,0,45,0,173,0,0,0,87,0,114,0,152,0,154,0,73,0,190,0,0,0,50,0,114,0,0,0,216,0,204,0,31,0,174,0,58,0,158,0,136,0,92,0,0,0,242,0,101,0,124,0,182,0,0,0,82,0,152,0,156,0,0,0,252,0,0,0,0,0,0,0,48,0,225,0,130,0,50,0,135,0,241,0,0,0,0,0,217,0,74,0,35,0,78,0,0,0,168,0,216,0,0,0,219,0,72,0,144,0,7,0,101,0,38,0,215,0,227,0,3,0,0,0,124,0,208,0,239,0,196,0,159,0,147,0,239,0,0,0,35,0,233,0,180,0,227,0,5,0,225,0,78,0,245,0,211,0,220,0,128,0,172,0,0,0,153,0,147,0,86,0,10,0,166,0,0,0,231,0,0,0,255,0,159,0,9,0,65,0,196,0,115,0,0,0,40,0,198,0,97,0,108,0,8,0,108,0,217,0,144,0,130,0,108,0,68,0,55,0,139,0,227,0,148,0,181,0,138,0,103,0,63,0,138,0,0,0,201,0,19,0,0,0,31,0,156,0,169,0,195,0,33,0,0,0,54,0,10,0,224,0,0,0,125,0,126,0,0,0,232,0,0,0,199,0,232,0,251,0,0,0,44,0,152,0,15,0,0,0,156,0,47,0,0,0,236,0,0,0,36,0,116,0,176,0,201,0,0,0,250,0,0,0,66,0,139,0,0,0,31,0,127,0,102,0,0,0,207,0,234,0,186,0,104,0,135,0,75,0,164,0,34,0,202,0,162,0,86,0,52,0,73,0,238,0,207,0,199,0,19,0,44,0,0,0,248,0,85,0,122,0,36,0,157,0,28,0,197,0,136,0,116,0,0,0,78,0,0,0,60,0,0,0,66,0,93,0,186,0,99,0,232,0,0,0,224,0,0,0,0,0,226,0,238,0,51,0,188,0,71,0,163,0,68,0,112,0,0,0,35,0,29,0,190,0,187,0,188,0,36,0,116,0,48,0,147,0,39,0,181,0,61,0,98,0,0,0,0,0,46,0,0,0,84,0,52,0,0,0,234,0,86,0,203,0,150,0,80,0,240,0,178,0,27,0,144,0,162,0,59,0,116,0,30,0,126,0,132,0,0,0,99,0,134,0,217,0,242,0,101,0,5,0,234,0,82,0,124,0,144,0,0,0,28,0,0,0,197,0,226,0,177,0,84,0,124,0,144,0,0,0,0,0,39,0,131,0,0,0,114,0,15,0,0,0,30,0,194,0,0,0,41,0,216,0,134,0,234,0,86,0,54,0,196,0,0,0,8,0,10,0,80,0,194,0,0,0,0,0,0,0,104,0,166,0,43,0,206,0,6,0,108,0,0,0,218,0,213,0,61,0,116,0,163,0,0,0,235,0,0,0,31,0,50,0,0,0,210,0,57,0,116,0,197,0,0,0,129,0,232,0,163,0,144,0,0,0,131,0,135,0,112,0,0,0,102,0,138,0,0,0,147,0,131,0,130,0,124,0,198,0,195,0,101,0,226,0,6,0,0,0,80,0,184,0,46,0,17,0,223,0,44,0,107,0,123,0,108,0,134,0,80,0,0,0,236,0,102,0,0,0,107,0,147,0,0,0,182,0,192,0,24,0,0,0,155,0,207,0,80,0,71,0,160,0,10,0,0,0,191,0,73,0,236,0,167,0,0,0,212,0,222,0,0,0,129,0,0,0,1,0,0,0,234,0,151,0,154,0,196,0,0,0,213,0,58,0,127,0,207,0,0,0,56,0,219,0,244,0,117,0,49,0,178,0,118,0,183,0,217,0,254,0,0,0,136,0,99,0,8,0,30,0,175,0,0,0,239,0,0,0,0,0,135,0,83,0,47,0,0,0,191,0,0,0,0,0,0,0,87,0,175,0,204,0,195,0,85,0,147,0,0,0,13,0,164,0,213,0,83,0,154,0,0,0,58,0,142,0,64,0,0,0,38,0,199,0,125,0,78,0,204,0,39,0,173,0,222,0,0,0);
signal scenario_full  : scenario_type := (11,31,223,31,129,31,129,30,30,31,190,31,90,31,39,31,62,31,83,31,172,31,172,30,108,31,108,30,186,31,186,30,186,29,110,31,113,31,6,31,159,31,211,31,78,31,29,31,224,31,224,30,107,31,116,31,238,31,246,31,246,30,246,29,224,31,79,31,195,31,195,30,82,31,82,30,224,31,224,30,241,31,53,31,67,31,79,31,79,30,139,31,91,31,91,30,91,29,17,31,219,31,243,31,131,31,131,30,131,29,86,31,86,30,190,31,112,31,171,31,95,31,233,31,133,31,169,31,101,31,3,31,3,30,3,29,177,31,244,31,119,31,119,30,100,31,8,31,54,31,244,31,138,31,162,31,162,30,162,29,193,31,208,31,196,31,196,30,96,31,96,30,96,29,96,28,99,31,114,31,37,31,114,31,171,31,74,31,182,31,182,30,41,31,142,31,1,31,45,31,181,31,162,31,162,30,162,29,169,31,70,31,119,31,190,31,190,30,246,31,41,31,195,31,123,31,57,31,153,31,153,30,141,31,104,31,177,31,131,31,104,31,206,31,226,31,147,31,38,31,39,31,184,31,108,31,136,31,136,30,234,31,54,31,206,31,163,31,163,30,8,31,78,31,78,30,78,29,38,31,152,31,150,31,89,31,133,31,127,31,127,30,195,31,18,31,218,31,60,31,195,31,165,31,165,30,75,31,232,31,236,31,144,31,98,31,98,30,84,31,167,31,167,30,26,31,82,31,172,31,31,31,197,31,197,30,197,29,197,28,123,31,58,31,58,30,249,31,249,30,138,31,86,31,86,30,126,31,249,31,192,31,107,31,40,31,79,31,58,31,155,31,155,30,46,31,46,30,229,31,229,30,248,31,232,31,66,31,19,31,248,31,119,31,119,30,176,31,129,31,34,31,205,31,205,30,205,29,179,31,42,31,194,31,174,31,181,31,107,31,232,31,232,30,223,31,148,31,101,31,178,31,46,31,228,31,211,31,211,30,196,31,19,31,192,31,30,31,183,31,94,31,94,30,93,31,93,30,24,31,13,31,116,31,136,31,45,31,173,31,173,30,87,31,114,31,152,31,154,31,73,31,190,31,190,30,50,31,114,31,114,30,216,31,204,31,31,31,174,31,58,31,158,31,136,31,92,31,92,30,242,31,101,31,124,31,182,31,182,30,82,31,152,31,156,31,156,30,252,31,252,30,252,29,252,28,48,31,225,31,130,31,50,31,135,31,241,31,241,30,241,29,217,31,74,31,35,31,78,31,78,30,168,31,216,31,216,30,219,31,72,31,144,31,7,31,101,31,38,31,215,31,227,31,3,31,3,30,124,31,208,31,239,31,196,31,159,31,147,31,239,31,239,30,35,31,233,31,180,31,227,31,5,31,225,31,78,31,245,31,211,31,220,31,128,31,172,31,172,30,153,31,147,31,86,31,10,31,166,31,166,30,231,31,231,30,255,31,159,31,9,31,65,31,196,31,115,31,115,30,40,31,198,31,97,31,108,31,8,31,108,31,217,31,144,31,130,31,108,31,68,31,55,31,139,31,227,31,148,31,181,31,138,31,103,31,63,31,138,31,138,30,201,31,19,31,19,30,31,31,156,31,169,31,195,31,33,31,33,30,54,31,10,31,224,31,224,30,125,31,126,31,126,30,232,31,232,30,199,31,232,31,251,31,251,30,44,31,152,31,15,31,15,30,156,31,47,31,47,30,236,31,236,30,36,31,116,31,176,31,201,31,201,30,250,31,250,30,66,31,139,31,139,30,31,31,127,31,102,31,102,30,207,31,234,31,186,31,104,31,135,31,75,31,164,31,34,31,202,31,162,31,86,31,52,31,73,31,238,31,207,31,199,31,19,31,44,31,44,30,248,31,85,31,122,31,36,31,157,31,28,31,197,31,136,31,116,31,116,30,78,31,78,30,60,31,60,30,66,31,93,31,186,31,99,31,232,31,232,30,224,31,224,30,224,29,226,31,238,31,51,31,188,31,71,31,163,31,68,31,112,31,112,30,35,31,29,31,190,31,187,31,188,31,36,31,116,31,48,31,147,31,39,31,181,31,61,31,98,31,98,30,98,29,46,31,46,30,84,31,52,31,52,30,234,31,86,31,203,31,150,31,80,31,240,31,178,31,27,31,144,31,162,31,59,31,116,31,30,31,126,31,132,31,132,30,99,31,134,31,217,31,242,31,101,31,5,31,234,31,82,31,124,31,144,31,144,30,28,31,28,30,197,31,226,31,177,31,84,31,124,31,144,31,144,30,144,29,39,31,131,31,131,30,114,31,15,31,15,30,30,31,194,31,194,30,41,31,216,31,134,31,234,31,86,31,54,31,196,31,196,30,8,31,10,31,80,31,194,31,194,30,194,29,194,28,104,31,166,31,43,31,206,31,6,31,108,31,108,30,218,31,213,31,61,31,116,31,163,31,163,30,235,31,235,30,31,31,50,31,50,30,210,31,57,31,116,31,197,31,197,30,129,31,232,31,163,31,144,31,144,30,131,31,135,31,112,31,112,30,102,31,138,31,138,30,147,31,131,31,130,31,124,31,198,31,195,31,101,31,226,31,6,31,6,30,80,31,184,31,46,31,17,31,223,31,44,31,107,31,123,31,108,31,134,31,80,31,80,30,236,31,102,31,102,30,107,31,147,31,147,30,182,31,192,31,24,31,24,30,155,31,207,31,80,31,71,31,160,31,10,31,10,30,191,31,73,31,236,31,167,31,167,30,212,31,222,31,222,30,129,31,129,30,1,31,1,30,234,31,151,31,154,31,196,31,196,30,213,31,58,31,127,31,207,31,207,30,56,31,219,31,244,31,117,31,49,31,178,31,118,31,183,31,217,31,254,31,254,30,136,31,99,31,8,31,30,31,175,31,175,30,239,31,239,30,239,29,135,31,83,31,47,31,47,30,191,31,191,30,191,29,191,28,87,31,175,31,204,31,195,31,85,31,147,31,147,30,13,31,164,31,213,31,83,31,154,31,154,30,58,31,142,31,64,31,64,30,38,31,199,31,125,31,78,31,204,31,39,31,173,31,222,31,222,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
