-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 399;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,179,0,44,0,18,0,184,0,0,0,167,0,75,0,222,0,206,0,201,0,0,0,89,0,47,0,63,0,0,0,136,0,0,0,197,0,0,0,31,0,10,0,35,0,0,0,5,0,44,0,1,0,0,0,178,0,125,0,180,0,4,0,148,0,0,0,175,0,38,0,104,0,91,0,0,0,0,0,182,0,247,0,0,0,44,0,0,0,1,0,226,0,99,0,87,0,212,0,117,0,0,0,17,0,203,0,223,0,52,0,181,0,126,0,47,0,0,0,0,0,0,0,251,0,0,0,214,0,166,0,17,0,0,0,0,0,0,0,211,0,175,0,241,0,25,0,0,0,0,0,0,0,126,0,0,0,39,0,139,0,0,0,131,0,252,0,58,0,32,0,0,0,29,0,227,0,75,0,251,0,117,0,255,0,200,0,8,0,56,0,99,0,6,0,0,0,103,0,201,0,55,0,118,0,217,0,34,0,107,0,44,0,43,0,0,0,0,0,0,0,0,0,3,0,119,0,0,0,0,0,102,0,89,0,25,0,150,0,226,0,0,0,118,0,0,0,134,0,83,0,201,0,90,0,12,0,227,0,32,0,77,0,16,0,0,0,151,0,0,0,0,0,162,0,0,0,232,0,233,0,161,0,76,0,60,0,214,0,194,0,236,0,48,0,72,0,67,0,104,0,205,0,186,0,135,0,30,0,215,0,200,0,0,0,172,0,234,0,33,0,17,0,127,0,209,0,2,0,159,0,153,0,224,0,252,0,0,0,157,0,161,0,73,0,235,0,27,0,0,0,100,0,208,0,186,0,129,0,193,0,51,0,169,0,5,0,164,0,0,0,18,0,3,0,71,0,154,0,0,0,87,0,166,0,141,0,0,0,29,0,0,0,80,0,0,0,243,0,86,0,179,0,37,0,70,0,151,0,79,0,68,0,130,0,0,0,0,0,33,0,29,0,99,0,28,0,0,0,117,0,0,0,93,0,59,0,61,0,57,0,0,0,72,0,203,0,0,0,90,0,84,0,0,0,169,0,136,0,241,0,198,0,83,0,98,0,0,0,104,0,241,0,28,0,184,0,252,0,136,0,0,0,40,0,46,0,90,0,191,0,56,0,84,0,94,0,124,0,12,0,59,0,0,0,127,0,181,0,0,0,59,0,13,0,54,0,246,0,25,0,0,0,168,0,12,0,232,0,105,0,37,0,2,0,217,0,200,0,236,0,58,0,182,0,86,0,83,0,0,0,110,0,129,0,0,0,18,0,31,0,122,0,0,0,0,0,185,0,122,0,160,0,161,0,130,0,178,0,103,0,249,0,171,0,0,0,215,0,41,0,95,0,16,0,0,0,167,0,93,0,238,0,222,0,86,0,10,0,51,0,127,0,0,0,56,0,0,0,27,0,145,0,33,0,16,0,127,0,152,0,58,0,157,0,51,0,0,0,93,0,25,0,0,0,89,0,76,0,214,0,221,0,51,0,209,0,126,0,221,0,6,0,152,0,35,0,7,0,0,0,208,0,189,0,139,0,98,0,0,0,90,0,40,0,40,0,62,0,114,0,0,0,32,0,20,0,212,0,182,0,0,0,0,0,153,0,207,0,0,0,243,0,184,0,161,0,161,0,63,0,134,0,0,0,179,0,66,0,114,0,222,0,73,0,92,0,8,0,173,0,244,0,74,0,0,0,207,0,48,0,160,0,176,0,50,0,123,0,35,0,186,0,181,0,141,0,100,0,215,0,140,0,84,0,0,0,0,0,35,0,62,0,0,0,224,0,240,0,0,0,221,0,165,0,14,0);
signal scenario_full  : scenario_type := (0,0,179,31,44,31,18,31,184,31,184,30,167,31,75,31,222,31,206,31,201,31,201,30,89,31,47,31,63,31,63,30,136,31,136,30,197,31,197,30,31,31,10,31,35,31,35,30,5,31,44,31,1,31,1,30,178,31,125,31,180,31,4,31,148,31,148,30,175,31,38,31,104,31,91,31,91,30,91,29,182,31,247,31,247,30,44,31,44,30,1,31,226,31,99,31,87,31,212,31,117,31,117,30,17,31,203,31,223,31,52,31,181,31,126,31,47,31,47,30,47,29,47,28,251,31,251,30,214,31,166,31,17,31,17,30,17,29,17,28,211,31,175,31,241,31,25,31,25,30,25,29,25,28,126,31,126,30,39,31,139,31,139,30,131,31,252,31,58,31,32,31,32,30,29,31,227,31,75,31,251,31,117,31,255,31,200,31,8,31,56,31,99,31,6,31,6,30,103,31,201,31,55,31,118,31,217,31,34,31,107,31,44,31,43,31,43,30,43,29,43,28,43,27,3,31,119,31,119,30,119,29,102,31,89,31,25,31,150,31,226,31,226,30,118,31,118,30,134,31,83,31,201,31,90,31,12,31,227,31,32,31,77,31,16,31,16,30,151,31,151,30,151,29,162,31,162,30,232,31,233,31,161,31,76,31,60,31,214,31,194,31,236,31,48,31,72,31,67,31,104,31,205,31,186,31,135,31,30,31,215,31,200,31,200,30,172,31,234,31,33,31,17,31,127,31,209,31,2,31,159,31,153,31,224,31,252,31,252,30,157,31,161,31,73,31,235,31,27,31,27,30,100,31,208,31,186,31,129,31,193,31,51,31,169,31,5,31,164,31,164,30,18,31,3,31,71,31,154,31,154,30,87,31,166,31,141,31,141,30,29,31,29,30,80,31,80,30,243,31,86,31,179,31,37,31,70,31,151,31,79,31,68,31,130,31,130,30,130,29,33,31,29,31,99,31,28,31,28,30,117,31,117,30,93,31,59,31,61,31,57,31,57,30,72,31,203,31,203,30,90,31,84,31,84,30,169,31,136,31,241,31,198,31,83,31,98,31,98,30,104,31,241,31,28,31,184,31,252,31,136,31,136,30,40,31,46,31,90,31,191,31,56,31,84,31,94,31,124,31,12,31,59,31,59,30,127,31,181,31,181,30,59,31,13,31,54,31,246,31,25,31,25,30,168,31,12,31,232,31,105,31,37,31,2,31,217,31,200,31,236,31,58,31,182,31,86,31,83,31,83,30,110,31,129,31,129,30,18,31,31,31,122,31,122,30,122,29,185,31,122,31,160,31,161,31,130,31,178,31,103,31,249,31,171,31,171,30,215,31,41,31,95,31,16,31,16,30,167,31,93,31,238,31,222,31,86,31,10,31,51,31,127,31,127,30,56,31,56,30,27,31,145,31,33,31,16,31,127,31,152,31,58,31,157,31,51,31,51,30,93,31,25,31,25,30,89,31,76,31,214,31,221,31,51,31,209,31,126,31,221,31,6,31,152,31,35,31,7,31,7,30,208,31,189,31,139,31,98,31,98,30,90,31,40,31,40,31,62,31,114,31,114,30,32,31,20,31,212,31,182,31,182,30,182,29,153,31,207,31,207,30,243,31,184,31,161,31,161,31,63,31,134,31,134,30,179,31,66,31,114,31,222,31,73,31,92,31,8,31,173,31,244,31,74,31,74,30,207,31,48,31,160,31,176,31,50,31,123,31,35,31,186,31,181,31,141,31,100,31,215,31,140,31,84,31,84,30,84,29,35,31,62,31,62,30,224,31,240,31,240,30,221,31,165,31,14,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
