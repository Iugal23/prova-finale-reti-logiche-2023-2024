-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 708;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (69,0,0,0,49,0,1,0,189,0,69,0,162,0,0,0,52,0,0,0,245,0,181,0,22,0,0,0,0,0,237,0,11,0,199,0,241,0,26,0,166,0,69,0,0,0,0,0,92,0,117,0,87,0,211,0,0,0,172,0,0,0,0,0,217,0,0,0,0,0,193,0,52,0,131,0,219,0,57,0,28,0,211,0,143,0,37,0,0,0,46,0,98,0,81,0,28,0,0,0,175,0,15,0,0,0,124,0,172,0,20,0,129,0,0,0,209,0,0,0,193,0,0,0,242,0,213,0,185,0,232,0,135,0,199,0,0,0,0,0,61,0,0,0,95,0,0,0,223,0,222,0,55,0,83,0,13,0,57,0,235,0,30,0,200,0,89,0,208,0,113,0,0,0,0,0,39,0,134,0,0,0,74,0,0,0,173,0,83,0,247,0,176,0,175,0,0,0,173,0,246,0,242,0,126,0,253,0,0,0,78,0,0,0,185,0,197,0,137,0,45,0,80,0,204,0,31,0,0,0,33,0,64,0,150,0,101,0,83,0,92,0,117,0,0,0,113,0,25,0,147,0,192,0,72,0,8,0,208,0,38,0,0,0,245,0,153,0,88,0,31,0,0,0,113,0,0,0,41,0,252,0,0,0,98,0,202,0,176,0,240,0,100,0,160,0,7,0,181,0,157,0,223,0,27,0,91,0,142,0,11,0,177,0,31,0,253,0,0,0,129,0,12,0,23,0,0,0,92,0,80,0,0,0,0,0,161,0,0,0,193,0,153,0,191,0,35,0,167,0,190,0,231,0,146,0,54,0,229,0,0,0,45,0,187,0,152,0,133,0,39,0,0,0,200,0,82,0,0,0,5,0,89,0,6,0,124,0,52,0,5,0,65,0,251,0,9,0,119,0,248,0,0,0,44,0,0,0,0,0,168,0,131,0,0,0,110,0,0,0,146,0,185,0,50,0,0,0,110,0,0,0,128,0,71,0,129,0,251,0,0,0,222,0,206,0,174,0,184,0,224,0,192,0,0,0,96,0,64,0,0,0,66,0,127,0,208,0,133,0,0,0,79,0,0,0,197,0,51,0,0,0,108,0,196,0,215,0,92,0,219,0,250,0,222,0,151,0,96,0,235,0,206,0,0,0,200,0,78,0,252,0,0,0,75,0,177,0,51,0,96,0,0,0,205,0,110,0,105,0,83,0,40,0,206,0,0,0,50,0,41,0,31,0,0,0,146,0,182,0,38,0,244,0,9,0,172,0,62,0,127,0,253,0,205,0,194,0,0,0,0,0,150,0,0,0,65,0,17,0,65,0,122,0,243,0,109,0,199,0,196,0,130,0,111,0,0,0,75,0,22,0,153,0,2,0,92,0,230,0,180,0,185,0,19,0,243,0,162,0,0,0,219,0,115,0,210,0,119,0,77,0,0,0,233,0,226,0,64,0,136,0,112,0,32,0,74,0,83,0,240,0,142,0,48,0,14,0,236,0,172,0,0,0,124,0,0,0,106,0,229,0,25,0,83,0,144,0,162,0,0,0,37,0,236,0,248,0,74,0,167,0,0,0,0,0,169,0,103,0,243,0,56,0,238,0,115,0,58,0,248,0,190,0,0,0,6,0,229,0,88,0,209,0,152,0,0,0,183,0,213,0,143,0,253,0,0,0,148,0,73,0,214,0,0,0,79,0,4,0,26,0,18,0,47,0,81,0,147,0,51,0,81,0,149,0,80,0,255,0,240,0,23,0,32,0,223,0,220,0,195,0,32,0,67,0,191,0,255,0,216,0,180,0,0,0,162,0,0,0,11,0,47,0,0,0,145,0,12,0,121,0,0,0,80,0,165,0,91,0,18,0,147,0,0,0,144,0,132,0,21,0,150,0,176,0,236,0,161,0,217,0,94,0,140,0,0,0,30,0,14,0,0,0,194,0,9,0,0,0,0,0,0,0,242,0,90,0,179,0,48,0,149,0,136,0,93,0,246,0,165,0,161,0,0,0,197,0,0,0,139,0,5,0,159,0,0,0,0,0,3,0,220,0,182,0,127,0,166,0,111,0,191,0,205,0,181,0,234,0,52,0,148,0,207,0,115,0,0,0,4,0,149,0,85,0,138,0,83,0,13,0,229,0,0,0,151,0,0,0,178,0,131,0,93,0,1,0,60,0,210,0,253,0,206,0,218,0,0,0,208,0,227,0,164,0,216,0,151,0,0,0,232,0,221,0,0,0,0,0,129,0,217,0,225,0,136,0,176,0,0,0,0,0,0,0,248,0,34,0,253,0,88,0,81,0,154,0,17,0,0,0,16,0,60,0,114,0,134,0,57,0,59,0,190,0,206,0,164,0,206,0,160,0,248,0,236,0,126,0,188,0,83,0,53,0,86,0,0,0,74,0,40,0,210,0,255,0,206,0,37,0,210,0,60,0,101,0,205,0,0,0,0,0,0,0,2,0,120,0,142,0,192,0,57,0,158,0,154,0,204,0,26,0,119,0,56,0,2,0,0,0,0,0,73,0,0,0,0,0,154,0,86,0,120,0,13,0,98,0,231,0,0,0,145,0,87,0,203,0,80,0,198,0,78,0,87,0,139,0,0,0,0,0,54,0,229,0,44,0,2,0,0,0,206,0,206,0,137,0,166,0,46,0,72,0,158,0,17,0,173,0,188,0,0,0,0,0,228,0,43,0,76,0,84,0,50,0,23,0,0,0,186,0,156,0,0,0,103,0,100,0,18,0,158,0,38,0,0,0,46,0,4,0,104,0,46,0,207,0,104,0,140,0,85,0,35,0,71,0,143,0,201,0,184,0,58,0,9,0,201,0,0,0,121,0,113,0,13,0,142,0,0,0,163,0,161,0,0,0,190,0,193,0,179,0,0,0,0,0,205,0,0,0,222,0,0,0,3,0,89,0,209,0,0,0,119,0,142,0,145,0,0,0,194,0,0,0,239,0,48,0,208,0,160,0,0,0,133,0,73,0,82,0,74,0,47,0,34,0,0,0,232,0,0,0,66,0,0,0,17,0,134,0,207,0,7,0,86,0,73,0,66,0,0,0,0,0,0,0,255,0,148,0,172,0,0,0,9,0,47,0,213,0,252,0,114,0,0,0,169,0,180,0,88,0,243,0,253,0,248,0,79,0,0,0,116,0,4,0,183,0,134,0,19,0,183,0,0,0,199,0,0,0,183,0);
signal scenario_full  : scenario_type := (69,31,69,30,49,31,1,31,189,31,69,31,162,31,162,30,52,31,52,30,245,31,181,31,22,31,22,30,22,29,237,31,11,31,199,31,241,31,26,31,166,31,69,31,69,30,69,29,92,31,117,31,87,31,211,31,211,30,172,31,172,30,172,29,217,31,217,30,217,29,193,31,52,31,131,31,219,31,57,31,28,31,211,31,143,31,37,31,37,30,46,31,98,31,81,31,28,31,28,30,175,31,15,31,15,30,124,31,172,31,20,31,129,31,129,30,209,31,209,30,193,31,193,30,242,31,213,31,185,31,232,31,135,31,199,31,199,30,199,29,61,31,61,30,95,31,95,30,223,31,222,31,55,31,83,31,13,31,57,31,235,31,30,31,200,31,89,31,208,31,113,31,113,30,113,29,39,31,134,31,134,30,74,31,74,30,173,31,83,31,247,31,176,31,175,31,175,30,173,31,246,31,242,31,126,31,253,31,253,30,78,31,78,30,185,31,197,31,137,31,45,31,80,31,204,31,31,31,31,30,33,31,64,31,150,31,101,31,83,31,92,31,117,31,117,30,113,31,25,31,147,31,192,31,72,31,8,31,208,31,38,31,38,30,245,31,153,31,88,31,31,31,31,30,113,31,113,30,41,31,252,31,252,30,98,31,202,31,176,31,240,31,100,31,160,31,7,31,181,31,157,31,223,31,27,31,91,31,142,31,11,31,177,31,31,31,253,31,253,30,129,31,12,31,23,31,23,30,92,31,80,31,80,30,80,29,161,31,161,30,193,31,153,31,191,31,35,31,167,31,190,31,231,31,146,31,54,31,229,31,229,30,45,31,187,31,152,31,133,31,39,31,39,30,200,31,82,31,82,30,5,31,89,31,6,31,124,31,52,31,5,31,65,31,251,31,9,31,119,31,248,31,248,30,44,31,44,30,44,29,168,31,131,31,131,30,110,31,110,30,146,31,185,31,50,31,50,30,110,31,110,30,128,31,71,31,129,31,251,31,251,30,222,31,206,31,174,31,184,31,224,31,192,31,192,30,96,31,64,31,64,30,66,31,127,31,208,31,133,31,133,30,79,31,79,30,197,31,51,31,51,30,108,31,196,31,215,31,92,31,219,31,250,31,222,31,151,31,96,31,235,31,206,31,206,30,200,31,78,31,252,31,252,30,75,31,177,31,51,31,96,31,96,30,205,31,110,31,105,31,83,31,40,31,206,31,206,30,50,31,41,31,31,31,31,30,146,31,182,31,38,31,244,31,9,31,172,31,62,31,127,31,253,31,205,31,194,31,194,30,194,29,150,31,150,30,65,31,17,31,65,31,122,31,243,31,109,31,199,31,196,31,130,31,111,31,111,30,75,31,22,31,153,31,2,31,92,31,230,31,180,31,185,31,19,31,243,31,162,31,162,30,219,31,115,31,210,31,119,31,77,31,77,30,233,31,226,31,64,31,136,31,112,31,32,31,74,31,83,31,240,31,142,31,48,31,14,31,236,31,172,31,172,30,124,31,124,30,106,31,229,31,25,31,83,31,144,31,162,31,162,30,37,31,236,31,248,31,74,31,167,31,167,30,167,29,169,31,103,31,243,31,56,31,238,31,115,31,58,31,248,31,190,31,190,30,6,31,229,31,88,31,209,31,152,31,152,30,183,31,213,31,143,31,253,31,253,30,148,31,73,31,214,31,214,30,79,31,4,31,26,31,18,31,47,31,81,31,147,31,51,31,81,31,149,31,80,31,255,31,240,31,23,31,32,31,223,31,220,31,195,31,32,31,67,31,191,31,255,31,216,31,180,31,180,30,162,31,162,30,11,31,47,31,47,30,145,31,12,31,121,31,121,30,80,31,165,31,91,31,18,31,147,31,147,30,144,31,132,31,21,31,150,31,176,31,236,31,161,31,217,31,94,31,140,31,140,30,30,31,14,31,14,30,194,31,9,31,9,30,9,29,9,28,242,31,90,31,179,31,48,31,149,31,136,31,93,31,246,31,165,31,161,31,161,30,197,31,197,30,139,31,5,31,159,31,159,30,159,29,3,31,220,31,182,31,127,31,166,31,111,31,191,31,205,31,181,31,234,31,52,31,148,31,207,31,115,31,115,30,4,31,149,31,85,31,138,31,83,31,13,31,229,31,229,30,151,31,151,30,178,31,131,31,93,31,1,31,60,31,210,31,253,31,206,31,218,31,218,30,208,31,227,31,164,31,216,31,151,31,151,30,232,31,221,31,221,30,221,29,129,31,217,31,225,31,136,31,176,31,176,30,176,29,176,28,248,31,34,31,253,31,88,31,81,31,154,31,17,31,17,30,16,31,60,31,114,31,134,31,57,31,59,31,190,31,206,31,164,31,206,31,160,31,248,31,236,31,126,31,188,31,83,31,53,31,86,31,86,30,74,31,40,31,210,31,255,31,206,31,37,31,210,31,60,31,101,31,205,31,205,30,205,29,205,28,2,31,120,31,142,31,192,31,57,31,158,31,154,31,204,31,26,31,119,31,56,31,2,31,2,30,2,29,73,31,73,30,73,29,154,31,86,31,120,31,13,31,98,31,231,31,231,30,145,31,87,31,203,31,80,31,198,31,78,31,87,31,139,31,139,30,139,29,54,31,229,31,44,31,2,31,2,30,206,31,206,31,137,31,166,31,46,31,72,31,158,31,17,31,173,31,188,31,188,30,188,29,228,31,43,31,76,31,84,31,50,31,23,31,23,30,186,31,156,31,156,30,103,31,100,31,18,31,158,31,38,31,38,30,46,31,4,31,104,31,46,31,207,31,104,31,140,31,85,31,35,31,71,31,143,31,201,31,184,31,58,31,9,31,201,31,201,30,121,31,113,31,13,31,142,31,142,30,163,31,161,31,161,30,190,31,193,31,179,31,179,30,179,29,205,31,205,30,222,31,222,30,3,31,89,31,209,31,209,30,119,31,142,31,145,31,145,30,194,31,194,30,239,31,48,31,208,31,160,31,160,30,133,31,73,31,82,31,74,31,47,31,34,31,34,30,232,31,232,30,66,31,66,30,17,31,134,31,207,31,7,31,86,31,73,31,66,31,66,30,66,29,66,28,255,31,148,31,172,31,172,30,9,31,47,31,213,31,252,31,114,31,114,30,169,31,180,31,88,31,243,31,253,31,248,31,79,31,79,30,116,31,4,31,183,31,134,31,19,31,183,31,183,30,199,31,199,30,183,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
