-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_325 is
end project_tb_325;

architecture project_tb_arch_325 of project_tb_325 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 329;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,122,0,0,0,81,0,0,0,0,0,250,0,80,0,198,0,129,0,195,0,233,0,236,0,72,0,127,0,68,0,0,0,75,0,142,0,108,0,204,0,0,0,0,0,26,0,182,0,46,0,111,0,176,0,0,0,0,0,55,0,191,0,210,0,0,0,234,0,119,0,28,0,0,0,232,0,125,0,76,0,117,0,0,0,159,0,222,0,142,0,80,0,4,0,0,0,235,0,119,0,203,0,230,0,147,0,0,0,211,0,57,0,169,0,245,0,169,0,82,0,76,0,93,0,161,0,0,0,0,0,84,0,116,0,99,0,237,0,209,0,0,0,168,0,109,0,61,0,153,0,147,0,0,0,226,0,108,0,158,0,33,0,164,0,0,0,0,0,36,0,41,0,5,0,206,0,0,0,54,0,98,0,54,0,0,0,218,0,162,0,70,0,250,0,156,0,0,0,59,0,205,0,174,0,138,0,67,0,0,0,19,0,0,0,104,0,107,0,0,0,140,0,255,0,18,0,220,0,144,0,73,0,15,0,117,0,136,0,192,0,215,0,106,0,124,0,0,0,208,0,2,0,0,0,23,0,143,0,222,0,150,0,126,0,0,0,67,0,161,0,115,0,42,0,53,0,85,0,157,0,0,0,122,0,219,0,68,0,165,0,146,0,0,0,85,0,139,0,36,0,1,0,0,0,207,0,233,0,144,0,99,0,0,0,149,0,0,0,217,0,247,0,0,0,0,0,15,0,240,0,109,0,0,0,0,0,68,0,0,0,63,0,52,0,20,0,218,0,191,0,156,0,0,0,14,0,203,0,239,0,218,0,0,0,0,0,237,0,128,0,228,0,226,0,0,0,172,0,21,0,161,0,241,0,0,0,204,0,0,0,127,0,0,0,0,0,123,0,72,0,174,0,185,0,0,0,0,0,120,0,69,0,0,0,160,0,117,0,0,0,0,0,252,0,0,0,150,0,30,0,0,0,150,0,113,0,0,0,20,0,0,0,104,0,0,0,207,0,0,0,115,0,235,0,121,0,104,0,208,0,31,0,169,0,207,0,122,0,77,0,99,0,233,0,30,0,251,0,230,0,0,0,161,0,200,0,92,0,0,0,15,0,0,0,213,0,0,0,131,0,75,0,244,0,213,0,253,0,0,0,0,0,4,0,30,0,213,0,200,0,3,0,253,0,95,0,108,0,0,0,93,0,144,0,103,0,171,0,164,0,67,0,204,0,194,0,22,0,0,0,132,0,177,0,83,0,203,0,131,0,0,0,114,0,170,0,149,0,151,0,0,0,0,0,57,0,218,0,0,0,98,0,253,0,112,0,109,0,167,0,202,0,132,0,0,0,52,0,253,0,0,0,15,0,216,0,0,0,70,0,142,0,241,0,0,0,78,0,0,0,84,0,73,0,12,0,0,0,0,0,234,0,0,0,43,0,47,0,0,0,0,0,231,0,148,0,0,0,0,0,153,0,231,0,203,0);
signal scenario_full  : scenario_type := (0,0,122,31,122,30,81,31,81,30,81,29,250,31,80,31,198,31,129,31,195,31,233,31,236,31,72,31,127,31,68,31,68,30,75,31,142,31,108,31,204,31,204,30,204,29,26,31,182,31,46,31,111,31,176,31,176,30,176,29,55,31,191,31,210,31,210,30,234,31,119,31,28,31,28,30,232,31,125,31,76,31,117,31,117,30,159,31,222,31,142,31,80,31,4,31,4,30,235,31,119,31,203,31,230,31,147,31,147,30,211,31,57,31,169,31,245,31,169,31,82,31,76,31,93,31,161,31,161,30,161,29,84,31,116,31,99,31,237,31,209,31,209,30,168,31,109,31,61,31,153,31,147,31,147,30,226,31,108,31,158,31,33,31,164,31,164,30,164,29,36,31,41,31,5,31,206,31,206,30,54,31,98,31,54,31,54,30,218,31,162,31,70,31,250,31,156,31,156,30,59,31,205,31,174,31,138,31,67,31,67,30,19,31,19,30,104,31,107,31,107,30,140,31,255,31,18,31,220,31,144,31,73,31,15,31,117,31,136,31,192,31,215,31,106,31,124,31,124,30,208,31,2,31,2,30,23,31,143,31,222,31,150,31,126,31,126,30,67,31,161,31,115,31,42,31,53,31,85,31,157,31,157,30,122,31,219,31,68,31,165,31,146,31,146,30,85,31,139,31,36,31,1,31,1,30,207,31,233,31,144,31,99,31,99,30,149,31,149,30,217,31,247,31,247,30,247,29,15,31,240,31,109,31,109,30,109,29,68,31,68,30,63,31,52,31,20,31,218,31,191,31,156,31,156,30,14,31,203,31,239,31,218,31,218,30,218,29,237,31,128,31,228,31,226,31,226,30,172,31,21,31,161,31,241,31,241,30,204,31,204,30,127,31,127,30,127,29,123,31,72,31,174,31,185,31,185,30,185,29,120,31,69,31,69,30,160,31,117,31,117,30,117,29,252,31,252,30,150,31,30,31,30,30,150,31,113,31,113,30,20,31,20,30,104,31,104,30,207,31,207,30,115,31,235,31,121,31,104,31,208,31,31,31,169,31,207,31,122,31,77,31,99,31,233,31,30,31,251,31,230,31,230,30,161,31,200,31,92,31,92,30,15,31,15,30,213,31,213,30,131,31,75,31,244,31,213,31,253,31,253,30,253,29,4,31,30,31,213,31,200,31,3,31,253,31,95,31,108,31,108,30,93,31,144,31,103,31,171,31,164,31,67,31,204,31,194,31,22,31,22,30,132,31,177,31,83,31,203,31,131,31,131,30,114,31,170,31,149,31,151,31,151,30,151,29,57,31,218,31,218,30,98,31,253,31,112,31,109,31,167,31,202,31,132,31,132,30,52,31,253,31,253,30,15,31,216,31,216,30,70,31,142,31,241,31,241,30,78,31,78,30,84,31,73,31,12,31,12,30,12,29,234,31,234,30,43,31,47,31,47,30,47,29,231,31,148,31,148,30,148,29,153,31,231,31,203,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
