-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_344 is
end project_tb_344;

architecture project_tb_arch_344 of project_tb_344 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 941;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (44,0,0,0,145,0,9,0,135,0,127,0,0,0,54,0,139,0,0,0,199,0,197,0,94,0,129,0,0,0,0,0,0,0,195,0,0,0,0,0,190,0,96,0,83,0,14,0,111,0,159,0,0,0,3,0,107,0,228,0,113,0,26,0,0,0,96,0,45,0,110,0,213,0,0,0,0,0,81,0,0,0,26,0,110,0,120,0,148,0,159,0,118,0,20,0,214,0,12,0,231,0,8,0,186,0,182,0,87,0,165,0,203,0,0,0,151,0,173,0,217,0,56,0,0,0,160,0,173,0,30,0,118,0,171,0,126,0,54,0,214,0,189,0,0,0,138,0,34,0,136,0,236,0,145,0,205,0,117,0,138,0,48,0,0,0,51,0,0,0,213,0,0,0,251,0,0,0,228,0,27,0,226,0,243,0,20,0,83,0,16,0,0,0,175,0,0,0,69,0,35,0,231,0,163,0,0,0,162,0,49,0,0,0,207,0,167,0,123,0,0,0,52,0,40,0,198,0,0,0,169,0,94,0,0,0,0,0,0,0,0,0,24,0,111,0,201,0,198,0,0,0,32,0,0,0,1,0,49,0,0,0,84,0,50,0,0,0,50,0,252,0,0,0,158,0,76,0,10,0,195,0,131,0,193,0,73,0,97,0,7,0,19,0,0,0,61,0,98,0,0,0,35,0,0,0,0,0,6,0,159,0,196,0,0,0,198,0,200,0,0,0,0,0,128,0,93,0,182,0,231,0,117,0,160,0,2,0,226,0,0,0,137,0,26,0,162,0,255,0,64,0,17,0,42,0,205,0,175,0,76,0,3,0,0,0,0,0,227,0,16,0,130,0,0,0,0,0,0,0,0,0,0,0,164,0,8,0,184,0,0,0,217,0,10,0,222,0,0,0,195,0,157,0,217,0,61,0,231,0,44,0,124,0,20,0,0,0,222,0,65,0,251,0,193,0,216,0,54,0,224,0,46,0,0,0,137,0,198,0,250,0,127,0,46,0,170,0,203,0,0,0,19,0,69,0,175,0,0,0,21,0,221,0,147,0,74,0,0,0,0,0,146,0,155,0,122,0,69,0,91,0,0,0,116,0,0,0,0,0,185,0,121,0,149,0,77,0,226,0,240,0,0,0,0,0,177,0,60,0,133,0,0,0,74,0,224,0,103,0,152,0,58,0,164,0,0,0,225,0,63,0,101,0,145,0,7,0,0,0,24,0,0,0,253,0,175,0,105,0,0,0,41,0,61,0,148,0,92,0,22,0,174,0,229,0,179,0,187,0,66,0,67,0,102,0,122,0,0,0,182,0,189,0,214,0,222,0,157,0,12,0,217,0,0,0,0,0,25,0,50,0,254,0,61,0,34,0,222,0,181,0,15,0,93,0,143,0,22,0,0,0,28,0,68,0,133,0,0,0,184,0,11,0,171,0,225,0,0,0,55,0,20,0,133,0,199,0,184,0,0,0,181,0,78,0,49,0,62,0,84,0,0,0,0,0,51,0,252,0,124,0,39,0,0,0,245,0,208,0,243,0,152,0,65,0,91,0,86,0,55,0,43,0,8,0,14,0,151,0,101,0,197,0,0,0,154,0,0,0,95,0,0,0,254,0,253,0,0,0,211,0,0,0,21,0,180,0,147,0,0,0,37,0,114,0,100,0,243,0,252,0,39,0,47,0,4,0,66,0,229,0,85,0,211,0,225,0,64,0,234,0,151,0,76,0,0,0,249,0,125,0,190,0,112,0,0,0,0,0,100,0,145,0,242,0,0,0,195,0,62,0,55,0,80,0,80,0,148,0,0,0,171,0,0,0,218,0,0,0,0,0,121,0,233,0,0,0,18,0,100,0,56,0,13,0,75,0,236,0,14,0,157,0,119,0,213,0,0,0,102,0,161,0,115,0,66,0,133,0,0,0,179,0,196,0,16,0,61,0,0,0,77,0,38,0,172,0,0,0,108,0,0,0,221,0,190,0,148,0,26,0,33,0,125,0,19,0,59,0,131,0,234,0,112,0,84,0,0,0,90,0,44,0,0,0,243,0,85,0,73,0,159,0,84,0,253,0,221,0,213,0,106,0,211,0,184,0,118,0,50,0,222,0,2,0,95,0,23,0,65,0,143,0,0,0,85,0,0,0,0,0,233,0,231,0,53,0,68,0,39,0,213,0,107,0,127,0,126,0,164,0,241,0,78,0,58,0,0,0,0,0,164,0,254,0,118,0,19,0,249,0,79,0,117,0,52,0,133,0,198,0,0,0,0,0,20,0,34,0,217,0,110,0,13,0,0,0,181,0,242,0,83,0,0,0,120,0,58,0,131,0,243,0,151,0,0,0,10,0,51,0,0,0,0,0,0,0,18,0,241,0,107,0,103,0,64,0,167,0,174,0,224,0,0,0,0,0,214,0,78,0,0,0,186,0,155,0,79,0,88,0,0,0,5,0,0,0,133,0,0,0,0,0,10,0,13,0,197,0,244,0,187,0,23,0,0,0,0,0,253,0,123,0,231,0,41,0,224,0,0,0,182,0,0,0,100,0,156,0,34,0,37,0,0,0,0,0,17,0,182,0,0,0,99,0,5,0,173,0,241,0,164,0,224,0,90,0,1,0,123,0,152,0,121,0,91,0,166,0,0,0,17,0,0,0,255,0,0,0,75,0,77,0,99,0,30,0,228,0,239,0,213,0,35,0,139,0,55,0,222,0,208,0,135,0,9,0,95,0,121,0,145,0,226,0,100,0,83,0,202,0,37,0,224,0,67,0,41,0,177,0,139,0,181,0,59,0,21,0,212,0,175,0,245,0,0,0,118,0,0,0,108,0,220,0,240,0,0,0,240,0,55,0,140,0,170,0,0,0,140,0,33,0,152,0,0,0,233,0,124,0,158,0,68,0,241,0,207,0,112,0,42,0,1,0,0,0,55,0,152,0,46,0,139,0,0,0,187,0,17,0,178,0,181,0,94,0,141,0,149,0,0,0,4,0,0,0,47,0,0,0,0,0,117,0,62,0,0,0,81,0,219,0,125,0,176,0,118,0,0,0,3,0,116,0,48,0,22,0,51,0,105,0,73,0,98,0,215,0,109,0,173,0,76,0,114,0,188,0,75,0,0,0,26,0,155,0,242,0,144,0,0,0,216,0,8,0,165,0,42,0,157,0,84,0,159,0,66,0,80,0,63,0,7,0,234,0,94,0,217,0,0,0,0,0,131,0,223,0,175,0,240,0,181,0,0,0,209,0,224,0,41,0,0,0,240,0,132,0,182,0,145,0,140,0,0,0,110,0,76,0,25,0,0,0,45,0,184,0,60,0,59,0,124,0,37,0,226,0,240,0,147,0,87,0,135,0,202,0,171,0,158,0,96,0,19,0,238,0,63,0,0,0,0,0,18,0,107,0,192,0,148,0,0,0,194,0,201,0,0,0,149,0,211,0,0,0,222,0,47,0,84,0,195,0,18,0,0,0,0,0,0,0,92,0,0,0,87,0,148,0,124,0,0,0,125,0,170,0,248,0,209,0,98,0,239,0,203,0,118,0,243,0,0,0,235,0,149,0,223,0,243,0,101,0,126,0,203,0,175,0,55,0,0,0,0,0,59,0,0,0,0,0,149,0,141,0,20,0,49,0,218,0,248,0,82,0,143,0,85,0,36,0,0,0,159,0,7,0,208,0,27,0,65,0,81,0,195,0,248,0,77,0,0,0,54,0,231,0,74,0,96,0,93,0,0,0,67,0,0,0,138,0,34,0,185,0,0,0,211,0,51,0,126,0,203,0,0,0,108,0,173,0,213,0,222,0,161,0,0,0,164,0,0,0,149,0,0,0,0,0,245,0,46,0,42,0,0,0,32,0,172,0,132,0,164,0,159,0,52,0,0,0,169,0,35,0,109,0,152,0,0,0,207,0,84,0,65,0,79,0,185,0,151,0,157,0,0,0,144,0,47,0,142,0,0,0,1,0,141,0,0,0,236,0,41,0,0,0,29,0,0,0,15,0,53,0,175,0,108,0,75,0,0,0,4,0,0,0,223,0,39,0,137,0,42,0,252,0,0,0,0,0,205,0,76,0,239,0,18,0,238,0,176,0,0,0,66,0,119,0,194,0,182,0,102,0,159,0,0,0,65,0,0,0,169,0,130,0,134,0,10,0,212,0,5,0,72,0,180,0,177,0,106,0,42,0,0,0,174,0,236,0,56,0,58,0,243,0,216,0,0,0,211,0,62,0,32,0,0,0);
signal scenario_full  : scenario_type := (44,31,44,30,145,31,9,31,135,31,127,31,127,30,54,31,139,31,139,30,199,31,197,31,94,31,129,31,129,30,129,29,129,28,195,31,195,30,195,29,190,31,96,31,83,31,14,31,111,31,159,31,159,30,3,31,107,31,228,31,113,31,26,31,26,30,96,31,45,31,110,31,213,31,213,30,213,29,81,31,81,30,26,31,110,31,120,31,148,31,159,31,118,31,20,31,214,31,12,31,231,31,8,31,186,31,182,31,87,31,165,31,203,31,203,30,151,31,173,31,217,31,56,31,56,30,160,31,173,31,30,31,118,31,171,31,126,31,54,31,214,31,189,31,189,30,138,31,34,31,136,31,236,31,145,31,205,31,117,31,138,31,48,31,48,30,51,31,51,30,213,31,213,30,251,31,251,30,228,31,27,31,226,31,243,31,20,31,83,31,16,31,16,30,175,31,175,30,69,31,35,31,231,31,163,31,163,30,162,31,49,31,49,30,207,31,167,31,123,31,123,30,52,31,40,31,198,31,198,30,169,31,94,31,94,30,94,29,94,28,94,27,24,31,111,31,201,31,198,31,198,30,32,31,32,30,1,31,49,31,49,30,84,31,50,31,50,30,50,31,252,31,252,30,158,31,76,31,10,31,195,31,131,31,193,31,73,31,97,31,7,31,19,31,19,30,61,31,98,31,98,30,35,31,35,30,35,29,6,31,159,31,196,31,196,30,198,31,200,31,200,30,200,29,128,31,93,31,182,31,231,31,117,31,160,31,2,31,226,31,226,30,137,31,26,31,162,31,255,31,64,31,17,31,42,31,205,31,175,31,76,31,3,31,3,30,3,29,227,31,16,31,130,31,130,30,130,29,130,28,130,27,130,26,164,31,8,31,184,31,184,30,217,31,10,31,222,31,222,30,195,31,157,31,217,31,61,31,231,31,44,31,124,31,20,31,20,30,222,31,65,31,251,31,193,31,216,31,54,31,224,31,46,31,46,30,137,31,198,31,250,31,127,31,46,31,170,31,203,31,203,30,19,31,69,31,175,31,175,30,21,31,221,31,147,31,74,31,74,30,74,29,146,31,155,31,122,31,69,31,91,31,91,30,116,31,116,30,116,29,185,31,121,31,149,31,77,31,226,31,240,31,240,30,240,29,177,31,60,31,133,31,133,30,74,31,224,31,103,31,152,31,58,31,164,31,164,30,225,31,63,31,101,31,145,31,7,31,7,30,24,31,24,30,253,31,175,31,105,31,105,30,41,31,61,31,148,31,92,31,22,31,174,31,229,31,179,31,187,31,66,31,67,31,102,31,122,31,122,30,182,31,189,31,214,31,222,31,157,31,12,31,217,31,217,30,217,29,25,31,50,31,254,31,61,31,34,31,222,31,181,31,15,31,93,31,143,31,22,31,22,30,28,31,68,31,133,31,133,30,184,31,11,31,171,31,225,31,225,30,55,31,20,31,133,31,199,31,184,31,184,30,181,31,78,31,49,31,62,31,84,31,84,30,84,29,51,31,252,31,124,31,39,31,39,30,245,31,208,31,243,31,152,31,65,31,91,31,86,31,55,31,43,31,8,31,14,31,151,31,101,31,197,31,197,30,154,31,154,30,95,31,95,30,254,31,253,31,253,30,211,31,211,30,21,31,180,31,147,31,147,30,37,31,114,31,100,31,243,31,252,31,39,31,47,31,4,31,66,31,229,31,85,31,211,31,225,31,64,31,234,31,151,31,76,31,76,30,249,31,125,31,190,31,112,31,112,30,112,29,100,31,145,31,242,31,242,30,195,31,62,31,55,31,80,31,80,31,148,31,148,30,171,31,171,30,218,31,218,30,218,29,121,31,233,31,233,30,18,31,100,31,56,31,13,31,75,31,236,31,14,31,157,31,119,31,213,31,213,30,102,31,161,31,115,31,66,31,133,31,133,30,179,31,196,31,16,31,61,31,61,30,77,31,38,31,172,31,172,30,108,31,108,30,221,31,190,31,148,31,26,31,33,31,125,31,19,31,59,31,131,31,234,31,112,31,84,31,84,30,90,31,44,31,44,30,243,31,85,31,73,31,159,31,84,31,253,31,221,31,213,31,106,31,211,31,184,31,118,31,50,31,222,31,2,31,95,31,23,31,65,31,143,31,143,30,85,31,85,30,85,29,233,31,231,31,53,31,68,31,39,31,213,31,107,31,127,31,126,31,164,31,241,31,78,31,58,31,58,30,58,29,164,31,254,31,118,31,19,31,249,31,79,31,117,31,52,31,133,31,198,31,198,30,198,29,20,31,34,31,217,31,110,31,13,31,13,30,181,31,242,31,83,31,83,30,120,31,58,31,131,31,243,31,151,31,151,30,10,31,51,31,51,30,51,29,51,28,18,31,241,31,107,31,103,31,64,31,167,31,174,31,224,31,224,30,224,29,214,31,78,31,78,30,186,31,155,31,79,31,88,31,88,30,5,31,5,30,133,31,133,30,133,29,10,31,13,31,197,31,244,31,187,31,23,31,23,30,23,29,253,31,123,31,231,31,41,31,224,31,224,30,182,31,182,30,100,31,156,31,34,31,37,31,37,30,37,29,17,31,182,31,182,30,99,31,5,31,173,31,241,31,164,31,224,31,90,31,1,31,123,31,152,31,121,31,91,31,166,31,166,30,17,31,17,30,255,31,255,30,75,31,77,31,99,31,30,31,228,31,239,31,213,31,35,31,139,31,55,31,222,31,208,31,135,31,9,31,95,31,121,31,145,31,226,31,100,31,83,31,202,31,37,31,224,31,67,31,41,31,177,31,139,31,181,31,59,31,21,31,212,31,175,31,245,31,245,30,118,31,118,30,108,31,220,31,240,31,240,30,240,31,55,31,140,31,170,31,170,30,140,31,33,31,152,31,152,30,233,31,124,31,158,31,68,31,241,31,207,31,112,31,42,31,1,31,1,30,55,31,152,31,46,31,139,31,139,30,187,31,17,31,178,31,181,31,94,31,141,31,149,31,149,30,4,31,4,30,47,31,47,30,47,29,117,31,62,31,62,30,81,31,219,31,125,31,176,31,118,31,118,30,3,31,116,31,48,31,22,31,51,31,105,31,73,31,98,31,215,31,109,31,173,31,76,31,114,31,188,31,75,31,75,30,26,31,155,31,242,31,144,31,144,30,216,31,8,31,165,31,42,31,157,31,84,31,159,31,66,31,80,31,63,31,7,31,234,31,94,31,217,31,217,30,217,29,131,31,223,31,175,31,240,31,181,31,181,30,209,31,224,31,41,31,41,30,240,31,132,31,182,31,145,31,140,31,140,30,110,31,76,31,25,31,25,30,45,31,184,31,60,31,59,31,124,31,37,31,226,31,240,31,147,31,87,31,135,31,202,31,171,31,158,31,96,31,19,31,238,31,63,31,63,30,63,29,18,31,107,31,192,31,148,31,148,30,194,31,201,31,201,30,149,31,211,31,211,30,222,31,47,31,84,31,195,31,18,31,18,30,18,29,18,28,92,31,92,30,87,31,148,31,124,31,124,30,125,31,170,31,248,31,209,31,98,31,239,31,203,31,118,31,243,31,243,30,235,31,149,31,223,31,243,31,101,31,126,31,203,31,175,31,55,31,55,30,55,29,59,31,59,30,59,29,149,31,141,31,20,31,49,31,218,31,248,31,82,31,143,31,85,31,36,31,36,30,159,31,7,31,208,31,27,31,65,31,81,31,195,31,248,31,77,31,77,30,54,31,231,31,74,31,96,31,93,31,93,30,67,31,67,30,138,31,34,31,185,31,185,30,211,31,51,31,126,31,203,31,203,30,108,31,173,31,213,31,222,31,161,31,161,30,164,31,164,30,149,31,149,30,149,29,245,31,46,31,42,31,42,30,32,31,172,31,132,31,164,31,159,31,52,31,52,30,169,31,35,31,109,31,152,31,152,30,207,31,84,31,65,31,79,31,185,31,151,31,157,31,157,30,144,31,47,31,142,31,142,30,1,31,141,31,141,30,236,31,41,31,41,30,29,31,29,30,15,31,53,31,175,31,108,31,75,31,75,30,4,31,4,30,223,31,39,31,137,31,42,31,252,31,252,30,252,29,205,31,76,31,239,31,18,31,238,31,176,31,176,30,66,31,119,31,194,31,182,31,102,31,159,31,159,30,65,31,65,30,169,31,130,31,134,31,10,31,212,31,5,31,72,31,180,31,177,31,106,31,42,31,42,30,174,31,236,31,56,31,58,31,243,31,216,31,216,30,211,31,62,31,32,31,32,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
