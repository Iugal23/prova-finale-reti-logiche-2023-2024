-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 949;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (162,0,178,0,0,0,0,0,44,0,84,0,6,0,22,0,200,0,226,0,24,0,179,0,23,0,28,0,0,0,99,0,154,0,0,0,139,0,110,0,59,0,165,0,40,0,87,0,0,0,36,0,61,0,91,0,73,0,124,0,7,0,0,0,26,0,59,0,129,0,226,0,69,0,0,0,80,0,1,0,0,0,209,0,160,0,83,0,0,0,152,0,137,0,236,0,0,0,29,0,203,0,184,0,243,0,0,0,208,0,220,0,164,0,19,0,0,0,147,0,173,0,2,0,189,0,0,0,0,0,114,0,0,0,236,0,182,0,39,0,67,0,129,0,0,0,0,0,221,0,0,0,0,0,62,0,94,0,195,0,203,0,23,0,179,0,220,0,0,0,217,0,125,0,89,0,163,0,117,0,155,0,163,0,235,0,55,0,67,0,189,0,16,0,104,0,41,0,99,0,54,0,158,0,154,0,133,0,69,0,12,0,80,0,222,0,0,0,87,0,47,0,24,0,70,0,197,0,190,0,192,0,192,0,0,0,73,0,0,0,98,0,107,0,134,0,134,0,16,0,0,0,7,0,44,0,154,0,11,0,176,0,219,0,71,0,224,0,253,0,0,0,0,0,192,0,0,0,0,0,140,0,156,0,215,0,31,0,44,0,195,0,68,0,30,0,144,0,157,0,36,0,45,0,184,0,29,0,128,0,0,0,46,0,85,0,0,0,71,0,120,0,168,0,0,0,179,0,43,0,177,0,0,0,147,0,0,0,0,0,0,0,165,0,251,0,32,0,36,0,249,0,22,0,198,0,0,0,0,0,21,0,31,0,9,0,0,0,0,0,124,0,176,0,175,0,154,0,247,0,163,0,243,0,57,0,86,0,216,0,221,0,250,0,132,0,135,0,169,0,0,0,146,0,162,0,0,0,72,0,69,0,116,0,8,0,169,0,186,0,206,0,0,0,0,0,177,0,8,0,79,0,115,0,89,0,179,0,123,0,255,0,34,0,0,0,71,0,59,0,0,0,31,0,55,0,242,0,25,0,0,0,93,0,0,0,188,0,18,0,0,0,187,0,0,0,34,0,158,0,111,0,0,0,140,0,0,0,0,0,0,0,99,0,0,0,230,0,235,0,114,0,117,0,69,0,136,0,63,0,11,0,154,0,9,0,0,0,26,0,54,0,124,0,139,0,68,0,172,0,195,0,0,0,14,0,116,0,96,0,0,0,176,0,0,0,210,0,206,0,223,0,46,0,191,0,0,0,89,0,196,0,104,0,0,0,0,0,0,0,34,0,200,0,94,0,0,0,160,0,0,0,96,0,0,0,0,0,149,0,21,0,90,0,128,0,0,0,0,0,0,0,0,0,80,0,187,0,0,0,36,0,0,0,109,0,108,0,121,0,190,0,125,0,27,0,102,0,19,0,194,0,3,0,4,0,254,0,111,0,122,0,62,0,132,0,90,0,201,0,217,0,102,0,231,0,245,0,137,0,27,0,44,0,191,0,69,0,57,0,0,0,9,0,93,0,193,0,233,0,175,0,0,0,41,0,158,0,169,0,88,0,191,0,229,0,32,0,179,0,92,0,205,0,123,0,0,0,211,0,215,0,150,0,0,0,48,0,235,0,32,0,207,0,0,0,21,0,243,0,36,0,229,0,175,0,181,0,108,0,238,0,183,0,32,0,247,0,174,0,93,0,0,0,219,0,41,0,110,0,212,0,0,0,14,0,189,0,198,0,25,0,35,0,0,0,72,0,0,0,254,0,3,0,190,0,155,0,12,0,33,0,52,0,121,0,117,0,170,0,0,0,53,0,121,0,0,0,133,0,229,0,110,0,240,0,112,0,248,0,0,0,41,0,64,0,28,0,243,0,0,0,0,0,142,0,92,0,79,0,209,0,137,0,240,0,0,0,0,0,0,0,0,0,0,0,23,0,25,0,33,0,63,0,241,0,176,0,123,0,238,0,65,0,110,0,138,0,0,0,0,0,1,0,201,0,73,0,88,0,0,0,0,0,65,0,134,0,143,0,52,0,20,0,61,0,61,0,103,0,36,0,99,0,0,0,214,0,232,0,139,0,142,0,0,0,75,0,12,0,183,0,0,0,73,0,240,0,175,0,0,0,87,0,58,0,198,0,56,0,151,0,250,0,235,0,118,0,0,0,100,0,149,0,225,0,251,0,38,0,0,0,0,0,0,0,4,0,163,0,68,0,119,0,78,0,118,0,0,0,232,0,0,0,139,0,76,0,52,0,11,0,135,0,180,0,0,0,232,0,157,0,239,0,0,0,79,0,205,0,0,0,89,0,197,0,99,0,247,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,70,0,119,0,163,0,247,0,249,0,0,0,112,0,251,0,125,0,63,0,20,0,22,0,0,0,0,0,0,0,49,0,194,0,227,0,0,0,146,0,100,0,0,0,0,0,214,0,161,0,0,0,243,0,76,0,173,0,160,0,191,0,17,0,142,0,250,0,228,0,100,0,65,0,137,0,0,0,51,0,48,0,31,0,0,0,58,0,65,0,180,0,210,0,0,0,0,0,44,0,123,0,206,0,242,0,86,0,0,0,196,0,157,0,0,0,0,0,243,0,118,0,95,0,0,0,0,0,114,0,0,0,0,0,182,0,96,0,130,0,0,0,71,0,154,0,21,0,0,0,0,0,25,0,100,0,244,0,8,0,198,0,0,0,93,0,16,0,178,0,102,0,159,0,6,0,5,0,0,0,0,0,252,0,0,0,171,0,148,0,252,0,0,0,236,0,181,0,160,0,189,0,81,0,167,0,107,0,33,0,0,0,242,0,0,0,0,0,210,0,0,0,101,0,0,0,5,0,0,0,0,0,211,0,132,0,0,0,172,0,0,0,145,0,76,0,54,0,0,0,43,0,160,0,0,0,248,0,50,0,156,0,178,0,177,0,0,0,6,0,0,0,228,0,117,0,162,0,192,0,89,0,234,0,0,0,22,0,213,0,119,0,52,0,90,0,150,0,153,0,211,0,155,0,131,0,81,0,112,0,251,0,207,0,67,0,178,0,150,0,0,0,92,0,61,0,0,0,0,0,197,0,0,0,28,0,0,0,72,0,0,0,198,0,213,0,0,0,140,0,35,0,4,0,90,0,109,0,15,0,94,0,232,0,233,0,42,0,0,0,19,0,0,0,36,0,172,0,8,0,31,0,100,0,139,0,172,0,33,0,0,0,0,0,130,0,190,0,39,0,169,0,67,0,0,0,84,0,52,0,221,0,125,0,22,0,93,0,14,0,245,0,37,0,2,0,62,0,161,0,86,0,54,0,142,0,79,0,188,0,223,0,89,0,184,0,144,0,199,0,51,0,0,0,85,0,35,0,251,0,161,0,198,0,98,0,179,0,106,0,147,0,106,0,251,0,69,0,2,0,173,0,193,0,71,0,187,0,201,0,229,0,115,0,212,0,247,0,70,0,167,0,96,0,152,0,199,0,41,0,13,0,114,0,157,0,0,0,0,0,199,0,231,0,253,0,41,0,168,0,181,0,188,0,0,0,38,0,211,0,0,0,119,0,152,0,180,0,0,0,0,0,13,0,20,0,97,0,246,0,102,0,72,0,104,0,172,0,220,0,19,0,206,0,0,0,89,0,22,0,0,0,233,0,171,0,0,0,22,0,92,0,252,0,131,0,217,0,39,0,189,0,64,0,112,0,126,0,0,0,44,0,45,0,0,0,91,0,0,0,29,0,137,0,249,0,241,0,219,0,118,0,231,0,244,0,166,0,138,0,191,0,100,0,66,0,96,0,11,0,210,0,246,0,5,0,211,0,0,0,199,0,209,0,111,0,177,0,0,0,161,0,198,0,0,0,93,0,184,0,162,0,176,0,96,0,196,0,188,0,201,0,67,0,238,0,0,0,157,0,222,0,102,0,12,0,0,0,221,0,0,0,32,0,192,0,250,0,178,0,212,0,55,0,242,0,176,0,0,0,119,0,0,0,23,0,44,0,0,0,76,0,203,0,100,0,72,0,99,0,163,0,0,0,79,0,161,0,197,0,109,0,193,0,0,0,84,0,7,0,223,0,0,0,0,0,0,0,101,0,250,0,164,0,125,0,40,0,95,0,197,0,32,0,0,0,82,0,227,0,185,0,232,0,120,0,0,0,230,0,0,0,27,0,0,0,160,0,3,0,171,0,128,0,0,0,103,0,115,0,49,0,73,0,0,0,55,0,115,0,51,0,75,0,143,0,0,0,123,0,144,0,147,0);
signal scenario_full  : scenario_type := (162,31,178,31,178,30,178,29,44,31,84,31,6,31,22,31,200,31,226,31,24,31,179,31,23,31,28,31,28,30,99,31,154,31,154,30,139,31,110,31,59,31,165,31,40,31,87,31,87,30,36,31,61,31,91,31,73,31,124,31,7,31,7,30,26,31,59,31,129,31,226,31,69,31,69,30,80,31,1,31,1,30,209,31,160,31,83,31,83,30,152,31,137,31,236,31,236,30,29,31,203,31,184,31,243,31,243,30,208,31,220,31,164,31,19,31,19,30,147,31,173,31,2,31,189,31,189,30,189,29,114,31,114,30,236,31,182,31,39,31,67,31,129,31,129,30,129,29,221,31,221,30,221,29,62,31,94,31,195,31,203,31,23,31,179,31,220,31,220,30,217,31,125,31,89,31,163,31,117,31,155,31,163,31,235,31,55,31,67,31,189,31,16,31,104,31,41,31,99,31,54,31,158,31,154,31,133,31,69,31,12,31,80,31,222,31,222,30,87,31,47,31,24,31,70,31,197,31,190,31,192,31,192,31,192,30,73,31,73,30,98,31,107,31,134,31,134,31,16,31,16,30,7,31,44,31,154,31,11,31,176,31,219,31,71,31,224,31,253,31,253,30,253,29,192,31,192,30,192,29,140,31,156,31,215,31,31,31,44,31,195,31,68,31,30,31,144,31,157,31,36,31,45,31,184,31,29,31,128,31,128,30,46,31,85,31,85,30,71,31,120,31,168,31,168,30,179,31,43,31,177,31,177,30,147,31,147,30,147,29,147,28,165,31,251,31,32,31,36,31,249,31,22,31,198,31,198,30,198,29,21,31,31,31,9,31,9,30,9,29,124,31,176,31,175,31,154,31,247,31,163,31,243,31,57,31,86,31,216,31,221,31,250,31,132,31,135,31,169,31,169,30,146,31,162,31,162,30,72,31,69,31,116,31,8,31,169,31,186,31,206,31,206,30,206,29,177,31,8,31,79,31,115,31,89,31,179,31,123,31,255,31,34,31,34,30,71,31,59,31,59,30,31,31,55,31,242,31,25,31,25,30,93,31,93,30,188,31,18,31,18,30,187,31,187,30,34,31,158,31,111,31,111,30,140,31,140,30,140,29,140,28,99,31,99,30,230,31,235,31,114,31,117,31,69,31,136,31,63,31,11,31,154,31,9,31,9,30,26,31,54,31,124,31,139,31,68,31,172,31,195,31,195,30,14,31,116,31,96,31,96,30,176,31,176,30,210,31,206,31,223,31,46,31,191,31,191,30,89,31,196,31,104,31,104,30,104,29,104,28,34,31,200,31,94,31,94,30,160,31,160,30,96,31,96,30,96,29,149,31,21,31,90,31,128,31,128,30,128,29,128,28,128,27,80,31,187,31,187,30,36,31,36,30,109,31,108,31,121,31,190,31,125,31,27,31,102,31,19,31,194,31,3,31,4,31,254,31,111,31,122,31,62,31,132,31,90,31,201,31,217,31,102,31,231,31,245,31,137,31,27,31,44,31,191,31,69,31,57,31,57,30,9,31,93,31,193,31,233,31,175,31,175,30,41,31,158,31,169,31,88,31,191,31,229,31,32,31,179,31,92,31,205,31,123,31,123,30,211,31,215,31,150,31,150,30,48,31,235,31,32,31,207,31,207,30,21,31,243,31,36,31,229,31,175,31,181,31,108,31,238,31,183,31,32,31,247,31,174,31,93,31,93,30,219,31,41,31,110,31,212,31,212,30,14,31,189,31,198,31,25,31,35,31,35,30,72,31,72,30,254,31,3,31,190,31,155,31,12,31,33,31,52,31,121,31,117,31,170,31,170,30,53,31,121,31,121,30,133,31,229,31,110,31,240,31,112,31,248,31,248,30,41,31,64,31,28,31,243,31,243,30,243,29,142,31,92,31,79,31,209,31,137,31,240,31,240,30,240,29,240,28,240,27,240,26,23,31,25,31,33,31,63,31,241,31,176,31,123,31,238,31,65,31,110,31,138,31,138,30,138,29,1,31,201,31,73,31,88,31,88,30,88,29,65,31,134,31,143,31,52,31,20,31,61,31,61,31,103,31,36,31,99,31,99,30,214,31,232,31,139,31,142,31,142,30,75,31,12,31,183,31,183,30,73,31,240,31,175,31,175,30,87,31,58,31,198,31,56,31,151,31,250,31,235,31,118,31,118,30,100,31,149,31,225,31,251,31,38,31,38,30,38,29,38,28,4,31,163,31,68,31,119,31,78,31,118,31,118,30,232,31,232,30,139,31,76,31,52,31,11,31,135,31,180,31,180,30,232,31,157,31,239,31,239,30,79,31,205,31,205,30,89,31,197,31,99,31,247,31,247,30,247,29,247,28,247,27,247,26,247,25,247,24,70,31,119,31,163,31,247,31,249,31,249,30,112,31,251,31,125,31,63,31,20,31,22,31,22,30,22,29,22,28,49,31,194,31,227,31,227,30,146,31,100,31,100,30,100,29,214,31,161,31,161,30,243,31,76,31,173,31,160,31,191,31,17,31,142,31,250,31,228,31,100,31,65,31,137,31,137,30,51,31,48,31,31,31,31,30,58,31,65,31,180,31,210,31,210,30,210,29,44,31,123,31,206,31,242,31,86,31,86,30,196,31,157,31,157,30,157,29,243,31,118,31,95,31,95,30,95,29,114,31,114,30,114,29,182,31,96,31,130,31,130,30,71,31,154,31,21,31,21,30,21,29,25,31,100,31,244,31,8,31,198,31,198,30,93,31,16,31,178,31,102,31,159,31,6,31,5,31,5,30,5,29,252,31,252,30,171,31,148,31,252,31,252,30,236,31,181,31,160,31,189,31,81,31,167,31,107,31,33,31,33,30,242,31,242,30,242,29,210,31,210,30,101,31,101,30,5,31,5,30,5,29,211,31,132,31,132,30,172,31,172,30,145,31,76,31,54,31,54,30,43,31,160,31,160,30,248,31,50,31,156,31,178,31,177,31,177,30,6,31,6,30,228,31,117,31,162,31,192,31,89,31,234,31,234,30,22,31,213,31,119,31,52,31,90,31,150,31,153,31,211,31,155,31,131,31,81,31,112,31,251,31,207,31,67,31,178,31,150,31,150,30,92,31,61,31,61,30,61,29,197,31,197,30,28,31,28,30,72,31,72,30,198,31,213,31,213,30,140,31,35,31,4,31,90,31,109,31,15,31,94,31,232,31,233,31,42,31,42,30,19,31,19,30,36,31,172,31,8,31,31,31,100,31,139,31,172,31,33,31,33,30,33,29,130,31,190,31,39,31,169,31,67,31,67,30,84,31,52,31,221,31,125,31,22,31,93,31,14,31,245,31,37,31,2,31,62,31,161,31,86,31,54,31,142,31,79,31,188,31,223,31,89,31,184,31,144,31,199,31,51,31,51,30,85,31,35,31,251,31,161,31,198,31,98,31,179,31,106,31,147,31,106,31,251,31,69,31,2,31,173,31,193,31,71,31,187,31,201,31,229,31,115,31,212,31,247,31,70,31,167,31,96,31,152,31,199,31,41,31,13,31,114,31,157,31,157,30,157,29,199,31,231,31,253,31,41,31,168,31,181,31,188,31,188,30,38,31,211,31,211,30,119,31,152,31,180,31,180,30,180,29,13,31,20,31,97,31,246,31,102,31,72,31,104,31,172,31,220,31,19,31,206,31,206,30,89,31,22,31,22,30,233,31,171,31,171,30,22,31,92,31,252,31,131,31,217,31,39,31,189,31,64,31,112,31,126,31,126,30,44,31,45,31,45,30,91,31,91,30,29,31,137,31,249,31,241,31,219,31,118,31,231,31,244,31,166,31,138,31,191,31,100,31,66,31,96,31,11,31,210,31,246,31,5,31,211,31,211,30,199,31,209,31,111,31,177,31,177,30,161,31,198,31,198,30,93,31,184,31,162,31,176,31,96,31,196,31,188,31,201,31,67,31,238,31,238,30,157,31,222,31,102,31,12,31,12,30,221,31,221,30,32,31,192,31,250,31,178,31,212,31,55,31,242,31,176,31,176,30,119,31,119,30,23,31,44,31,44,30,76,31,203,31,100,31,72,31,99,31,163,31,163,30,79,31,161,31,197,31,109,31,193,31,193,30,84,31,7,31,223,31,223,30,223,29,223,28,101,31,250,31,164,31,125,31,40,31,95,31,197,31,32,31,32,30,82,31,227,31,185,31,232,31,120,31,120,30,230,31,230,30,27,31,27,30,160,31,3,31,171,31,128,31,128,30,103,31,115,31,49,31,73,31,73,30,55,31,115,31,51,31,75,31,143,31,143,30,123,31,144,31,147,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
