-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 317;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (49,0,0,0,0,0,185,0,2,0,79,0,240,0,0,0,210,0,6,0,199,0,1,0,0,0,4,0,116,0,0,0,45,0,199,0,0,0,232,0,230,0,0,0,251,0,158,0,63,0,25,0,85,0,101,0,160,0,105,0,0,0,56,0,135,0,0,0,182,0,107,0,183,0,96,0,0,0,66,0,60,0,0,0,32,0,164,0,129,0,98,0,0,0,0,0,105,0,137,0,182,0,0,0,130,0,140,0,24,0,0,0,232,0,45,0,252,0,108,0,220,0,185,0,254,0,0,0,83,0,60,0,167,0,0,0,34,0,78,0,17,0,101,0,252,0,153,0,172,0,126,0,102,0,251,0,0,0,0,0,46,0,0,0,212,0,198,0,0,0,54,0,54,0,216,0,115,0,142,0,128,0,189,0,0,0,231,0,0,0,20,0,227,0,15,0,154,0,215,0,22,0,215,0,0,0,187,0,0,0,206,0,92,0,249,0,0,0,136,0,13,0,106,0,0,0,0,0,59,0,112,0,74,0,251,0,0,0,70,0,0,0,125,0,254,0,181,0,0,0,137,0,217,0,27,0,2,0,100,0,49,0,89,0,0,0,0,0,0,0,14,0,221,0,151,0,30,0,0,0,112,0,32,0,153,0,134,0,78,0,235,0,132,0,130,0,141,0,89,0,2,0,0,0,216,0,98,0,186,0,65,0,0,0,157,0,111,0,114,0,116,0,0,0,135,0,124,0,102,0,178,0,0,0,6,0,57,0,127,0,108,0,212,0,100,0,32,0,0,0,247,0,188,0,220,0,226,0,232,0,208,0,66,0,235,0,144,0,109,0,38,0,200,0,47,0,55,0,66,0,249,0,173,0,214,0,104,0,113,0,0,0,0,0,11,0,44,0,250,0,53,0,90,0,160,0,118,0,31,0,167,0,109,0,0,0,191,0,145,0,160,0,238,0,0,0,105,0,0,0,245,0,229,0,124,0,0,0,188,0,241,0,227,0,241,0,145,0,0,0,39,0,187,0,0,0,0,0,128,0,0,0,0,0,104,0,139,0,237,0,43,0,56,0,183,0,215,0,0,0,16,0,200,0,70,0,117,0,43,0,0,0,0,0,146,0,0,0,243,0,205,0,173,0,0,0,0,0,219,0,0,0,0,0,42,0,192,0,77,0,51,0,60,0,239,0,106,0,9,0,5,0,0,0,0,0,216,0,26,0,0,0,112,0,207,0,199,0,132,0,10,0,219,0,226,0,112,0,179,0,85,0,214,0,165,0,0,0,0,0,40,0,180,0,75,0,229,0,37,0,0,0,207,0,96,0,28,0,201,0,0,0,147,0,221,0,164,0,215,0,0,0,252,0,189,0,190,0,226,0,138,0,154,0,0,0,79,0,79,0,105,0,121,0,154,0,35,0,16,0,33,0,181,0);
signal scenario_full  : scenario_type := (49,31,49,30,49,29,185,31,2,31,79,31,240,31,240,30,210,31,6,31,199,31,1,31,1,30,4,31,116,31,116,30,45,31,199,31,199,30,232,31,230,31,230,30,251,31,158,31,63,31,25,31,85,31,101,31,160,31,105,31,105,30,56,31,135,31,135,30,182,31,107,31,183,31,96,31,96,30,66,31,60,31,60,30,32,31,164,31,129,31,98,31,98,30,98,29,105,31,137,31,182,31,182,30,130,31,140,31,24,31,24,30,232,31,45,31,252,31,108,31,220,31,185,31,254,31,254,30,83,31,60,31,167,31,167,30,34,31,78,31,17,31,101,31,252,31,153,31,172,31,126,31,102,31,251,31,251,30,251,29,46,31,46,30,212,31,198,31,198,30,54,31,54,31,216,31,115,31,142,31,128,31,189,31,189,30,231,31,231,30,20,31,227,31,15,31,154,31,215,31,22,31,215,31,215,30,187,31,187,30,206,31,92,31,249,31,249,30,136,31,13,31,106,31,106,30,106,29,59,31,112,31,74,31,251,31,251,30,70,31,70,30,125,31,254,31,181,31,181,30,137,31,217,31,27,31,2,31,100,31,49,31,89,31,89,30,89,29,89,28,14,31,221,31,151,31,30,31,30,30,112,31,32,31,153,31,134,31,78,31,235,31,132,31,130,31,141,31,89,31,2,31,2,30,216,31,98,31,186,31,65,31,65,30,157,31,111,31,114,31,116,31,116,30,135,31,124,31,102,31,178,31,178,30,6,31,57,31,127,31,108,31,212,31,100,31,32,31,32,30,247,31,188,31,220,31,226,31,232,31,208,31,66,31,235,31,144,31,109,31,38,31,200,31,47,31,55,31,66,31,249,31,173,31,214,31,104,31,113,31,113,30,113,29,11,31,44,31,250,31,53,31,90,31,160,31,118,31,31,31,167,31,109,31,109,30,191,31,145,31,160,31,238,31,238,30,105,31,105,30,245,31,229,31,124,31,124,30,188,31,241,31,227,31,241,31,145,31,145,30,39,31,187,31,187,30,187,29,128,31,128,30,128,29,104,31,139,31,237,31,43,31,56,31,183,31,215,31,215,30,16,31,200,31,70,31,117,31,43,31,43,30,43,29,146,31,146,30,243,31,205,31,173,31,173,30,173,29,219,31,219,30,219,29,42,31,192,31,77,31,51,31,60,31,239,31,106,31,9,31,5,31,5,30,5,29,216,31,26,31,26,30,112,31,207,31,199,31,132,31,10,31,219,31,226,31,112,31,179,31,85,31,214,31,165,31,165,30,165,29,40,31,180,31,75,31,229,31,37,31,37,30,207,31,96,31,28,31,201,31,201,30,147,31,221,31,164,31,215,31,215,30,252,31,189,31,190,31,226,31,138,31,154,31,154,30,79,31,79,31,105,31,121,31,154,31,35,31,16,31,33,31,181,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
