-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_123 is
end project_tb_123;

architecture project_tb_arch_123 of project_tb_123 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 946;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (71,0,0,0,79,0,151,0,125,0,28,0,29,0,160,0,129,0,73,0,31,0,243,0,0,0,205,0,3,0,125,0,0,0,117,0,219,0,0,0,247,0,49,0,48,0,8,0,0,0,0,0,28,0,0,0,8,0,240,0,18,0,0,0,126,0,0,0,173,0,71,0,249,0,117,0,102,0,212,0,35,0,0,0,52,0,61,0,201,0,10,0,55,0,176,0,218,0,63,0,243,0,117,0,170,0,0,0,26,0,83,0,197,0,36,0,229,0,0,0,0,0,0,0,198,0,226,0,197,0,143,0,145,0,93,0,66,0,0,0,92,0,21,0,73,0,192,0,61,0,178,0,125,0,0,0,22,0,0,0,163,0,22,0,24,0,0,0,171,0,0,0,124,0,180,0,203,0,0,0,0,0,59,0,0,0,216,0,0,0,91,0,178,0,135,0,180,0,0,0,166,0,196,0,239,0,251,0,238,0,225,0,162,0,152,0,0,0,211,0,94,0,249,0,69,0,101,0,72,0,118,0,0,0,0,0,0,0,139,0,0,0,28,0,177,0,0,0,90,0,90,0,0,0,73,0,170,0,0,0,103,0,16,0,102,0,132,0,0,0,0,0,249,0,171,0,212,0,69,0,78,0,17,0,0,0,122,0,27,0,54,0,106,0,76,0,153,0,166,0,129,0,223,0,153,0,248,0,28,0,110,0,214,0,214,0,47,0,20,0,162,0,136,0,202,0,74,0,105,0,0,0,61,0,130,0,96,0,0,0,25,0,192,0,120,0,0,0,52,0,0,0,15,0,249,0,47,0,238,0,86,0,99,0,207,0,0,0,80,0,0,0,42,0,224,0,99,0,66,0,109,0,0,0,180,0,0,0,0,0,50,0,28,0,159,0,72,0,53,0,0,0,90,0,224,0,0,0,152,0,0,0,0,0,102,0,105,0,103,0,86,0,232,0,78,0,127,0,148,0,21,0,209,0,101,0,237,0,203,0,140,0,221,0,194,0,128,0,182,0,157,0,254,0,0,0,0,0,0,0,86,0,235,0,183,0,58,0,80,0,253,0,62,0,86,0,0,0,157,0,17,0,97,0,203,0,62,0,0,0,118,0,149,0,64,0,156,0,83,0,250,0,135,0,48,0,0,0,0,0,0,0,0,0,179,0,244,0,143,0,0,0,13,0,143,0,145,0,65,0,143,0,250,0,240,0,231,0,171,0,0,0,84,0,173,0,0,0,236,0,117,0,33,0,135,0,190,0,43,0,96,0,141,0,15,0,170,0,99,0,0,0,0,0,125,0,84,0,235,0,77,0,72,0,159,0,74,0,176,0,88,0,150,0,134,0,231,0,92,0,27,0,228,0,0,0,140,0,190,0,135,0,54,0,152,0,186,0,191,0,0,0,110,0,0,0,34,0,0,0,0,0,60,0,44,0,56,0,12,0,249,0,55,0,71,0,209,0,69,0,14,0,105,0,101,0,4,0,0,0,93,0,38,0,247,0,210,0,172,0,224,0,12,0,143,0,254,0,98,0,214,0,52,0,0,0,76,0,67,0,74,0,21,0,254,0,198,0,232,0,59,0,67,0,0,0,0,0,248,0,0,0,17,0,0,0,0,0,66,0,71,0,37,0,39,0,0,0,108,0,0,0,47,0,45,0,0,0,212,0,0,0,0,0,200,0,133,0,135,0,66,0,196,0,63,0,0,0,178,0,0,0,158,0,0,0,249,0,45,0,34,0,158,0,0,0,134,0,130,0,204,0,102,0,96,0,0,0,70,0,33,0,0,0,33,0,0,0,34,0,230,0,0,0,50,0,57,0,166,0,0,0,248,0,200,0,142,0,101,0,219,0,111,0,63,0,39,0,108,0,172,0,70,0,31,0,0,0,82,0,132,0,230,0,34,0,163,0,39,0,214,0,166,0,24,0,63,0,0,0,0,0,164,0,236,0,174,0,69,0,171,0,0,0,0,0,99,0,0,0,0,0,186,0,75,0,187,0,52,0,41,0,138,0,179,0,83,0,241,0,218,0,0,0,220,0,15,0,118,0,0,0,0,0,11,0,172,0,89,0,144,0,35,0,233,0,13,0,66,0,185,0,156,0,23,0,200,0,197,0,149,0,0,0,116,0,203,0,134,0,130,0,173,0,139,0,218,0,193,0,110,0,91,0,64,0,233,0,161,0,115,0,244,0,132,0,0,0,242,0,200,0,232,0,106,0,35,0,0,0,140,0,158,0,27,0,0,0,123,0,215,0,0,0,210,0,144,0,0,0,155,0,1,0,42,0,118,0,209,0,155,0,0,0,201,0,94,0,0,0,19,0,27,0,115,0,244,0,255,0,73,0,182,0,20,0,69,0,106,0,36,0,252,0,203,0,137,0,225,0,144,0,68,0,178,0,0,0,250,0,15,0,0,0,1,0,181,0,118,0,0,0,231,0,137,0,243,0,174,0,180,0,3,0,0,0,239,0,131,0,58,0,24,0,182,0,7,0,84,0,6,0,178,0,109,0,163,0,0,0,131,0,183,0,0,0,174,0,119,0,17,0,50,0,46,0,212,0,24,0,98,0,176,0,203,0,0,0,54,0,58,0,49,0,109,0,15,0,14,0,0,0,21,0,159,0,181,0,51,0,164,0,218,0,101,0,105,0,0,0,188,0,80,0,221,0,97,0,0,0,45,0,0,0,200,0,107,0,57,0,52,0,0,0,0,0,0,0,248,0,92,0,92,0,119,0,71,0,96,0,0,0,232,0,0,0,122,0,143,0,231,0,0,0,0,0,172,0,115,0,201,0,218,0,42,0,195,0,68,0,0,0,166,0,225,0,67,0,112,0,246,0,46,0,196,0,191,0,0,0,0,0,126,0,163,0,194,0,130,0,235,0,227,0,157,0,91,0,10,0,100,0,202,0,137,0,204,0,213,0,214,0,0,0,149,0,0,0,167,0,83,0,0,0,211,0,150,0,255,0,0,0,11,0,15,0,204,0,2,0,0,0,197,0,136,0,15,0,154,0,57,0,221,0,90,0,94,0,1,0,108,0,217,0,127,0,139,0,177,0,149,0,97,0,19,0,0,0,0,0,54,0,117,0,0,0,222,0,218,0,146,0,160,0,199,0,0,0,0,0,241,0,196,0,101,0,139,0,181,0,227,0,209,0,31,0,0,0,18,0,46,0,94,0,150,0,18,0,89,0,224,0,108,0,94,0,109,0,107,0,179,0,175,0,0,0,2,0,176,0,21,0,153,0,193,0,20,0,137,0,125,0,100,0,212,0,26,0,0,0,213,0,200,0,189,0,0,0,12,0,135,0,28,0,0,0,129,0,178,0,96,0,25,0,146,0,108,0,11,0,0,0,58,0,154,0,151,0,2,0,107,0,210,0,86,0,0,0,85,0,17,0,29,0,30,0,42,0,175,0,109,0,128,0,26,0,192,0,106,0,238,0,223,0,65,0,0,0,35,0,168,0,211,0,65,0,195,0,59,0,197,0,175,0,61,0,66,0,88,0,69,0,84,0,210,0,193,0,0,0,0,0,0,0,241,0,21,0,0,0,143,0,110,0,94,0,0,0,0,0,125,0,8,0,37,0,239,0,200,0,137,0,0,0,122,0,247,0,5,0,0,0,124,0,0,0,3,0,192,0,58,0,229,0,60,0,0,0,47,0,167,0,109,0,184,0,98,0,47,0,42,0,0,0,0,0,183,0,100,0,150,0,0,0,120,0,253,0,40,0,108,0,177,0,243,0,0,0,239,0,217,0,52,0,134,0,216,0,135,0,249,0,69,0,77,0,186,0,154,0,66,0,198,0,160,0,0,0,0,0,214,0,0,0,96,0,175,0,2,0,182,0,181,0,227,0,0,0,0,0,104,0,0,0,16,0,26,0,47,0,36,0,0,0,251,0,0,0,0,0,215,0,130,0,115,0,213,0,59,0,223,0,33,0,44,0,194,0,0,0,221,0,104,0,194,0,0,0,0,0,0,0,0,0,40,0,229,0,0,0,133,0,183,0,40,0,39,0,0,0,197,0,119,0,216,0,48,0,78,0,159,0,53,0,120,0,182,0,71,0,60,0,69,0,129,0,112,0,0,0,217,0,70,0,6,0,0,0,148,0,181,0,0,0,72,0,116,0,0,0,252,0,228,0,225,0,85,0,79,0,15,0,111,0,2,0,0,0,186,0,0,0,125,0,53,0,154,0,12,0,44,0,0,0,206,0,0,0,67,0,30,0,76,0,190,0,164,0,0,0,181,0);
signal scenario_full  : scenario_type := (71,31,71,30,79,31,151,31,125,31,28,31,29,31,160,31,129,31,73,31,31,31,243,31,243,30,205,31,3,31,125,31,125,30,117,31,219,31,219,30,247,31,49,31,48,31,8,31,8,30,8,29,28,31,28,30,8,31,240,31,18,31,18,30,126,31,126,30,173,31,71,31,249,31,117,31,102,31,212,31,35,31,35,30,52,31,61,31,201,31,10,31,55,31,176,31,218,31,63,31,243,31,117,31,170,31,170,30,26,31,83,31,197,31,36,31,229,31,229,30,229,29,229,28,198,31,226,31,197,31,143,31,145,31,93,31,66,31,66,30,92,31,21,31,73,31,192,31,61,31,178,31,125,31,125,30,22,31,22,30,163,31,22,31,24,31,24,30,171,31,171,30,124,31,180,31,203,31,203,30,203,29,59,31,59,30,216,31,216,30,91,31,178,31,135,31,180,31,180,30,166,31,196,31,239,31,251,31,238,31,225,31,162,31,152,31,152,30,211,31,94,31,249,31,69,31,101,31,72,31,118,31,118,30,118,29,118,28,139,31,139,30,28,31,177,31,177,30,90,31,90,31,90,30,73,31,170,31,170,30,103,31,16,31,102,31,132,31,132,30,132,29,249,31,171,31,212,31,69,31,78,31,17,31,17,30,122,31,27,31,54,31,106,31,76,31,153,31,166,31,129,31,223,31,153,31,248,31,28,31,110,31,214,31,214,31,47,31,20,31,162,31,136,31,202,31,74,31,105,31,105,30,61,31,130,31,96,31,96,30,25,31,192,31,120,31,120,30,52,31,52,30,15,31,249,31,47,31,238,31,86,31,99,31,207,31,207,30,80,31,80,30,42,31,224,31,99,31,66,31,109,31,109,30,180,31,180,30,180,29,50,31,28,31,159,31,72,31,53,31,53,30,90,31,224,31,224,30,152,31,152,30,152,29,102,31,105,31,103,31,86,31,232,31,78,31,127,31,148,31,21,31,209,31,101,31,237,31,203,31,140,31,221,31,194,31,128,31,182,31,157,31,254,31,254,30,254,29,254,28,86,31,235,31,183,31,58,31,80,31,253,31,62,31,86,31,86,30,157,31,17,31,97,31,203,31,62,31,62,30,118,31,149,31,64,31,156,31,83,31,250,31,135,31,48,31,48,30,48,29,48,28,48,27,179,31,244,31,143,31,143,30,13,31,143,31,145,31,65,31,143,31,250,31,240,31,231,31,171,31,171,30,84,31,173,31,173,30,236,31,117,31,33,31,135,31,190,31,43,31,96,31,141,31,15,31,170,31,99,31,99,30,99,29,125,31,84,31,235,31,77,31,72,31,159,31,74,31,176,31,88,31,150,31,134,31,231,31,92,31,27,31,228,31,228,30,140,31,190,31,135,31,54,31,152,31,186,31,191,31,191,30,110,31,110,30,34,31,34,30,34,29,60,31,44,31,56,31,12,31,249,31,55,31,71,31,209,31,69,31,14,31,105,31,101,31,4,31,4,30,93,31,38,31,247,31,210,31,172,31,224,31,12,31,143,31,254,31,98,31,214,31,52,31,52,30,76,31,67,31,74,31,21,31,254,31,198,31,232,31,59,31,67,31,67,30,67,29,248,31,248,30,17,31,17,30,17,29,66,31,71,31,37,31,39,31,39,30,108,31,108,30,47,31,45,31,45,30,212,31,212,30,212,29,200,31,133,31,135,31,66,31,196,31,63,31,63,30,178,31,178,30,158,31,158,30,249,31,45,31,34,31,158,31,158,30,134,31,130,31,204,31,102,31,96,31,96,30,70,31,33,31,33,30,33,31,33,30,34,31,230,31,230,30,50,31,57,31,166,31,166,30,248,31,200,31,142,31,101,31,219,31,111,31,63,31,39,31,108,31,172,31,70,31,31,31,31,30,82,31,132,31,230,31,34,31,163,31,39,31,214,31,166,31,24,31,63,31,63,30,63,29,164,31,236,31,174,31,69,31,171,31,171,30,171,29,99,31,99,30,99,29,186,31,75,31,187,31,52,31,41,31,138,31,179,31,83,31,241,31,218,31,218,30,220,31,15,31,118,31,118,30,118,29,11,31,172,31,89,31,144,31,35,31,233,31,13,31,66,31,185,31,156,31,23,31,200,31,197,31,149,31,149,30,116,31,203,31,134,31,130,31,173,31,139,31,218,31,193,31,110,31,91,31,64,31,233,31,161,31,115,31,244,31,132,31,132,30,242,31,200,31,232,31,106,31,35,31,35,30,140,31,158,31,27,31,27,30,123,31,215,31,215,30,210,31,144,31,144,30,155,31,1,31,42,31,118,31,209,31,155,31,155,30,201,31,94,31,94,30,19,31,27,31,115,31,244,31,255,31,73,31,182,31,20,31,69,31,106,31,36,31,252,31,203,31,137,31,225,31,144,31,68,31,178,31,178,30,250,31,15,31,15,30,1,31,181,31,118,31,118,30,231,31,137,31,243,31,174,31,180,31,3,31,3,30,239,31,131,31,58,31,24,31,182,31,7,31,84,31,6,31,178,31,109,31,163,31,163,30,131,31,183,31,183,30,174,31,119,31,17,31,50,31,46,31,212,31,24,31,98,31,176,31,203,31,203,30,54,31,58,31,49,31,109,31,15,31,14,31,14,30,21,31,159,31,181,31,51,31,164,31,218,31,101,31,105,31,105,30,188,31,80,31,221,31,97,31,97,30,45,31,45,30,200,31,107,31,57,31,52,31,52,30,52,29,52,28,248,31,92,31,92,31,119,31,71,31,96,31,96,30,232,31,232,30,122,31,143,31,231,31,231,30,231,29,172,31,115,31,201,31,218,31,42,31,195,31,68,31,68,30,166,31,225,31,67,31,112,31,246,31,46,31,196,31,191,31,191,30,191,29,126,31,163,31,194,31,130,31,235,31,227,31,157,31,91,31,10,31,100,31,202,31,137,31,204,31,213,31,214,31,214,30,149,31,149,30,167,31,83,31,83,30,211,31,150,31,255,31,255,30,11,31,15,31,204,31,2,31,2,30,197,31,136,31,15,31,154,31,57,31,221,31,90,31,94,31,1,31,108,31,217,31,127,31,139,31,177,31,149,31,97,31,19,31,19,30,19,29,54,31,117,31,117,30,222,31,218,31,146,31,160,31,199,31,199,30,199,29,241,31,196,31,101,31,139,31,181,31,227,31,209,31,31,31,31,30,18,31,46,31,94,31,150,31,18,31,89,31,224,31,108,31,94,31,109,31,107,31,179,31,175,31,175,30,2,31,176,31,21,31,153,31,193,31,20,31,137,31,125,31,100,31,212,31,26,31,26,30,213,31,200,31,189,31,189,30,12,31,135,31,28,31,28,30,129,31,178,31,96,31,25,31,146,31,108,31,11,31,11,30,58,31,154,31,151,31,2,31,107,31,210,31,86,31,86,30,85,31,17,31,29,31,30,31,42,31,175,31,109,31,128,31,26,31,192,31,106,31,238,31,223,31,65,31,65,30,35,31,168,31,211,31,65,31,195,31,59,31,197,31,175,31,61,31,66,31,88,31,69,31,84,31,210,31,193,31,193,30,193,29,193,28,241,31,21,31,21,30,143,31,110,31,94,31,94,30,94,29,125,31,8,31,37,31,239,31,200,31,137,31,137,30,122,31,247,31,5,31,5,30,124,31,124,30,3,31,192,31,58,31,229,31,60,31,60,30,47,31,167,31,109,31,184,31,98,31,47,31,42,31,42,30,42,29,183,31,100,31,150,31,150,30,120,31,253,31,40,31,108,31,177,31,243,31,243,30,239,31,217,31,52,31,134,31,216,31,135,31,249,31,69,31,77,31,186,31,154,31,66,31,198,31,160,31,160,30,160,29,214,31,214,30,96,31,175,31,2,31,182,31,181,31,227,31,227,30,227,29,104,31,104,30,16,31,26,31,47,31,36,31,36,30,251,31,251,30,251,29,215,31,130,31,115,31,213,31,59,31,223,31,33,31,44,31,194,31,194,30,221,31,104,31,194,31,194,30,194,29,194,28,194,27,40,31,229,31,229,30,133,31,183,31,40,31,39,31,39,30,197,31,119,31,216,31,48,31,78,31,159,31,53,31,120,31,182,31,71,31,60,31,69,31,129,31,112,31,112,30,217,31,70,31,6,31,6,30,148,31,181,31,181,30,72,31,116,31,116,30,252,31,228,31,225,31,85,31,79,31,15,31,111,31,2,31,2,30,186,31,186,30,125,31,53,31,154,31,12,31,44,31,44,30,206,31,206,30,67,31,30,31,76,31,190,31,164,31,164,30,181,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
