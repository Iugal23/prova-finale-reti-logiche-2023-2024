-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1003;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (56,0,0,0,151,0,174,0,218,0,75,0,152,0,114,0,158,0,215,0,204,0,0,0,0,0,113,0,12,0,87,0,72,0,46,0,91,0,53,0,0,0,0,0,48,0,31,0,14,0,0,0,249,0,144,0,137,0,113,0,69,0,175,0,0,0,226,0,37,0,245,0,0,0,73,0,106,0,4,0,10,0,0,0,0,0,181,0,21,0,200,0,0,0,0,0,0,0,1,0,33,0,36,0,96,0,187,0,38,0,244,0,184,0,174,0,49,0,206,0,0,0,24,0,27,0,50,0,138,0,204,0,0,0,92,0,43,0,0,0,131,0,0,0,92,0,50,0,49,0,104,0,61,0,135,0,140,0,159,0,0,0,183,0,99,0,0,0,201,0,181,0,130,0,0,0,0,0,0,0,242,0,88,0,0,0,59,0,224,0,226,0,224,0,242,0,174,0,6,0,0,0,45,0,183,0,0,0,180,0,97,0,108,0,52,0,115,0,33,0,241,0,0,0,193,0,144,0,12,0,0,0,191,0,27,0,78,0,48,0,93,0,60,0,235,0,48,0,0,0,0,0,5,0,224,0,120,0,237,0,136,0,0,0,0,0,28,0,190,0,230,0,236,0,230,0,83,0,68,0,0,0,215,0,0,0,247,0,99,0,149,0,208,0,0,0,22,0,226,0,0,0,175,0,0,0,128,0,0,0,96,0,195,0,0,0,19,0,121,0,84,0,79,0,63,0,35,0,192,0,111,0,225,0,128,0,0,0,0,0,240,0,79,0,194,0,103,0,76,0,48,0,114,0,13,0,8,0,202,0,248,0,190,0,154,0,150,0,29,0,74,0,59,0,96,0,81,0,171,0,0,0,155,0,8,0,46,0,39,0,113,0,31,0,1,0,0,0,239,0,54,0,65,0,225,0,114,0,105,0,0,0,0,0,103,0,11,0,117,0,201,0,0,0,111,0,53,0,57,0,141,0,31,0,178,0,0,0,16,0,0,0,206,0,53,0,216,0,96,0,0,0,1,0,0,0,0,0,253,0,0,0,66,0,173,0,20,0,114,0,0,0,0,0,15,0,0,0,219,0,211,0,163,0,173,0,217,0,223,0,105,0,0,0,163,0,64,0,0,0,77,0,203,0,33,0,72,0,0,0,178,0,0,0,67,0,186,0,88,0,154,0,149,0,0,0,0,0,0,0,0,0,0,0,245,0,97,0,0,0,0,0,0,0,156,0,106,0,29,0,72,0,0,0,215,0,144,0,57,0,213,0,183,0,0,0,153,0,121,0,29,0,0,0,131,0,149,0,123,0,100,0,0,0,0,0,66,0,122,0,150,0,10,0,83,0,65,0,80,0,238,0,161,0,207,0,0,0,0,0,2,0,0,0,127,0,177,0,0,0,163,0,0,0,198,0,176,0,135,0,85,0,66,0,81,0,174,0,213,0,0,0,0,0,29,0,92,0,179,0,30,0,91,0,191,0,151,0,0,0,82,0,230,0,53,0,4,0,15,0,207,0,142,0,114,0,160,0,49,0,144,0,3,0,0,0,102,0,132,0,216,0,55,0,0,0,0,0,52,0,12,0,0,0,44,0,16,0,160,0,39,0,227,0,155,0,66,0,195,0,51,0,14,0,180,0,103,0,122,0,0,0,0,0,179,0,78,0,85,0,130,0,125,0,132,0,0,0,186,0,100,0,0,0,242,0,243,0,168,0,107,0,78,0,18,0,0,0,26,0,99,0,230,0,71,0,227,0,123,0,70,0,20,0,216,0,156,0,106,0,161,0,95,0,0,0,30,0,180,0,168,0,209,0,19,0,207,0,0,0,134,0,88,0,122,0,5,0,0,0,123,0,121,0,28,0,212,0,134,0,0,0,18,0,0,0,64,0,0,0,131,0,49,0,69,0,154,0,38,0,156,0,0,0,153,0,236,0,159,0,128,0,23,0,133,0,0,0,49,0,92,0,186,0,59,0,147,0,80,0,181,0,0,0,12,0,112,0,180,0,179,0,107,0,0,0,112,0,3,0,119,0,43,0,192,0,96,0,83,0,185,0,88,0,24,0,164,0,59,0,112,0,79,0,16,0,101,0,174,0,177,0,27,0,178,0,123,0,161,0,68,0,119,0,0,0,0,0,107,0,252,0,30,0,0,0,0,0,201,0,156,0,79,0,23,0,0,0,219,0,0,0,206,0,0,0,0,0,127,0,116,0,45,0,0,0,90,0,71,0,199,0,12,0,142,0,106,0,197,0,51,0,30,0,201,0,38,0,186,0,86,0,0,0,100,0,0,0,7,0,226,0,49,0,132,0,216,0,8,0,49,0,0,0,95,0,148,0,40,0,153,0,177,0,231,0,0,0,163,0,3,0,230,0,5,0,95,0,107,0,0,0,9,0,13,0,230,0,0,0,239,0,187,0,88,0,0,0,159,0,199,0,61,0,0,0,27,0,89,0,171,0,42,0,0,0,0,0,89,0,85,0,195,0,212,0,13,0,147,0,116,0,0,0,0,0,141,0,253,0,0,0,158,0,58,0,149,0,166,0,0,0,0,0,13,0,0,0,22,0,220,0,0,0,31,0,102,0,133,0,22,0,105,0,76,0,143,0,124,0,0,0,34,0,12,0,76,0,21,0,222,0,129,0,250,0,34,0,139,0,74,0,9,0,141,0,4,0,93,0,15,0,178,0,252,0,64,0,29,0,17,0,252,0,209,0,8,0,0,0,237,0,68,0,191,0,201,0,106,0,139,0,35,0,167,0,169,0,42,0,240,0,224,0,14,0,0,0,186,0,48,0,113,0,243,0,32,0,227,0,0,0,125,0,46,0,0,0,0,0,231,0,27,0,223,0,68,0,0,0,247,0,17,0,0,0,225,0,68,0,174,0,230,0,87,0,130,0,205,0,209,0,157,0,226,0,0,0,85,0,15,0,0,0,101,0,213,0,41,0,0,0,45,0,239,0,144,0,54,0,30,0,172,0,225,0,75,0,11,0,245,0,223,0,62,0,37,0,0,0,209,0,31,0,208,0,207,0,146,0,35,0,41,0,182,0,131,0,118,0,151,0,98,0,96,0,178,0,128,0,51,0,163,0,29,0,0,0,98,0,149,0,113,0,0,0,222,0,0,0,15,0,57,0,0,0,56,0,95,0,182,0,0,0,0,0,96,0,159,0,252,0,57,0,128,0,23,0,94,0,135,0,210,0,10,0,178,0,228,0,236,0,0,0,18,0,0,0,220,0,245,0,146,0,228,0,63,0,0,0,128,0,255,0,117,0,149,0,192,0,0,0,93,0,164,0,216,0,40,0,217,0,153,0,0,0,0,0,131,0,0,0,92,0,126,0,44,0,144,0,0,0,101,0,185,0,15,0,125,0,0,0,126,0,0,0,0,0,66,0,243,0,73,0,0,0,107,0,0,0,0,0,77,0,213,0,238,0,208,0,0,0,20,0,159,0,137,0,32,0,93,0,0,0,247,0,137,0,232,0,0,0,54,0,243,0,168,0,121,0,113,0,82,0,135,0,21,0,105,0,105,0,22,0,90,0,0,0,224,0,234,0,196,0,40,0,69,0,0,0,105,0,0,0,30,0,198,0,213,0,41,0,0,0,206,0,0,0,110,0,79,0,0,0,139,0,63,0,202,0,244,0,229,0,8,0,184,0,27,0,25,0,152,0,120,0,255,0,26,0,218,0,141,0,241,0,49,0,173,0,247,0,16,0,49,0,169,0,142,0,209,0,161,0,70,0,192,0,197,0,85,0,49,0,46,0,0,0,70,0,88,0,243,0,50,0,253,0,221,0,0,0,31,0,0,0,11,0,0,0,72,0,165,0,1,0,48,0,0,0,195,0,29,0,10,0,129,0,177,0,225,0,94,0,39,0,188,0,239,0,124,0,45,0,134,0,28,0,27,0,48,0,91,0,128,0,0,0,213,0,0,0,25,0,59,0,1,0,128,0,218,0,28,0,41,0,0,0,136,0,227,0,0,0,238,0,50,0,139,0,0,0,128,0,82,0,85,0,56,0,61,0,56,0,142,0,0,0,193,0,180,0,114,0,0,0,0,0,120,0,130,0,72,0,15,0,49,0,199,0,184,0,54,0,142,0,67,0,41,0,211,0,117,0,133,0,148,0,66,0,53,0,124,0,24,0,2,0,129,0,130,0,0,0,82,0,63,0,162,0,0,0,27,0,0,0,0,0,245,0,225,0,78,0,0,0,124,0,40,0,13,0,204,0,156,0,230,0,5,0,147,0,55,0,204,0,188,0,209,0,86,0,77,0,53,0,199,0,30,0,0,0,184,0,49,0,39,0,210,0,52,0,235,0,22,0,84,0,20,0,25,0,1,0,1,0,33,0,34,0,3,0,203,0,0,0,0,0,180,0,190,0,252,0,228,0,0,0,58,0,144,0,182,0,0,0,238,0,0,0,92,0,244,0,205,0,245,0,161,0,45,0,147,0,118,0,250,0,239,0,0,0,149,0,0,0,164,0,225,0,51,0,101,0,106,0);
signal scenario_full  : scenario_type := (56,31,56,30,151,31,174,31,218,31,75,31,152,31,114,31,158,31,215,31,204,31,204,30,204,29,113,31,12,31,87,31,72,31,46,31,91,31,53,31,53,30,53,29,48,31,31,31,14,31,14,30,249,31,144,31,137,31,113,31,69,31,175,31,175,30,226,31,37,31,245,31,245,30,73,31,106,31,4,31,10,31,10,30,10,29,181,31,21,31,200,31,200,30,200,29,200,28,1,31,33,31,36,31,96,31,187,31,38,31,244,31,184,31,174,31,49,31,206,31,206,30,24,31,27,31,50,31,138,31,204,31,204,30,92,31,43,31,43,30,131,31,131,30,92,31,50,31,49,31,104,31,61,31,135,31,140,31,159,31,159,30,183,31,99,31,99,30,201,31,181,31,130,31,130,30,130,29,130,28,242,31,88,31,88,30,59,31,224,31,226,31,224,31,242,31,174,31,6,31,6,30,45,31,183,31,183,30,180,31,97,31,108,31,52,31,115,31,33,31,241,31,241,30,193,31,144,31,12,31,12,30,191,31,27,31,78,31,48,31,93,31,60,31,235,31,48,31,48,30,48,29,5,31,224,31,120,31,237,31,136,31,136,30,136,29,28,31,190,31,230,31,236,31,230,31,83,31,68,31,68,30,215,31,215,30,247,31,99,31,149,31,208,31,208,30,22,31,226,31,226,30,175,31,175,30,128,31,128,30,96,31,195,31,195,30,19,31,121,31,84,31,79,31,63,31,35,31,192,31,111,31,225,31,128,31,128,30,128,29,240,31,79,31,194,31,103,31,76,31,48,31,114,31,13,31,8,31,202,31,248,31,190,31,154,31,150,31,29,31,74,31,59,31,96,31,81,31,171,31,171,30,155,31,8,31,46,31,39,31,113,31,31,31,1,31,1,30,239,31,54,31,65,31,225,31,114,31,105,31,105,30,105,29,103,31,11,31,117,31,201,31,201,30,111,31,53,31,57,31,141,31,31,31,178,31,178,30,16,31,16,30,206,31,53,31,216,31,96,31,96,30,1,31,1,30,1,29,253,31,253,30,66,31,173,31,20,31,114,31,114,30,114,29,15,31,15,30,219,31,211,31,163,31,173,31,217,31,223,31,105,31,105,30,163,31,64,31,64,30,77,31,203,31,33,31,72,31,72,30,178,31,178,30,67,31,186,31,88,31,154,31,149,31,149,30,149,29,149,28,149,27,149,26,245,31,97,31,97,30,97,29,97,28,156,31,106,31,29,31,72,31,72,30,215,31,144,31,57,31,213,31,183,31,183,30,153,31,121,31,29,31,29,30,131,31,149,31,123,31,100,31,100,30,100,29,66,31,122,31,150,31,10,31,83,31,65,31,80,31,238,31,161,31,207,31,207,30,207,29,2,31,2,30,127,31,177,31,177,30,163,31,163,30,198,31,176,31,135,31,85,31,66,31,81,31,174,31,213,31,213,30,213,29,29,31,92,31,179,31,30,31,91,31,191,31,151,31,151,30,82,31,230,31,53,31,4,31,15,31,207,31,142,31,114,31,160,31,49,31,144,31,3,31,3,30,102,31,132,31,216,31,55,31,55,30,55,29,52,31,12,31,12,30,44,31,16,31,160,31,39,31,227,31,155,31,66,31,195,31,51,31,14,31,180,31,103,31,122,31,122,30,122,29,179,31,78,31,85,31,130,31,125,31,132,31,132,30,186,31,100,31,100,30,242,31,243,31,168,31,107,31,78,31,18,31,18,30,26,31,99,31,230,31,71,31,227,31,123,31,70,31,20,31,216,31,156,31,106,31,161,31,95,31,95,30,30,31,180,31,168,31,209,31,19,31,207,31,207,30,134,31,88,31,122,31,5,31,5,30,123,31,121,31,28,31,212,31,134,31,134,30,18,31,18,30,64,31,64,30,131,31,49,31,69,31,154,31,38,31,156,31,156,30,153,31,236,31,159,31,128,31,23,31,133,31,133,30,49,31,92,31,186,31,59,31,147,31,80,31,181,31,181,30,12,31,112,31,180,31,179,31,107,31,107,30,112,31,3,31,119,31,43,31,192,31,96,31,83,31,185,31,88,31,24,31,164,31,59,31,112,31,79,31,16,31,101,31,174,31,177,31,27,31,178,31,123,31,161,31,68,31,119,31,119,30,119,29,107,31,252,31,30,31,30,30,30,29,201,31,156,31,79,31,23,31,23,30,219,31,219,30,206,31,206,30,206,29,127,31,116,31,45,31,45,30,90,31,71,31,199,31,12,31,142,31,106,31,197,31,51,31,30,31,201,31,38,31,186,31,86,31,86,30,100,31,100,30,7,31,226,31,49,31,132,31,216,31,8,31,49,31,49,30,95,31,148,31,40,31,153,31,177,31,231,31,231,30,163,31,3,31,230,31,5,31,95,31,107,31,107,30,9,31,13,31,230,31,230,30,239,31,187,31,88,31,88,30,159,31,199,31,61,31,61,30,27,31,89,31,171,31,42,31,42,30,42,29,89,31,85,31,195,31,212,31,13,31,147,31,116,31,116,30,116,29,141,31,253,31,253,30,158,31,58,31,149,31,166,31,166,30,166,29,13,31,13,30,22,31,220,31,220,30,31,31,102,31,133,31,22,31,105,31,76,31,143,31,124,31,124,30,34,31,12,31,76,31,21,31,222,31,129,31,250,31,34,31,139,31,74,31,9,31,141,31,4,31,93,31,15,31,178,31,252,31,64,31,29,31,17,31,252,31,209,31,8,31,8,30,237,31,68,31,191,31,201,31,106,31,139,31,35,31,167,31,169,31,42,31,240,31,224,31,14,31,14,30,186,31,48,31,113,31,243,31,32,31,227,31,227,30,125,31,46,31,46,30,46,29,231,31,27,31,223,31,68,31,68,30,247,31,17,31,17,30,225,31,68,31,174,31,230,31,87,31,130,31,205,31,209,31,157,31,226,31,226,30,85,31,15,31,15,30,101,31,213,31,41,31,41,30,45,31,239,31,144,31,54,31,30,31,172,31,225,31,75,31,11,31,245,31,223,31,62,31,37,31,37,30,209,31,31,31,208,31,207,31,146,31,35,31,41,31,182,31,131,31,118,31,151,31,98,31,96,31,178,31,128,31,51,31,163,31,29,31,29,30,98,31,149,31,113,31,113,30,222,31,222,30,15,31,57,31,57,30,56,31,95,31,182,31,182,30,182,29,96,31,159,31,252,31,57,31,128,31,23,31,94,31,135,31,210,31,10,31,178,31,228,31,236,31,236,30,18,31,18,30,220,31,245,31,146,31,228,31,63,31,63,30,128,31,255,31,117,31,149,31,192,31,192,30,93,31,164,31,216,31,40,31,217,31,153,31,153,30,153,29,131,31,131,30,92,31,126,31,44,31,144,31,144,30,101,31,185,31,15,31,125,31,125,30,126,31,126,30,126,29,66,31,243,31,73,31,73,30,107,31,107,30,107,29,77,31,213,31,238,31,208,31,208,30,20,31,159,31,137,31,32,31,93,31,93,30,247,31,137,31,232,31,232,30,54,31,243,31,168,31,121,31,113,31,82,31,135,31,21,31,105,31,105,31,22,31,90,31,90,30,224,31,234,31,196,31,40,31,69,31,69,30,105,31,105,30,30,31,198,31,213,31,41,31,41,30,206,31,206,30,110,31,79,31,79,30,139,31,63,31,202,31,244,31,229,31,8,31,184,31,27,31,25,31,152,31,120,31,255,31,26,31,218,31,141,31,241,31,49,31,173,31,247,31,16,31,49,31,169,31,142,31,209,31,161,31,70,31,192,31,197,31,85,31,49,31,46,31,46,30,70,31,88,31,243,31,50,31,253,31,221,31,221,30,31,31,31,30,11,31,11,30,72,31,165,31,1,31,48,31,48,30,195,31,29,31,10,31,129,31,177,31,225,31,94,31,39,31,188,31,239,31,124,31,45,31,134,31,28,31,27,31,48,31,91,31,128,31,128,30,213,31,213,30,25,31,59,31,1,31,128,31,218,31,28,31,41,31,41,30,136,31,227,31,227,30,238,31,50,31,139,31,139,30,128,31,82,31,85,31,56,31,61,31,56,31,142,31,142,30,193,31,180,31,114,31,114,30,114,29,120,31,130,31,72,31,15,31,49,31,199,31,184,31,54,31,142,31,67,31,41,31,211,31,117,31,133,31,148,31,66,31,53,31,124,31,24,31,2,31,129,31,130,31,130,30,82,31,63,31,162,31,162,30,27,31,27,30,27,29,245,31,225,31,78,31,78,30,124,31,40,31,13,31,204,31,156,31,230,31,5,31,147,31,55,31,204,31,188,31,209,31,86,31,77,31,53,31,199,31,30,31,30,30,184,31,49,31,39,31,210,31,52,31,235,31,22,31,84,31,20,31,25,31,1,31,1,31,33,31,34,31,3,31,203,31,203,30,203,29,180,31,190,31,252,31,228,31,228,30,58,31,144,31,182,31,182,30,238,31,238,30,92,31,244,31,205,31,245,31,161,31,45,31,147,31,118,31,250,31,239,31,239,30,149,31,149,30,164,31,225,31,51,31,101,31,106,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
