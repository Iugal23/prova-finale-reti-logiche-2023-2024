-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 302;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (127,0,0,0,47,0,153,0,0,0,0,0,59,0,26,0,0,0,184,0,201,0,199,0,57,0,0,0,8,0,19,0,43,0,117,0,171,0,74,0,24,0,248,0,225,0,0,0,152,0,244,0,6,0,213,0,199,0,145,0,150,0,0,0,1,0,65,0,149,0,201,0,1,0,0,0,97,0,0,0,29,0,127,0,0,0,203,0,0,0,0,0,218,0,0,0,216,0,155,0,0,0,0,0,67,0,0,0,44,0,95,0,187,0,156,0,24,0,100,0,32,0,230,0,25,0,75,0,72,0,51,0,0,0,157,0,0,0,255,0,142,0,145,0,0,0,0,0,137,0,39,0,20,0,0,0,0,0,236,0,33,0,141,0,129,0,37,0,250,0,122,0,187,0,222,0,0,0,251,0,242,0,0,0,244,0,36,0,22,0,21,0,9,0,0,0,0,0,55,0,4,0,168,0,112,0,79,0,181,0,215,0,119,0,66,0,75,0,26,0,34,0,177,0,68,0,215,0,225,0,103,0,0,0,202,0,0,0,178,0,241,0,200,0,0,0,1,0,97,0,112,0,218,0,132,0,180,0,0,0,0,0,123,0,192,0,168,0,0,0,42,0,69,0,107,0,16,0,12,0,47,0,212,0,94,0,160,0,36,0,192,0,73,0,0,0,243,0,124,0,0,0,189,0,83,0,43,0,80,0,155,0,120,0,10,0,183,0,206,0,91,0,129,0,120,0,108,0,42,0,59,0,52,0,0,0,139,0,199,0,0,0,246,0,20,0,179,0,0,0,177,0,228,0,0,0,99,0,109,0,61,0,42,0,0,0,131,0,161,0,37,0,0,0,0,0,4,0,33,0,119,0,189,0,162,0,56,0,0,0,253,0,249,0,0,0,0,0,78,0,0,0,95,0,96,0,11,0,13,0,142,0,96,0,0,0,80,0,0,0,99,0,0,0,0,0,216,0,171,0,206,0,0,0,0,0,230,0,186,0,122,0,31,0,18,0,85,0,175,0,207,0,4,0,250,0,179,0,205,0,113,0,0,0,18,0,47,0,247,0,73,0,68,0,146,0,0,0,235,0,243,0,0,0,178,0,19,0,150,0,179,0,0,0,186,0,0,0,3,0,87,0,59,0,21,0,174,0,232,0,36,0,0,0,170,0,38,0,0,0,250,0,118,0,0,0,0,0,97,0,132,0,98,0,20,0,238,0,176,0,61,0,0,0,201,0,36,0,151,0,0,0,209,0,145,0,0,0,74,0,0,0,0,0,24,0,0,0,73,0,0,0,0,0,55,0,106,0,145,0,22,0,157,0,183,0,59,0,228,0,183,0,252,0,144,0,250,0,70,0,150,0,220,0);
signal scenario_full  : scenario_type := (127,31,127,30,47,31,153,31,153,30,153,29,59,31,26,31,26,30,184,31,201,31,199,31,57,31,57,30,8,31,19,31,43,31,117,31,171,31,74,31,24,31,248,31,225,31,225,30,152,31,244,31,6,31,213,31,199,31,145,31,150,31,150,30,1,31,65,31,149,31,201,31,1,31,1,30,97,31,97,30,29,31,127,31,127,30,203,31,203,30,203,29,218,31,218,30,216,31,155,31,155,30,155,29,67,31,67,30,44,31,95,31,187,31,156,31,24,31,100,31,32,31,230,31,25,31,75,31,72,31,51,31,51,30,157,31,157,30,255,31,142,31,145,31,145,30,145,29,137,31,39,31,20,31,20,30,20,29,236,31,33,31,141,31,129,31,37,31,250,31,122,31,187,31,222,31,222,30,251,31,242,31,242,30,244,31,36,31,22,31,21,31,9,31,9,30,9,29,55,31,4,31,168,31,112,31,79,31,181,31,215,31,119,31,66,31,75,31,26,31,34,31,177,31,68,31,215,31,225,31,103,31,103,30,202,31,202,30,178,31,241,31,200,31,200,30,1,31,97,31,112,31,218,31,132,31,180,31,180,30,180,29,123,31,192,31,168,31,168,30,42,31,69,31,107,31,16,31,12,31,47,31,212,31,94,31,160,31,36,31,192,31,73,31,73,30,243,31,124,31,124,30,189,31,83,31,43,31,80,31,155,31,120,31,10,31,183,31,206,31,91,31,129,31,120,31,108,31,42,31,59,31,52,31,52,30,139,31,199,31,199,30,246,31,20,31,179,31,179,30,177,31,228,31,228,30,99,31,109,31,61,31,42,31,42,30,131,31,161,31,37,31,37,30,37,29,4,31,33,31,119,31,189,31,162,31,56,31,56,30,253,31,249,31,249,30,249,29,78,31,78,30,95,31,96,31,11,31,13,31,142,31,96,31,96,30,80,31,80,30,99,31,99,30,99,29,216,31,171,31,206,31,206,30,206,29,230,31,186,31,122,31,31,31,18,31,85,31,175,31,207,31,4,31,250,31,179,31,205,31,113,31,113,30,18,31,47,31,247,31,73,31,68,31,146,31,146,30,235,31,243,31,243,30,178,31,19,31,150,31,179,31,179,30,186,31,186,30,3,31,87,31,59,31,21,31,174,31,232,31,36,31,36,30,170,31,38,31,38,30,250,31,118,31,118,30,118,29,97,31,132,31,98,31,20,31,238,31,176,31,61,31,61,30,201,31,36,31,151,31,151,30,209,31,145,31,145,30,74,31,74,30,74,29,24,31,24,30,73,31,73,30,73,29,55,31,106,31,145,31,22,31,157,31,183,31,59,31,228,31,183,31,252,31,144,31,250,31,70,31,150,31,220,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
