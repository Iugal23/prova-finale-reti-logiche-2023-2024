-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_960 is
end project_tb_960;

architecture project_tb_arch_960 of project_tb_960 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 973;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (171,0,114,0,182,0,53,0,0,0,0,0,221,0,186,0,0,0,217,0,78,0,143,0,189,0,147,0,232,0,60,0,186,0,51,0,52,0,0,0,220,0,161,0,153,0,250,0,8,0,91,0,250,0,0,0,0,0,88,0,215,0,255,0,229,0,0,0,173,0,108,0,15,0,97,0,18,0,188,0,225,0,133,0,0,0,105,0,128,0,102,0,31,0,60,0,144,0,0,0,124,0,144,0,0,0,98,0,171,0,30,0,218,0,225,0,52,0,116,0,4,0,126,0,119,0,220,0,224,0,0,0,111,0,222,0,150,0,0,0,0,0,71,0,38,0,0,0,0,0,46,0,214,0,236,0,44,0,0,0,0,0,151,0,190,0,162,0,151,0,9,0,41,0,209,0,41,0,0,0,191,0,234,0,0,0,81,0,69,0,87,0,84,0,46,0,190,0,0,0,0,0,180,0,74,0,253,0,104,0,0,0,27,0,232,0,199,0,219,0,16,0,0,0,0,0,122,0,88,0,0,0,253,0,57,0,16,0,0,0,19,0,29,0,99,0,120,0,89,0,53,0,212,0,0,0,121,0,67,0,134,0,164,0,0,0,198,0,166,0,131,0,35,0,182,0,253,0,229,0,169,0,133,0,107,0,250,0,21,0,0,0,211,0,148,0,125,0,57,0,137,0,188,0,98,0,96,0,105,0,0,0,55,0,16,0,15,0,78,0,133,0,3,0,65,0,191,0,79,0,40,0,0,0,0,0,241,0,183,0,26,0,226,0,15,0,0,0,31,0,0,0,0,0,45,0,0,0,173,0,94,0,50,0,120,0,67,0,48,0,136,0,15,0,40,0,252,0,0,0,215,0,0,0,237,0,230,0,121,0,242,0,142,0,255,0,222,0,165,0,56,0,91,0,20,0,74,0,117,0,0,0,0,0,79,0,88,0,112,0,252,0,207,0,36,0,138,0,8,0,208,0,0,0,168,0,207,0,67,0,155,0,193,0,203,0,171,0,50,0,251,0,0,0,227,0,137,0,116,0,182,0,132,0,32,0,53,0,238,0,161,0,143,0,193,0,240,0,0,0,0,0,56,0,46,0,139,0,0,0,0,0,0,0,133,0,164,0,111,0,134,0,65,0,236,0,187,0,190,0,169,0,89,0,182,0,130,0,0,0,185,0,199,0,243,0,88,0,250,0,247,0,0,0,81,0,255,0,68,0,41,0,201,0,0,0,198,0,0,0,51,0,12,0,46,0,117,0,129,0,94,0,41,0,197,0,74,0,0,0,60,0,106,0,112,0,237,0,91,0,104,0,47,0,50,0,166,0,239,0,148,0,0,0,44,0,225,0,56,0,0,0,244,0,40,0,52,0,33,0,0,0,227,0,184,0,252,0,210,0,0,0,0,0,0,0,0,0,79,0,249,0,25,0,0,0,211,0,0,0,233,0,55,0,47,0,175,0,149,0,0,0,143,0,245,0,0,0,120,0,6,0,0,0,26,0,25,0,224,0,125,0,230,0,222,0,181,0,114,0,0,0,117,0,148,0,164,0,0,0,0,0,224,0,0,0,43,0,34,0,62,0,74,0,162,0,199,0,172,0,126,0,52,0,141,0,174,0,232,0,0,0,191,0,195,0,220,0,135,0,46,0,51,0,39,0,73,0,0,0,167,0,234,0,105,0,0,0,29,0,0,0,203,0,111,0,206,0,130,0,0,0,188,0,239,0,145,0,87,0,32,0,0,0,131,0,40,0,33,0,135,0,0,0,0,0,136,0,183,0,32,0,150,0,150,0,54,0,70,0,83,0,218,0,255,0,85,0,82,0,62,0,87,0,200,0,85,0,139,0,6,0,189,0,0,0,247,0,223,0,127,0,24,0,241,0,110,0,0,0,12,0,155,0,20,0,0,0,69,0,0,0,52,0,236,0,0,0,176,0,0,0,155,0,0,0,255,0,89,0,80,0,0,0,10,0,220,0,175,0,152,0,61,0,0,0,57,0,180,0,148,0,69,0,0,0,143,0,201,0,0,0,205,0,131,0,216,0,178,0,189,0,47,0,74,0,34,0,215,0,217,0,164,0,250,0,237,0,225,0,31,0,98,0,233,0,49,0,0,0,0,0,32,0,0,0,252,0,91,0,141,0,24,0,121,0,0,0,0,0,0,0,0,0,7,0,0,0,0,0,0,0,225,0,0,0,134,0,0,0,0,0,95,0,133,0,246,0,232,0,103,0,27,0,37,0,105,0,0,0,0,0,133,0,130,0,59,0,22,0,193,0,0,0,74,0,4,0,52,0,156,0,134,0,224,0,0,0,175,0,71,0,63,0,96,0,230,0,224,0,79,0,102,0,135,0,71,0,0,0,99,0,253,0,245,0,168,0,0,0,144,0,243,0,0,0,127,0,221,0,186,0,125,0,0,0,97,0,107,0,24,0,233,0,147,0,200,0,36,0,30,0,88,0,239,0,58,0,187,0,190,0,76,0,175,0,182,0,170,0,0,0,0,0,132,0,205,0,230,0,133,0,178,0,190,0,62,0,216,0,22,0,137,0,100,0,247,0,14,0,102,0,140,0,114,0,0,0,166,0,61,0,77,0,22,0,111,0,171,0,54,0,20,0,253,0,141,0,175,0,227,0,239,0,96,0,206,0,136,0,189,0,98,0,188,0,172,0,60,0,21,0,186,0,190,0,153,0,159,0,135,0,227,0,0,0,19,0,32,0,66,0,0,0,32,0,0,0,53,0,28,0,0,0,189,0,162,0,144,0,192,0,60,0,96,0,168,0,0,0,192,0,232,0,180,0,132,0,0,0,207,0,91,0,186,0,0,0,5,0,176,0,102,0,139,0,241,0,5,0,99,0,225,0,148,0,0,0,0,0,13,0,214,0,72,0,169,0,69,0,90,0,228,0,0,0,122,0,171,0,98,0,150,0,48,0,90,0,211,0,37,0,0,0,78,0,106,0,179,0,97,0,0,0,0,0,252,0,35,0,140,0,0,0,26,0,194,0,60,0,235,0,131,0,79,0,195,0,45,0,121,0,180,0,66,0,0,0,180,0,113,0,0,0,194,0,68,0,0,0,0,0,42,0,186,0,0,0,81,0,0,0,141,0,30,0,0,0,108,0,252,0,123,0,114,0,112,0,191,0,241,0,234,0,35,0,0,0,0,0,83,0,0,0,132,0,133,0,71,0,0,0,0,0,0,0,0,0,84,0,123,0,189,0,0,0,0,0,242,0,0,0,0,0,73,0,0,0,139,0,0,0,0,0,94,0,0,0,65,0,165,0,112,0,200,0,33,0,203,0,0,0,197,0,0,0,39,0,42,0,0,0,135,0,190,0,140,0,210,0,49,0,156,0,167,0,14,0,0,0,230,0,65,0,237,0,162,0,203,0,108,0,56,0,34,0,0,0,196,0,73,0,73,0,93,0,53,0,202,0,17,0,205,0,97,0,219,0,16,0,166,0,0,0,194,0,245,0,0,0,0,0,0,0,0,0,83,0,50,0,120,0,130,0,200,0,243,0,162,0,239,0,0,0,199,0,82,0,223,0,20,0,250,0,98,0,0,0,160,0,193,0,220,0,23,0,77,0,98,0,43,0,0,0,0,0,43,0,0,0,208,0,0,0,3,0,0,0,0,0,0,0,100,0,70,0,110,0,0,0,10,0,132,0,98,0,6,0,165,0,132,0,248,0,34,0,102,0,198,0,200,0,9,0,28,0,65,0,162,0,208,0,20,0,0,0,128,0,22,0,245,0,26,0,40,0,153,0,64,0,249,0,0,0,47,0,208,0,223,0,221,0,0,0,0,0,213,0,0,0,0,0,13,0,155,0,79,0,0,0,239,0,17,0,113,0,192,0,0,0,20,0,42,0,106,0,207,0,0,0,121,0,0,0,92,0,214,0,247,0,0,0,226,0,241,0,132,0,92,0,115,0,60,0,84,0,253,0,126,0,241,0,0,0,3,0,0,0,0,0,0,0,39,0,82,0,0,0,59,0,59,0,243,0,217,0,183,0,122,0,144,0,100,0,146,0,197,0,0,0,202,0,62,0,214,0,196,0,45,0,147,0,239,0,198,0,75,0,0,0,29,0,215,0,181,0,0,0,0,0,136,0,29,0,175,0,54,0,8,0,53,0,0,0,0,0,188,0,88,0,15,0,0,0,0,0,0,0,94,0,0,0,90,0,153,0,153,0,189,0,129,0,209,0,247,0,0,0,95,0,0,0,120,0,0,0,53,0,3,0,0,0,45,0,0,0,0,0,46,0,125,0,56,0,50,0,36,0,44,0,91,0,207,0,194,0,24,0,174,0,249,0,127,0,39,0,68,0,0,0,192,0,102,0,252,0,161,0,148,0,0,0,255,0,0,0);
signal scenario_full  : scenario_type := (171,31,114,31,182,31,53,31,53,30,53,29,221,31,186,31,186,30,217,31,78,31,143,31,189,31,147,31,232,31,60,31,186,31,51,31,52,31,52,30,220,31,161,31,153,31,250,31,8,31,91,31,250,31,250,30,250,29,88,31,215,31,255,31,229,31,229,30,173,31,108,31,15,31,97,31,18,31,188,31,225,31,133,31,133,30,105,31,128,31,102,31,31,31,60,31,144,31,144,30,124,31,144,31,144,30,98,31,171,31,30,31,218,31,225,31,52,31,116,31,4,31,126,31,119,31,220,31,224,31,224,30,111,31,222,31,150,31,150,30,150,29,71,31,38,31,38,30,38,29,46,31,214,31,236,31,44,31,44,30,44,29,151,31,190,31,162,31,151,31,9,31,41,31,209,31,41,31,41,30,191,31,234,31,234,30,81,31,69,31,87,31,84,31,46,31,190,31,190,30,190,29,180,31,74,31,253,31,104,31,104,30,27,31,232,31,199,31,219,31,16,31,16,30,16,29,122,31,88,31,88,30,253,31,57,31,16,31,16,30,19,31,29,31,99,31,120,31,89,31,53,31,212,31,212,30,121,31,67,31,134,31,164,31,164,30,198,31,166,31,131,31,35,31,182,31,253,31,229,31,169,31,133,31,107,31,250,31,21,31,21,30,211,31,148,31,125,31,57,31,137,31,188,31,98,31,96,31,105,31,105,30,55,31,16,31,15,31,78,31,133,31,3,31,65,31,191,31,79,31,40,31,40,30,40,29,241,31,183,31,26,31,226,31,15,31,15,30,31,31,31,30,31,29,45,31,45,30,173,31,94,31,50,31,120,31,67,31,48,31,136,31,15,31,40,31,252,31,252,30,215,31,215,30,237,31,230,31,121,31,242,31,142,31,255,31,222,31,165,31,56,31,91,31,20,31,74,31,117,31,117,30,117,29,79,31,88,31,112,31,252,31,207,31,36,31,138,31,8,31,208,31,208,30,168,31,207,31,67,31,155,31,193,31,203,31,171,31,50,31,251,31,251,30,227,31,137,31,116,31,182,31,132,31,32,31,53,31,238,31,161,31,143,31,193,31,240,31,240,30,240,29,56,31,46,31,139,31,139,30,139,29,139,28,133,31,164,31,111,31,134,31,65,31,236,31,187,31,190,31,169,31,89,31,182,31,130,31,130,30,185,31,199,31,243,31,88,31,250,31,247,31,247,30,81,31,255,31,68,31,41,31,201,31,201,30,198,31,198,30,51,31,12,31,46,31,117,31,129,31,94,31,41,31,197,31,74,31,74,30,60,31,106,31,112,31,237,31,91,31,104,31,47,31,50,31,166,31,239,31,148,31,148,30,44,31,225,31,56,31,56,30,244,31,40,31,52,31,33,31,33,30,227,31,184,31,252,31,210,31,210,30,210,29,210,28,210,27,79,31,249,31,25,31,25,30,211,31,211,30,233,31,55,31,47,31,175,31,149,31,149,30,143,31,245,31,245,30,120,31,6,31,6,30,26,31,25,31,224,31,125,31,230,31,222,31,181,31,114,31,114,30,117,31,148,31,164,31,164,30,164,29,224,31,224,30,43,31,34,31,62,31,74,31,162,31,199,31,172,31,126,31,52,31,141,31,174,31,232,31,232,30,191,31,195,31,220,31,135,31,46,31,51,31,39,31,73,31,73,30,167,31,234,31,105,31,105,30,29,31,29,30,203,31,111,31,206,31,130,31,130,30,188,31,239,31,145,31,87,31,32,31,32,30,131,31,40,31,33,31,135,31,135,30,135,29,136,31,183,31,32,31,150,31,150,31,54,31,70,31,83,31,218,31,255,31,85,31,82,31,62,31,87,31,200,31,85,31,139,31,6,31,189,31,189,30,247,31,223,31,127,31,24,31,241,31,110,31,110,30,12,31,155,31,20,31,20,30,69,31,69,30,52,31,236,31,236,30,176,31,176,30,155,31,155,30,255,31,89,31,80,31,80,30,10,31,220,31,175,31,152,31,61,31,61,30,57,31,180,31,148,31,69,31,69,30,143,31,201,31,201,30,205,31,131,31,216,31,178,31,189,31,47,31,74,31,34,31,215,31,217,31,164,31,250,31,237,31,225,31,31,31,98,31,233,31,49,31,49,30,49,29,32,31,32,30,252,31,91,31,141,31,24,31,121,31,121,30,121,29,121,28,121,27,7,31,7,30,7,29,7,28,225,31,225,30,134,31,134,30,134,29,95,31,133,31,246,31,232,31,103,31,27,31,37,31,105,31,105,30,105,29,133,31,130,31,59,31,22,31,193,31,193,30,74,31,4,31,52,31,156,31,134,31,224,31,224,30,175,31,71,31,63,31,96,31,230,31,224,31,79,31,102,31,135,31,71,31,71,30,99,31,253,31,245,31,168,31,168,30,144,31,243,31,243,30,127,31,221,31,186,31,125,31,125,30,97,31,107,31,24,31,233,31,147,31,200,31,36,31,30,31,88,31,239,31,58,31,187,31,190,31,76,31,175,31,182,31,170,31,170,30,170,29,132,31,205,31,230,31,133,31,178,31,190,31,62,31,216,31,22,31,137,31,100,31,247,31,14,31,102,31,140,31,114,31,114,30,166,31,61,31,77,31,22,31,111,31,171,31,54,31,20,31,253,31,141,31,175,31,227,31,239,31,96,31,206,31,136,31,189,31,98,31,188,31,172,31,60,31,21,31,186,31,190,31,153,31,159,31,135,31,227,31,227,30,19,31,32,31,66,31,66,30,32,31,32,30,53,31,28,31,28,30,189,31,162,31,144,31,192,31,60,31,96,31,168,31,168,30,192,31,232,31,180,31,132,31,132,30,207,31,91,31,186,31,186,30,5,31,176,31,102,31,139,31,241,31,5,31,99,31,225,31,148,31,148,30,148,29,13,31,214,31,72,31,169,31,69,31,90,31,228,31,228,30,122,31,171,31,98,31,150,31,48,31,90,31,211,31,37,31,37,30,78,31,106,31,179,31,97,31,97,30,97,29,252,31,35,31,140,31,140,30,26,31,194,31,60,31,235,31,131,31,79,31,195,31,45,31,121,31,180,31,66,31,66,30,180,31,113,31,113,30,194,31,68,31,68,30,68,29,42,31,186,31,186,30,81,31,81,30,141,31,30,31,30,30,108,31,252,31,123,31,114,31,112,31,191,31,241,31,234,31,35,31,35,30,35,29,83,31,83,30,132,31,133,31,71,31,71,30,71,29,71,28,71,27,84,31,123,31,189,31,189,30,189,29,242,31,242,30,242,29,73,31,73,30,139,31,139,30,139,29,94,31,94,30,65,31,165,31,112,31,200,31,33,31,203,31,203,30,197,31,197,30,39,31,42,31,42,30,135,31,190,31,140,31,210,31,49,31,156,31,167,31,14,31,14,30,230,31,65,31,237,31,162,31,203,31,108,31,56,31,34,31,34,30,196,31,73,31,73,31,93,31,53,31,202,31,17,31,205,31,97,31,219,31,16,31,166,31,166,30,194,31,245,31,245,30,245,29,245,28,245,27,83,31,50,31,120,31,130,31,200,31,243,31,162,31,239,31,239,30,199,31,82,31,223,31,20,31,250,31,98,31,98,30,160,31,193,31,220,31,23,31,77,31,98,31,43,31,43,30,43,29,43,31,43,30,208,31,208,30,3,31,3,30,3,29,3,28,100,31,70,31,110,31,110,30,10,31,132,31,98,31,6,31,165,31,132,31,248,31,34,31,102,31,198,31,200,31,9,31,28,31,65,31,162,31,208,31,20,31,20,30,128,31,22,31,245,31,26,31,40,31,153,31,64,31,249,31,249,30,47,31,208,31,223,31,221,31,221,30,221,29,213,31,213,30,213,29,13,31,155,31,79,31,79,30,239,31,17,31,113,31,192,31,192,30,20,31,42,31,106,31,207,31,207,30,121,31,121,30,92,31,214,31,247,31,247,30,226,31,241,31,132,31,92,31,115,31,60,31,84,31,253,31,126,31,241,31,241,30,3,31,3,30,3,29,3,28,39,31,82,31,82,30,59,31,59,31,243,31,217,31,183,31,122,31,144,31,100,31,146,31,197,31,197,30,202,31,62,31,214,31,196,31,45,31,147,31,239,31,198,31,75,31,75,30,29,31,215,31,181,31,181,30,181,29,136,31,29,31,175,31,54,31,8,31,53,31,53,30,53,29,188,31,88,31,15,31,15,30,15,29,15,28,94,31,94,30,90,31,153,31,153,31,189,31,129,31,209,31,247,31,247,30,95,31,95,30,120,31,120,30,53,31,3,31,3,30,45,31,45,30,45,29,46,31,125,31,56,31,50,31,36,31,44,31,91,31,207,31,194,31,24,31,174,31,249,31,127,31,39,31,68,31,68,30,192,31,102,31,252,31,161,31,148,31,148,30,255,31,255,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
