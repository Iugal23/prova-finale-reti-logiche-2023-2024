-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 707;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (159,0,85,0,90,0,210,0,23,0,70,0,192,0,237,0,78,0,71,0,145,0,203,0,64,0,105,0,0,0,117,0,167,0,0,0,143,0,0,0,176,0,18,0,99,0,26,0,99,0,0,0,236,0,0,0,72,0,0,0,33,0,214,0,106,0,227,0,0,0,153,0,129,0,97,0,89,0,0,0,41,0,233,0,52,0,168,0,65,0,64,0,206,0,79,0,16,0,103,0,166,0,135,0,27,0,123,0,35,0,0,0,176,0,0,0,245,0,90,0,0,0,186,0,208,0,31,0,232,0,98,0,172,0,150,0,0,0,173,0,2,0,152,0,6,0,136,0,42,0,244,0,0,0,0,0,0,0,33,0,84,0,144,0,219,0,144,0,32,0,221,0,0,0,65,0,211,0,0,0,235,0,41,0,208,0,74,0,203,0,3,0,86,0,228,0,0,0,0,0,199,0,171,0,60,0,31,0,189,0,0,0,0,0,3,0,107,0,9,0,120,0,217,0,92,0,101,0,96,0,0,0,175,0,8,0,0,0,0,0,0,0,5,0,122,0,172,0,128,0,0,0,198,0,183,0,9,0,48,0,0,0,229,0,166,0,0,0,0,0,203,0,45,0,3,0,200,0,164,0,161,0,30,0,36,0,145,0,188,0,0,0,152,0,0,0,28,0,183,0,208,0,0,0,185,0,201,0,0,0,210,0,107,0,183,0,174,0,89,0,218,0,183,0,200,0,0,0,103,0,174,0,115,0,0,0,243,0,61,0,15,0,4,0,118,0,61,0,192,0,204,0,111,0,119,0,214,0,79,0,9,0,170,0,126,0,221,0,38,0,39,0,129,0,168,0,16,0,0,0,130,0,0,0,116,0,71,0,243,0,120,0,0,0,156,0,95,0,155,0,0,0,0,0,51,0,31,0,0,0,248,0,36,0,0,0,94,0,102,0,248,0,76,0,47,0,0,0,90,0,203,0,207,0,79,0,36,0,72,0,129,0,151,0,51,0,28,0,186,0,108,0,0,0,93,0,227,0,132,0,18,0,20,0,222,0,180,0,14,0,0,0,20,0,0,0,19,0,122,0,173,0,174,0,61,0,0,0,59,0,0,0,154,0,191,0,171,0,240,0,4,0,227,0,0,0,29,0,40,0,164,0,0,0,0,0,3,0,43,0,10,0,28,0,105,0,21,0,89,0,138,0,0,0,94,0,7,0,75,0,208,0,78,0,34,0,10,0,216,0,9,0,235,0,0,0,146,0,168,0,0,0,230,0,43,0,210,0,117,0,81,0,79,0,99,0,171,0,50,0,75,0,44,0,204,0,0,0,214,0,0,0,67,0,20,0,12,0,184,0,185,0,197,0,194,0,80,0,236,0,59,0,137,0,126,0,128,0,96,0,0,0,0,0,0,0,168,0,12,0,188,0,0,0,129,0,242,0,178,0,116,0,39,0,21,0,101,0,78,0,160,0,250,0,0,0,16,0,17,0,223,0,250,0,115,0,71,0,193,0,131,0,0,0,78,0,0,0,0,0,177,0,243,0,58,0,0,0,35,0,61,0,69,0,15,0,53,0,191,0,137,0,186,0,83,0,0,0,89,0,213,0,80,0,174,0,70,0,169,0,107,0,0,0,190,0,131,0,14,0,52,0,203,0,99,0,190,0,94,0,207,0,227,0,9,0,41,0,94,0,1,0,0,0,115,0,95,0,193,0,227,0,158,0,179,0,27,0,160,0,249,0,108,0,94,0,48,0,141,0,160,0,220,0,0,0,20,0,27,0,247,0,0,0,0,0,139,0,0,0,0,0,61,0,36,0,0,0,30,0,224,0,0,0,175,0,134,0,128,0,213,0,92,0,0,0,0,0,230,0,16,0,48,0,201,0,0,0,71,0,218,0,0,0,74,0,85,0,235,0,177,0,216,0,85,0,111,0,231,0,218,0,229,0,253,0,30,0,149,0,25,0,5,0,0,0,0,0,81,0,0,0,29,0,0,0,11,0,0,0,0,0,191,0,140,0,0,0,244,0,221,0,93,0,59,0,67,0,133,0,11,0,11,0,0,0,143,0,0,0,238,0,15,0,206,0,97,0,39,0,136,0,238,0,135,0,245,0,62,0,47,0,0,0,0,0,0,0,126,0,60,0,195,0,246,0,0,0,238,0,148,0,165,0,144,0,54,0,135,0,190,0,0,0,187,0,81,0,208,0,88,0,0,0,70,0,206,0,0,0,168,0,128,0,118,0,0,0,134,0,131,0,94,0,140,0,135,0,128,0,90,0,200,0,115,0,78,0,227,0,242,0,130,0,230,0,13,0,188,0,252,0,0,0,243,0,39,0,237,0,186,0,11,0,178,0,253,0,193,0,72,0,193,0,249,0,6,0,0,0,0,0,0,0,240,0,207,0,90,0,0,0,121,0,60,0,18,0,211,0,0,0,0,0,0,0,163,0,77,0,89,0,0,0,8,0,173,0,226,0,129,0,195,0,0,0,148,0,156,0,254,0,0,0,174,0,0,0,185,0,132,0,246,0,66,0,181,0,186,0,101,0,105,0,104,0,0,0,172,0,142,0,92,0,0,0,22,0,17,0,116,0,106,0,52,0,179,0,247,0,75,0,0,0,88,0,0,0,0,0,230,0,197,0,124,0,133,0,218,0,159,0,105,0,236,0,0,0,101,0,102,0,103,0,150,0,7,0,216,0,175,0,130,0,164,0,240,0,225,0,3,0,33,0,38,0,229,0,0,0,226,0,211,0,54,0,165,0,50,0,239,0,231,0,0,0,88,0,44,0,19,0,83,0,0,0,6,0,115,0,100,0,214,0,102,0,0,0,194,0,113,0,0,0,192,0,0,0,54,0,58,0,168,0,51,0,209,0,105,0,193,0,206,0,240,0,121,0,200,0,222,0,0,0,73,0,183,0,229,0,198,0,132,0,0,0,0,0,119,0,234,0,106,0,0,0,218,0,33,0,142,0,17,0,164,0,0,0,42,0,74,0,100,0,223,0,0,0,0,0,0,0,238,0,194,0,129,0,207,0,158,0,64,0,0,0,0,0,216,0,202,0,0,0,39,0,2,0,106,0,115,0,0,0,0,0,139,0,250,0,201,0,19,0,0,0,146,0,152,0,0,0,0,0,207,0,118,0,0,0,121,0,137,0,219,0,2,0,64,0,141,0,136,0);
signal scenario_full  : scenario_type := (159,31,85,31,90,31,210,31,23,31,70,31,192,31,237,31,78,31,71,31,145,31,203,31,64,31,105,31,105,30,117,31,167,31,167,30,143,31,143,30,176,31,18,31,99,31,26,31,99,31,99,30,236,31,236,30,72,31,72,30,33,31,214,31,106,31,227,31,227,30,153,31,129,31,97,31,89,31,89,30,41,31,233,31,52,31,168,31,65,31,64,31,206,31,79,31,16,31,103,31,166,31,135,31,27,31,123,31,35,31,35,30,176,31,176,30,245,31,90,31,90,30,186,31,208,31,31,31,232,31,98,31,172,31,150,31,150,30,173,31,2,31,152,31,6,31,136,31,42,31,244,31,244,30,244,29,244,28,33,31,84,31,144,31,219,31,144,31,32,31,221,31,221,30,65,31,211,31,211,30,235,31,41,31,208,31,74,31,203,31,3,31,86,31,228,31,228,30,228,29,199,31,171,31,60,31,31,31,189,31,189,30,189,29,3,31,107,31,9,31,120,31,217,31,92,31,101,31,96,31,96,30,175,31,8,31,8,30,8,29,8,28,5,31,122,31,172,31,128,31,128,30,198,31,183,31,9,31,48,31,48,30,229,31,166,31,166,30,166,29,203,31,45,31,3,31,200,31,164,31,161,31,30,31,36,31,145,31,188,31,188,30,152,31,152,30,28,31,183,31,208,31,208,30,185,31,201,31,201,30,210,31,107,31,183,31,174,31,89,31,218,31,183,31,200,31,200,30,103,31,174,31,115,31,115,30,243,31,61,31,15,31,4,31,118,31,61,31,192,31,204,31,111,31,119,31,214,31,79,31,9,31,170,31,126,31,221,31,38,31,39,31,129,31,168,31,16,31,16,30,130,31,130,30,116,31,71,31,243,31,120,31,120,30,156,31,95,31,155,31,155,30,155,29,51,31,31,31,31,30,248,31,36,31,36,30,94,31,102,31,248,31,76,31,47,31,47,30,90,31,203,31,207,31,79,31,36,31,72,31,129,31,151,31,51,31,28,31,186,31,108,31,108,30,93,31,227,31,132,31,18,31,20,31,222,31,180,31,14,31,14,30,20,31,20,30,19,31,122,31,173,31,174,31,61,31,61,30,59,31,59,30,154,31,191,31,171,31,240,31,4,31,227,31,227,30,29,31,40,31,164,31,164,30,164,29,3,31,43,31,10,31,28,31,105,31,21,31,89,31,138,31,138,30,94,31,7,31,75,31,208,31,78,31,34,31,10,31,216,31,9,31,235,31,235,30,146,31,168,31,168,30,230,31,43,31,210,31,117,31,81,31,79,31,99,31,171,31,50,31,75,31,44,31,204,31,204,30,214,31,214,30,67,31,20,31,12,31,184,31,185,31,197,31,194,31,80,31,236,31,59,31,137,31,126,31,128,31,96,31,96,30,96,29,96,28,168,31,12,31,188,31,188,30,129,31,242,31,178,31,116,31,39,31,21,31,101,31,78,31,160,31,250,31,250,30,16,31,17,31,223,31,250,31,115,31,71,31,193,31,131,31,131,30,78,31,78,30,78,29,177,31,243,31,58,31,58,30,35,31,61,31,69,31,15,31,53,31,191,31,137,31,186,31,83,31,83,30,89,31,213,31,80,31,174,31,70,31,169,31,107,31,107,30,190,31,131,31,14,31,52,31,203,31,99,31,190,31,94,31,207,31,227,31,9,31,41,31,94,31,1,31,1,30,115,31,95,31,193,31,227,31,158,31,179,31,27,31,160,31,249,31,108,31,94,31,48,31,141,31,160,31,220,31,220,30,20,31,27,31,247,31,247,30,247,29,139,31,139,30,139,29,61,31,36,31,36,30,30,31,224,31,224,30,175,31,134,31,128,31,213,31,92,31,92,30,92,29,230,31,16,31,48,31,201,31,201,30,71,31,218,31,218,30,74,31,85,31,235,31,177,31,216,31,85,31,111,31,231,31,218,31,229,31,253,31,30,31,149,31,25,31,5,31,5,30,5,29,81,31,81,30,29,31,29,30,11,31,11,30,11,29,191,31,140,31,140,30,244,31,221,31,93,31,59,31,67,31,133,31,11,31,11,31,11,30,143,31,143,30,238,31,15,31,206,31,97,31,39,31,136,31,238,31,135,31,245,31,62,31,47,31,47,30,47,29,47,28,126,31,60,31,195,31,246,31,246,30,238,31,148,31,165,31,144,31,54,31,135,31,190,31,190,30,187,31,81,31,208,31,88,31,88,30,70,31,206,31,206,30,168,31,128,31,118,31,118,30,134,31,131,31,94,31,140,31,135,31,128,31,90,31,200,31,115,31,78,31,227,31,242,31,130,31,230,31,13,31,188,31,252,31,252,30,243,31,39,31,237,31,186,31,11,31,178,31,253,31,193,31,72,31,193,31,249,31,6,31,6,30,6,29,6,28,240,31,207,31,90,31,90,30,121,31,60,31,18,31,211,31,211,30,211,29,211,28,163,31,77,31,89,31,89,30,8,31,173,31,226,31,129,31,195,31,195,30,148,31,156,31,254,31,254,30,174,31,174,30,185,31,132,31,246,31,66,31,181,31,186,31,101,31,105,31,104,31,104,30,172,31,142,31,92,31,92,30,22,31,17,31,116,31,106,31,52,31,179,31,247,31,75,31,75,30,88,31,88,30,88,29,230,31,197,31,124,31,133,31,218,31,159,31,105,31,236,31,236,30,101,31,102,31,103,31,150,31,7,31,216,31,175,31,130,31,164,31,240,31,225,31,3,31,33,31,38,31,229,31,229,30,226,31,211,31,54,31,165,31,50,31,239,31,231,31,231,30,88,31,44,31,19,31,83,31,83,30,6,31,115,31,100,31,214,31,102,31,102,30,194,31,113,31,113,30,192,31,192,30,54,31,58,31,168,31,51,31,209,31,105,31,193,31,206,31,240,31,121,31,200,31,222,31,222,30,73,31,183,31,229,31,198,31,132,31,132,30,132,29,119,31,234,31,106,31,106,30,218,31,33,31,142,31,17,31,164,31,164,30,42,31,74,31,100,31,223,31,223,30,223,29,223,28,238,31,194,31,129,31,207,31,158,31,64,31,64,30,64,29,216,31,202,31,202,30,39,31,2,31,106,31,115,31,115,30,115,29,139,31,250,31,201,31,19,31,19,30,146,31,152,31,152,30,152,29,207,31,118,31,118,30,121,31,137,31,219,31,2,31,64,31,141,31,136,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
