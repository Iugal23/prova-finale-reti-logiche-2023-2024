-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_271 is
end project_tb_271;

architecture project_tb_arch_271 of project_tb_271 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 332;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (219,0,68,0,2,0,185,0,34,0,153,0,162,0,190,0,228,0,56,0,0,0,177,0,0,0,159,0,205,0,231,0,50,0,123,0,81,0,184,0,28,0,0,0,0,0,36,0,118,0,201,0,61,0,60,0,113,0,91,0,0,0,167,0,202,0,17,0,157,0,76,0,196,0,21,0,30,0,132,0,228,0,1,0,180,0,227,0,251,0,106,0,153,0,29,0,160,0,33,0,104,0,248,0,245,0,161,0,0,0,179,0,56,0,157,0,44,0,44,0,214,0,144,0,186,0,0,0,0,0,80,0,223,0,109,0,16,0,184,0,144,0,239,0,208,0,35,0,196,0,39,0,163,0,0,0,247,0,54,0,150,0,0,0,251,0,81,0,0,0,68,0,193,0,0,0,0,0,93,0,169,0,162,0,188,0,222,0,0,0,0,0,22,0,70,0,167,0,25,0,87,0,0,0,82,0,169,0,0,0,169,0,233,0,73,0,57,0,220,0,0,0,43,0,36,0,0,0,4,0,193,0,235,0,38,0,221,0,252,0,100,0,0,0,0,0,34,0,101,0,250,0,76,0,38,0,55,0,164,0,197,0,179,0,219,0,108,0,253,0,244,0,125,0,144,0,62,0,242,0,156,0,146,0,254,0,210,0,123,0,126,0,160,0,205,0,37,0,106,0,206,0,88,0,0,0,18,0,60,0,185,0,0,0,14,0,0,0,21,0,172,0,40,0,0,0,56,0,0,0,232,0,114,0,186,0,2,0,158,0,200,0,210,0,14,0,56,0,9,0,17,0,15,0,0,0,129,0,76,0,190,0,131,0,138,0,116,0,76,0,0,0,0,0,89,0,199,0,0,0,42,0,0,0,158,0,246,0,19,0,174,0,82,0,184,0,224,0,102,0,0,0,65,0,164,0,132,0,241,0,70,0,10,0,80,0,42,0,145,0,229,0,0,0,210,0,140,0,36,0,10,0,187,0,124,0,0,0,246,0,50,0,150,0,0,0,83,0,0,0,0,0,174,0,161,0,134,0,0,0,9,0,0,0,247,0,247,0,226,0,64,0,53,0,38,0,15,0,116,0,12,0,244,0,19,0,0,0,121,0,224,0,0,0,14,0,17,0,29,0,0,0,77,0,0,0,21,0,0,0,151,0,96,0,131,0,94,0,21,0,150,0,157,0,247,0,208,0,190,0,227,0,141,0,219,0,151,0,180,0,222,0,0,0,0,0,197,0,8,0,137,0,254,0,107,0,240,0,0,0,131,0,172,0,62,0,29,0,56,0,57,0,0,0,34,0,215,0,29,0,187,0,172,0,249,0,207,0,201,0,119,0,14,0,118,0,0,0,107,0,248,0,150,0,236,0,0,0,0,0,0,0,0,0,128,0,0,0,207,0,48,0,233,0,109,0,0,0,239,0,215,0,45,0,19,0,199,0,125,0,10,0,0,0,106,0,102,0,0,0,237,0,72,0,5,0,194,0,111,0,0,0,176,0);
signal scenario_full  : scenario_type := (219,31,68,31,2,31,185,31,34,31,153,31,162,31,190,31,228,31,56,31,56,30,177,31,177,30,159,31,205,31,231,31,50,31,123,31,81,31,184,31,28,31,28,30,28,29,36,31,118,31,201,31,61,31,60,31,113,31,91,31,91,30,167,31,202,31,17,31,157,31,76,31,196,31,21,31,30,31,132,31,228,31,1,31,180,31,227,31,251,31,106,31,153,31,29,31,160,31,33,31,104,31,248,31,245,31,161,31,161,30,179,31,56,31,157,31,44,31,44,31,214,31,144,31,186,31,186,30,186,29,80,31,223,31,109,31,16,31,184,31,144,31,239,31,208,31,35,31,196,31,39,31,163,31,163,30,247,31,54,31,150,31,150,30,251,31,81,31,81,30,68,31,193,31,193,30,193,29,93,31,169,31,162,31,188,31,222,31,222,30,222,29,22,31,70,31,167,31,25,31,87,31,87,30,82,31,169,31,169,30,169,31,233,31,73,31,57,31,220,31,220,30,43,31,36,31,36,30,4,31,193,31,235,31,38,31,221,31,252,31,100,31,100,30,100,29,34,31,101,31,250,31,76,31,38,31,55,31,164,31,197,31,179,31,219,31,108,31,253,31,244,31,125,31,144,31,62,31,242,31,156,31,146,31,254,31,210,31,123,31,126,31,160,31,205,31,37,31,106,31,206,31,88,31,88,30,18,31,60,31,185,31,185,30,14,31,14,30,21,31,172,31,40,31,40,30,56,31,56,30,232,31,114,31,186,31,2,31,158,31,200,31,210,31,14,31,56,31,9,31,17,31,15,31,15,30,129,31,76,31,190,31,131,31,138,31,116,31,76,31,76,30,76,29,89,31,199,31,199,30,42,31,42,30,158,31,246,31,19,31,174,31,82,31,184,31,224,31,102,31,102,30,65,31,164,31,132,31,241,31,70,31,10,31,80,31,42,31,145,31,229,31,229,30,210,31,140,31,36,31,10,31,187,31,124,31,124,30,246,31,50,31,150,31,150,30,83,31,83,30,83,29,174,31,161,31,134,31,134,30,9,31,9,30,247,31,247,31,226,31,64,31,53,31,38,31,15,31,116,31,12,31,244,31,19,31,19,30,121,31,224,31,224,30,14,31,17,31,29,31,29,30,77,31,77,30,21,31,21,30,151,31,96,31,131,31,94,31,21,31,150,31,157,31,247,31,208,31,190,31,227,31,141,31,219,31,151,31,180,31,222,31,222,30,222,29,197,31,8,31,137,31,254,31,107,31,240,31,240,30,131,31,172,31,62,31,29,31,56,31,57,31,57,30,34,31,215,31,29,31,187,31,172,31,249,31,207,31,201,31,119,31,14,31,118,31,118,30,107,31,248,31,150,31,236,31,236,30,236,29,236,28,236,27,128,31,128,30,207,31,48,31,233,31,109,31,109,30,239,31,215,31,45,31,19,31,199,31,125,31,10,31,10,30,106,31,102,31,102,30,237,31,72,31,5,31,194,31,111,31,111,30,176,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
