-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_655 is
end project_tb_655;

architecture project_tb_arch_655 of project_tb_655 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 816;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (229,0,41,0,246,0,24,0,91,0,49,0,0,0,126,0,31,0,146,0,0,0,212,0,0,0,0,0,87,0,130,0,189,0,122,0,0,0,0,0,174,0,194,0,13,0,96,0,194,0,147,0,28,0,226,0,217,0,139,0,187,0,70,0,249,0,220,0,242,0,143,0,93,0,211,0,0,0,37,0,246,0,194,0,0,0,80,0,76,0,254,0,0,0,203,0,106,0,182,0,150,0,7,0,96,0,236,0,138,0,37,0,0,0,149,0,230,0,207,0,206,0,37,0,44,0,0,0,0,0,234,0,233,0,94,0,121,0,54,0,145,0,134,0,0,0,221,0,204,0,194,0,247,0,130,0,113,0,14,0,0,0,0,0,0,0,93,0,0,0,42,0,205,0,84,0,58,0,130,0,86,0,0,0,47,0,0,0,0,0,201,0,0,0,119,0,251,0,119,0,168,0,0,0,14,0,0,0,182,0,248,0,204,0,39,0,138,0,0,0,168,0,233,0,172,0,126,0,162,0,210,0,99,0,0,0,102,0,150,0,175,0,3,0,109,0,88,0,78,0,0,0,0,0,250,0,0,0,241,0,204,0,176,0,22,0,243,0,0,0,49,0,46,0,59,0,203,0,52,0,0,0,161,0,17,0,80,0,0,0,175,0,134,0,130,0,26,0,0,0,20,0,199,0,75,0,75,0,38,0,218,0,243,0,245,0,65,0,0,0,0,0,234,0,0,0,68,0,183,0,207,0,222,0,171,0,178,0,221,0,34,0,91,0,24,0,0,0,0,0,209,0,3,0,97,0,245,0,228,0,6,0,0,0,239,0,19,0,107,0,64,0,240,0,142,0,139,0,0,0,177,0,199,0,37,0,154,0,231,0,0,0,0,0,236,0,155,0,0,0,96,0,183,0,0,0,0,0,139,0,14,0,137,0,215,0,45,0,88,0,0,0,149,0,139,0,143,0,73,0,245,0,127,0,0,0,0,0,222,0,127,0,129,0,0,0,92,0,0,0,150,0,37,0,185,0,0,0,208,0,196,0,124,0,0,0,0,0,69,0,243,0,178,0,34,0,143,0,225,0,173,0,110,0,203,0,233,0,70,0,0,0,191,0,199,0,228,0,239,0,55,0,156,0,188,0,0,0,108,0,101,0,149,0,240,0,141,0,83,0,30,0,0,0,188,0,138,0,2,0,130,0,0,0,53,0,0,0,0,0,57,0,225,0,116,0,0,0,103,0,0,0,151,0,241,0,104,0,0,0,244,0,169,0,0,0,211,0,132,0,0,0,252,0,0,0,168,0,188,0,188,0,147,0,118,0,92,0,58,0,109,0,0,0,10,0,200,0,211,0,89,0,92,0,0,0,48,0,127,0,0,0,53,0,205,0,55,0,0,0,130,0,70,0,207,0,0,0,229,0,144,0,70,0,0,0,157,0,199,0,241,0,174,0,0,0,161,0,69,0,0,0,224,0,73,0,0,0,0,0,198,0,32,0,145,0,0,0,136,0,246,0,88,0,0,0,199,0,0,0,79,0,82,0,218,0,92,0,41,0,0,0,168,0,16,0,0,0,45,0,27,0,54,0,0,0,0,0,0,0,123,0,207,0,152,0,0,0,11,0,225,0,225,0,189,0,246,0,66,0,75,0,0,0,50,0,89,0,96,0,57,0,104,0,216,0,220,0,171,0,59,0,0,0,233,0,0,0,0,0,0,0,0,0,213,0,209,0,255,0,169,0,64,0,0,0,167,0,211,0,18,0,153,0,0,0,52,0,196,0,68,0,175,0,155,0,206,0,0,0,0,0,0,0,215,0,169,0,255,0,0,0,0,0,188,0,152,0,0,0,247,0,48,0,132,0,0,0,103,0,158,0,117,0,170,0,152,0,0,0,36,0,0,0,230,0,0,0,191,0,25,0,120,0,0,0,151,0,168,0,146,0,0,0,52,0,139,0,101,0,190,0,197,0,0,0,6,0,241,0,81,0,213,0,27,0,84,0,23,0,0,0,143,0,0,0,54,0,40,0,149,0,98,0,0,0,0,0,114,0,207,0,0,0,70,0,222,0,0,0,0,0,0,0,189,0,179,0,17,0,146,0,0,0,156,0,122,0,129,0,67,0,138,0,230,0,170,0,245,0,239,0,134,0,172,0,61,0,139,0,0,0,136,0,78,0,103,0,57,0,172,0,152,0,0,0,91,0,58,0,33,0,255,0,0,0,78,0,216,0,51,0,173,0,30,0,45,0,148,0,0,0,47,0,148,0,22,0,88,0,172,0,189,0,165,0,201,0,32,0,238,0,164,0,152,0,88,0,105,0,65,0,76,0,246,0,146,0,38,0,65,0,97,0,166,0,0,0,190,0,136,0,137,0,44,0,16,0,148,0,247,0,0,0,0,0,247,0,161,0,0,0,124,0,16,0,95,0,125,0,66,0,245,0,169,0,177,0,0,0,173,0,216,0,81,0,54,0,2,0,0,0,114,0,246,0,98,0,225,0,14,0,121,0,90,0,254,0,138,0,74,0,82,0,0,0,6,0,186,0,55,0,0,0,210,0,93,0,244,0,195,0,57,0,124,0,182,0,82,0,5,0,187,0,133,0,202,0,94,0,115,0,123,0,83,0,0,0,0,0,230,0,232,0,173,0,104,0,165,0,190,0,163,0,0,0,54,0,232,0,56,0,36,0,16,0,1,0,95,0,91,0,106,0,32,0,254,0,203,0,0,0,53,0,191,0,0,0,154,0,59,0,82,0,56,0,40,0,0,0,230,0,0,0,150,0,0,0,134,0,89,0,0,0,108,0,223,0,136,0,0,0,227,0,0,0,192,0,147,0,0,0,0,0,166,0,0,0,0,0,30,0,121,0,191,0,64,0,85,0,97,0,56,0,36,0,107,0,90,0,133,0,227,0,52,0,190,0,238,0,28,0,80,0,76,0,145,0,44,0,0,0,157,0,214,0,154,0,166,0,140,0,53,0,0,0,17,0,0,0,0,0,247,0,16,0,51,0,52,0,0,0,177,0,230,0,0,0,209,0,186,0,80,0,27,0,0,0,233,0,217,0,188,0,45,0,0,0,144,0,131,0,20,0,9,0,104,0,10,0,228,0,86,0,78,0,0,0,243,0,40,0,12,0,228,0,16,0,236,0,238,0,0,0,0,0,146,0,237,0,197,0,199,0,97,0,215,0,0,0,240,0,232,0,254,0,30,0,137,0,109,0,254,0,0,0,0,0,0,0,0,0,234,0,109,0,15,0,0,0,209,0,27,0,0,0,0,0,27,0,114,0,192,0,0,0,120,0,6,0,164,0,4,0,159,0,0,0,189,0,0,0,71,0,13,0,0,0,0,0,186,0,0,0,225,0,171,0,175,0,122,0,0,0,82,0,63,0,203,0,101,0,77,0,32,0,83,0,141,0,0,0,184,0,28,0,0,0,2,0,103,0,42,0,242,0,149,0,116,0,0,0,0,0,181,0,186,0,47,0,130,0,0,0,129,0,111,0,24,0,0,0,143,0,0,0,135,0,94,0,0,0,209,0,0,0,74,0,7,0,0,0,0,0,233,0,166,0,188,0,215,0,159,0,41,0,106,0,62,0,135,0,187,0,32,0,136,0,47,0,0,0,82,0,225,0,0,0,40,0,46,0,25,0,0,0,57,0,76,0,0,0);
signal scenario_full  : scenario_type := (229,31,41,31,246,31,24,31,91,31,49,31,49,30,126,31,31,31,146,31,146,30,212,31,212,30,212,29,87,31,130,31,189,31,122,31,122,30,122,29,174,31,194,31,13,31,96,31,194,31,147,31,28,31,226,31,217,31,139,31,187,31,70,31,249,31,220,31,242,31,143,31,93,31,211,31,211,30,37,31,246,31,194,31,194,30,80,31,76,31,254,31,254,30,203,31,106,31,182,31,150,31,7,31,96,31,236,31,138,31,37,31,37,30,149,31,230,31,207,31,206,31,37,31,44,31,44,30,44,29,234,31,233,31,94,31,121,31,54,31,145,31,134,31,134,30,221,31,204,31,194,31,247,31,130,31,113,31,14,31,14,30,14,29,14,28,93,31,93,30,42,31,205,31,84,31,58,31,130,31,86,31,86,30,47,31,47,30,47,29,201,31,201,30,119,31,251,31,119,31,168,31,168,30,14,31,14,30,182,31,248,31,204,31,39,31,138,31,138,30,168,31,233,31,172,31,126,31,162,31,210,31,99,31,99,30,102,31,150,31,175,31,3,31,109,31,88,31,78,31,78,30,78,29,250,31,250,30,241,31,204,31,176,31,22,31,243,31,243,30,49,31,46,31,59,31,203,31,52,31,52,30,161,31,17,31,80,31,80,30,175,31,134,31,130,31,26,31,26,30,20,31,199,31,75,31,75,31,38,31,218,31,243,31,245,31,65,31,65,30,65,29,234,31,234,30,68,31,183,31,207,31,222,31,171,31,178,31,221,31,34,31,91,31,24,31,24,30,24,29,209,31,3,31,97,31,245,31,228,31,6,31,6,30,239,31,19,31,107,31,64,31,240,31,142,31,139,31,139,30,177,31,199,31,37,31,154,31,231,31,231,30,231,29,236,31,155,31,155,30,96,31,183,31,183,30,183,29,139,31,14,31,137,31,215,31,45,31,88,31,88,30,149,31,139,31,143,31,73,31,245,31,127,31,127,30,127,29,222,31,127,31,129,31,129,30,92,31,92,30,150,31,37,31,185,31,185,30,208,31,196,31,124,31,124,30,124,29,69,31,243,31,178,31,34,31,143,31,225,31,173,31,110,31,203,31,233,31,70,31,70,30,191,31,199,31,228,31,239,31,55,31,156,31,188,31,188,30,108,31,101,31,149,31,240,31,141,31,83,31,30,31,30,30,188,31,138,31,2,31,130,31,130,30,53,31,53,30,53,29,57,31,225,31,116,31,116,30,103,31,103,30,151,31,241,31,104,31,104,30,244,31,169,31,169,30,211,31,132,31,132,30,252,31,252,30,168,31,188,31,188,31,147,31,118,31,92,31,58,31,109,31,109,30,10,31,200,31,211,31,89,31,92,31,92,30,48,31,127,31,127,30,53,31,205,31,55,31,55,30,130,31,70,31,207,31,207,30,229,31,144,31,70,31,70,30,157,31,199,31,241,31,174,31,174,30,161,31,69,31,69,30,224,31,73,31,73,30,73,29,198,31,32,31,145,31,145,30,136,31,246,31,88,31,88,30,199,31,199,30,79,31,82,31,218,31,92,31,41,31,41,30,168,31,16,31,16,30,45,31,27,31,54,31,54,30,54,29,54,28,123,31,207,31,152,31,152,30,11,31,225,31,225,31,189,31,246,31,66,31,75,31,75,30,50,31,89,31,96,31,57,31,104,31,216,31,220,31,171,31,59,31,59,30,233,31,233,30,233,29,233,28,233,27,213,31,209,31,255,31,169,31,64,31,64,30,167,31,211,31,18,31,153,31,153,30,52,31,196,31,68,31,175,31,155,31,206,31,206,30,206,29,206,28,215,31,169,31,255,31,255,30,255,29,188,31,152,31,152,30,247,31,48,31,132,31,132,30,103,31,158,31,117,31,170,31,152,31,152,30,36,31,36,30,230,31,230,30,191,31,25,31,120,31,120,30,151,31,168,31,146,31,146,30,52,31,139,31,101,31,190,31,197,31,197,30,6,31,241,31,81,31,213,31,27,31,84,31,23,31,23,30,143,31,143,30,54,31,40,31,149,31,98,31,98,30,98,29,114,31,207,31,207,30,70,31,222,31,222,30,222,29,222,28,189,31,179,31,17,31,146,31,146,30,156,31,122,31,129,31,67,31,138,31,230,31,170,31,245,31,239,31,134,31,172,31,61,31,139,31,139,30,136,31,78,31,103,31,57,31,172,31,152,31,152,30,91,31,58,31,33,31,255,31,255,30,78,31,216,31,51,31,173,31,30,31,45,31,148,31,148,30,47,31,148,31,22,31,88,31,172,31,189,31,165,31,201,31,32,31,238,31,164,31,152,31,88,31,105,31,65,31,76,31,246,31,146,31,38,31,65,31,97,31,166,31,166,30,190,31,136,31,137,31,44,31,16,31,148,31,247,31,247,30,247,29,247,31,161,31,161,30,124,31,16,31,95,31,125,31,66,31,245,31,169,31,177,31,177,30,173,31,216,31,81,31,54,31,2,31,2,30,114,31,246,31,98,31,225,31,14,31,121,31,90,31,254,31,138,31,74,31,82,31,82,30,6,31,186,31,55,31,55,30,210,31,93,31,244,31,195,31,57,31,124,31,182,31,82,31,5,31,187,31,133,31,202,31,94,31,115,31,123,31,83,31,83,30,83,29,230,31,232,31,173,31,104,31,165,31,190,31,163,31,163,30,54,31,232,31,56,31,36,31,16,31,1,31,95,31,91,31,106,31,32,31,254,31,203,31,203,30,53,31,191,31,191,30,154,31,59,31,82,31,56,31,40,31,40,30,230,31,230,30,150,31,150,30,134,31,89,31,89,30,108,31,223,31,136,31,136,30,227,31,227,30,192,31,147,31,147,30,147,29,166,31,166,30,166,29,30,31,121,31,191,31,64,31,85,31,97,31,56,31,36,31,107,31,90,31,133,31,227,31,52,31,190,31,238,31,28,31,80,31,76,31,145,31,44,31,44,30,157,31,214,31,154,31,166,31,140,31,53,31,53,30,17,31,17,30,17,29,247,31,16,31,51,31,52,31,52,30,177,31,230,31,230,30,209,31,186,31,80,31,27,31,27,30,233,31,217,31,188,31,45,31,45,30,144,31,131,31,20,31,9,31,104,31,10,31,228,31,86,31,78,31,78,30,243,31,40,31,12,31,228,31,16,31,236,31,238,31,238,30,238,29,146,31,237,31,197,31,199,31,97,31,215,31,215,30,240,31,232,31,254,31,30,31,137,31,109,31,254,31,254,30,254,29,254,28,254,27,234,31,109,31,15,31,15,30,209,31,27,31,27,30,27,29,27,31,114,31,192,31,192,30,120,31,6,31,164,31,4,31,159,31,159,30,189,31,189,30,71,31,13,31,13,30,13,29,186,31,186,30,225,31,171,31,175,31,122,31,122,30,82,31,63,31,203,31,101,31,77,31,32,31,83,31,141,31,141,30,184,31,28,31,28,30,2,31,103,31,42,31,242,31,149,31,116,31,116,30,116,29,181,31,186,31,47,31,130,31,130,30,129,31,111,31,24,31,24,30,143,31,143,30,135,31,94,31,94,30,209,31,209,30,74,31,7,31,7,30,7,29,233,31,166,31,188,31,215,31,159,31,41,31,106,31,62,31,135,31,187,31,32,31,136,31,47,31,47,30,82,31,225,31,225,30,40,31,46,31,25,31,25,30,57,31,76,31,76,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
