-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 244;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (224,0,111,0,0,0,180,0,197,0,225,0,200,0,155,0,130,0,225,0,0,0,0,0,0,0,74,0,238,0,48,0,170,0,0,0,76,0,148,0,0,0,167,0,10,0,0,0,150,0,7,0,222,0,0,0,0,0,9,0,21,0,0,0,96,0,232,0,17,0,131,0,246,0,201,0,182,0,0,0,7,0,248,0,25,0,0,0,208,0,213,0,64,0,171,0,99,0,64,0,171,0,210,0,40,0,0,0,139,0,0,0,138,0,213,0,64,0,134,0,78,0,136,0,42,0,0,0,163,0,0,0,0,0,0,0,33,0,210,0,77,0,27,0,104,0,0,0,198,0,61,0,159,0,0,0,214,0,208,0,0,0,93,0,0,0,91,0,56,0,0,0,219,0,135,0,155,0,0,0,178,0,211,0,64,0,183,0,132,0,138,0,168,0,183,0,0,0,0,0,201,0,0,0,231,0,0,0,178,0,0,0,60,0,134,0,143,0,114,0,233,0,225,0,15,0,153,0,1,0,0,0,125,0,0,0,0,0,59,0,22,0,175,0,144,0,26,0,230,0,16,0,108,0,0,0,9,0,21,0,208,0,11,0,67,0,0,0,0,0,195,0,0,0,62,0,48,0,0,0,218,0,0,0,23,0,147,0,135,0,0,0,58,0,64,0,236,0,172,0,185,0,125,0,126,0,134,0,0,0,125,0,0,0,153,0,195,0,200,0,125,0,87,0,0,0,54,0,0,0,232,0,213,0,230,0,219,0,55,0,123,0,163,0,0,0,210,0,0,0,99,0,179,0,0,0,250,0,0,0,178,0,214,0,163,0,194,0,0,0,0,0,0,0,154,0,0,0,13,0,0,0,146,0,77,0,0,0,0,0,239,0,204,0,196,0,0,0,0,0,135,0,189,0,0,0,79,0,0,0,0,0,8,0,216,0,255,0,0,0,223,0,190,0,255,0,124,0,0,0,0,0,226,0,155,0,75,0,0,0,122,0,60,0,0,0,209,0,251,0,0,0,105,0,127,0,0,0,68,0,107,0,9,0,173,0,226,0,0,0,0,0,0,0,82,0,125,0,228,0,237,0,252,0,143,0,122,0);
signal scenario_full  : scenario_type := (224,31,111,31,111,30,180,31,197,31,225,31,200,31,155,31,130,31,225,31,225,30,225,29,225,28,74,31,238,31,48,31,170,31,170,30,76,31,148,31,148,30,167,31,10,31,10,30,150,31,7,31,222,31,222,30,222,29,9,31,21,31,21,30,96,31,232,31,17,31,131,31,246,31,201,31,182,31,182,30,7,31,248,31,25,31,25,30,208,31,213,31,64,31,171,31,99,31,64,31,171,31,210,31,40,31,40,30,139,31,139,30,138,31,213,31,64,31,134,31,78,31,136,31,42,31,42,30,163,31,163,30,163,29,163,28,33,31,210,31,77,31,27,31,104,31,104,30,198,31,61,31,159,31,159,30,214,31,208,31,208,30,93,31,93,30,91,31,56,31,56,30,219,31,135,31,155,31,155,30,178,31,211,31,64,31,183,31,132,31,138,31,168,31,183,31,183,30,183,29,201,31,201,30,231,31,231,30,178,31,178,30,60,31,134,31,143,31,114,31,233,31,225,31,15,31,153,31,1,31,1,30,125,31,125,30,125,29,59,31,22,31,175,31,144,31,26,31,230,31,16,31,108,31,108,30,9,31,21,31,208,31,11,31,67,31,67,30,67,29,195,31,195,30,62,31,48,31,48,30,218,31,218,30,23,31,147,31,135,31,135,30,58,31,64,31,236,31,172,31,185,31,125,31,126,31,134,31,134,30,125,31,125,30,153,31,195,31,200,31,125,31,87,31,87,30,54,31,54,30,232,31,213,31,230,31,219,31,55,31,123,31,163,31,163,30,210,31,210,30,99,31,179,31,179,30,250,31,250,30,178,31,214,31,163,31,194,31,194,30,194,29,194,28,154,31,154,30,13,31,13,30,146,31,77,31,77,30,77,29,239,31,204,31,196,31,196,30,196,29,135,31,189,31,189,30,79,31,79,30,79,29,8,31,216,31,255,31,255,30,223,31,190,31,255,31,124,31,124,30,124,29,226,31,155,31,75,31,75,30,122,31,60,31,60,30,209,31,251,31,251,30,105,31,127,31,127,30,68,31,107,31,9,31,173,31,226,31,226,30,226,29,226,28,82,31,125,31,228,31,237,31,252,31,143,31,122,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
