-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 194;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (171,0,72,0,237,0,210,0,0,0,3,0,0,0,230,0,67,0,131,0,158,0,192,0,233,0,90,0,35,0,153,0,66,0,2,0,83,0,125,0,0,0,169,0,52,0,200,0,33,0,159,0,181,0,227,0,0,0,0,0,127,0,99,0,125,0,47,0,0,0,0,0,235,0,0,0,140,0,217,0,197,0,127,0,0,0,0,0,58,0,195,0,78,0,0,0,50,0,223,0,36,0,141,0,109,0,233,0,7,0,183,0,135,0,145,0,47,0,108,0,129,0,93,0,85,0,80,0,0,0,0,0,64,0,0,0,62,0,247,0,147,0,154,0,47,0,198,0,184,0,0,0,0,0,0,0,50,0,134,0,8,0,50,0,208,0,49,0,48,0,235,0,127,0,0,0,0,0,90,0,158,0,157,0,175,0,136,0,213,0,42,0,120,0,58,0,156,0,106,0,32,0,175,0,208,0,0,0,93,0,250,0,243,0,198,0,168,0,60,0,109,0,26,0,0,0,0,0,0,0,225,0,0,0,176,0,11,0,153,0,198,0,133,0,0,0,0,0,0,0,253,0,116,0,85,0,188,0,41,0,37,0,252,0,172,0,180,0,76,0,0,0,254,0,0,0,0,0,0,0,78,0,153,0,0,0,26,0,0,0,0,0,121,0,145,0,0,0,3,0,70,0,162,0,0,0,90,0,0,0,0,0,81,0,213,0,88,0,200,0,133,0,74,0,43,0,0,0,105,0,0,0,170,0,222,0,78,0,53,0,121,0,112,0,109,0,222,0,89,0,65,0,128,0,0,0,140,0,121,0,0,0,96,0,244,0,207,0,151,0,37,0,172,0,114,0,0,0,82,0,32,0,101,0,88,0,84,0);
signal scenario_full  : scenario_type := (171,31,72,31,237,31,210,31,210,30,3,31,3,30,230,31,67,31,131,31,158,31,192,31,233,31,90,31,35,31,153,31,66,31,2,31,83,31,125,31,125,30,169,31,52,31,200,31,33,31,159,31,181,31,227,31,227,30,227,29,127,31,99,31,125,31,47,31,47,30,47,29,235,31,235,30,140,31,217,31,197,31,127,31,127,30,127,29,58,31,195,31,78,31,78,30,50,31,223,31,36,31,141,31,109,31,233,31,7,31,183,31,135,31,145,31,47,31,108,31,129,31,93,31,85,31,80,31,80,30,80,29,64,31,64,30,62,31,247,31,147,31,154,31,47,31,198,31,184,31,184,30,184,29,184,28,50,31,134,31,8,31,50,31,208,31,49,31,48,31,235,31,127,31,127,30,127,29,90,31,158,31,157,31,175,31,136,31,213,31,42,31,120,31,58,31,156,31,106,31,32,31,175,31,208,31,208,30,93,31,250,31,243,31,198,31,168,31,60,31,109,31,26,31,26,30,26,29,26,28,225,31,225,30,176,31,11,31,153,31,198,31,133,31,133,30,133,29,133,28,253,31,116,31,85,31,188,31,41,31,37,31,252,31,172,31,180,31,76,31,76,30,254,31,254,30,254,29,254,28,78,31,153,31,153,30,26,31,26,30,26,29,121,31,145,31,145,30,3,31,70,31,162,31,162,30,90,31,90,30,90,29,81,31,213,31,88,31,200,31,133,31,74,31,43,31,43,30,105,31,105,30,170,31,222,31,78,31,53,31,121,31,112,31,109,31,222,31,89,31,65,31,128,31,128,30,140,31,121,31,121,30,96,31,244,31,207,31,151,31,37,31,172,31,114,31,114,30,82,31,32,31,101,31,88,31,84,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
