-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 482;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,166,0,0,0,114,0,210,0,0,0,0,0,218,0,0,0,0,0,110,0,0,0,0,0,30,0,74,0,0,0,0,0,154,0,71,0,0,0,113,0,133,0,188,0,0,0,0,0,0,0,142,0,0,0,39,0,132,0,237,0,66,0,86,0,73,0,45,0,112,0,140,0,0,0,73,0,227,0,0,0,239,0,122,0,153,0,15,0,80,0,122,0,179,0,71,0,58,0,0,0,153,0,139,0,151,0,0,0,49,0,165,0,141,0,0,0,9,0,246,0,0,0,45,0,186,0,77,0,0,0,198,0,163,0,33,0,85,0,211,0,28,0,6,0,11,0,0,0,79,0,236,0,0,0,25,0,98,0,246,0,121,0,190,0,59,0,207,0,138,0,163,0,68,0,202,0,249,0,102,0,220,0,12,0,72,0,198,0,73,0,0,0,0,0,105,0,9,0,252,0,21,0,0,0,0,0,213,0,155,0,66,0,161,0,252,0,0,0,178,0,239,0,108,0,45,0,247,0,48,0,118,0,123,0,68,0,2,0,2,0,0,0,24,0,19,0,84,0,7,0,0,0,137,0,20,0,0,0,64,0,102,0,253,0,250,0,0,0,47,0,82,0,69,0,47,0,0,0,134,0,227,0,89,0,86,0,130,0,0,0,127,0,130,0,127,0,47,0,68,0,0,0,156,0,0,0,0,0,54,0,0,0,150,0,0,0,85,0,30,0,0,0,4,0,69,0,122,0,184,0,249,0,113,0,0,0,0,0,220,0,57,0,57,0,13,0,16,0,121,0,59,0,82,0,86,0,102,0,33,0,252,0,212,0,0,0,245,0,93,0,0,0,244,0,195,0,60,0,165,0,116,0,37,0,0,0,0,0,203,0,24,0,55,0,39,0,134,0,246,0,96,0,244,0,21,0,48,0,195,0,0,0,217,0,105,0,59,0,77,0,24,0,224,0,50,0,0,0,118,0,139,0,0,0,45,0,182,0,208,0,166,0,148,0,164,0,223,0,222,0,24,0,0,0,0,0,217,0,241,0,110,0,42,0,133,0,152,0,9,0,98,0,118,0,97,0,90,0,72,0,92,0,149,0,146,0,0,0,99,0,59,0,0,0,0,0,30,0,76,0,0,0,73,0,146,0,143,0,0,0,29,0,243,0,168,0,0,0,131,0,115,0,0,0,147,0,12,0,157,0,189,0,221,0,93,0,161,0,100,0,0,0,179,0,0,0,0,0,202,0,97,0,166,0,164,0,194,0,0,0,32,0,101,0,0,0,189,0,218,0,82,0,13,0,120,0,11,0,189,0,247,0,239,0,41,0,122,0,192,0,16,0,47,0,108,0,82,0,130,0,252,0,0,0,54,0,86,0,162,0,3,0,58,0,223,0,80,0,155,0,194,0,29,0,0,0,248,0,82,0,73,0,49,0,94,0,0,0,0,0,64,0,21,0,120,0,0,0,123,0,1,0,0,0,128,0,186,0,0,0,0,0,206,0,178,0,142,0,38,0,122,0,90,0,102,0,0,0,114,0,122,0,45,0,67,0,40,0,30,0,0,0,29,0,132,0,241,0,135,0,173,0,0,0,18,0,82,0,38,0,95,0,91,0,29,0,186,0,186,0,0,0,224,0,225,0,112,0,223,0,173,0,219,0,247,0,190,0,34,0,24,0,205,0,218,0,51,0,99,0,0,0,0,0,45,0,32,0,169,0,166,0,217,0,10,0,76,0,24,0,121,0,44,0,0,0,168,0,221,0,244,0,216,0,73,0,0,0,77,0,73,0,204,0,114,0,221,0,185,0,102,0,0,0,221,0,45,0,121,0,0,0,4,0,9,0,111,0,128,0,217,0,60,0,57,0,74,0,92,0,15,0,0,0,198,0,31,0,46,0,0,0,140,0,112,0,141,0,101,0,27,0,250,0,227,0,233,0,239,0,238,0,198,0,0,0,165,0,225,0,248,0,81,0,126,0,186,0,76,0,55,0,203,0,149,0,216,0,90,0,163,0,220,0,237,0,185,0,77,0,158,0,85,0,177,0,167,0,190,0,223,0,129,0,167,0,13,0,160,0,135,0,52,0,64,0,0,0,211,0,63,0,223,0,48,0,0,0,0,0,79,0,82,0,96,0,235,0,109,0,227,0,137,0,158,0,107,0,108,0,48,0);
signal scenario_full  : scenario_type := (0,0,166,31,166,30,114,31,210,31,210,30,210,29,218,31,218,30,218,29,110,31,110,30,110,29,30,31,74,31,74,30,74,29,154,31,71,31,71,30,113,31,133,31,188,31,188,30,188,29,188,28,142,31,142,30,39,31,132,31,237,31,66,31,86,31,73,31,45,31,112,31,140,31,140,30,73,31,227,31,227,30,239,31,122,31,153,31,15,31,80,31,122,31,179,31,71,31,58,31,58,30,153,31,139,31,151,31,151,30,49,31,165,31,141,31,141,30,9,31,246,31,246,30,45,31,186,31,77,31,77,30,198,31,163,31,33,31,85,31,211,31,28,31,6,31,11,31,11,30,79,31,236,31,236,30,25,31,98,31,246,31,121,31,190,31,59,31,207,31,138,31,163,31,68,31,202,31,249,31,102,31,220,31,12,31,72,31,198,31,73,31,73,30,73,29,105,31,9,31,252,31,21,31,21,30,21,29,213,31,155,31,66,31,161,31,252,31,252,30,178,31,239,31,108,31,45,31,247,31,48,31,118,31,123,31,68,31,2,31,2,31,2,30,24,31,19,31,84,31,7,31,7,30,137,31,20,31,20,30,64,31,102,31,253,31,250,31,250,30,47,31,82,31,69,31,47,31,47,30,134,31,227,31,89,31,86,31,130,31,130,30,127,31,130,31,127,31,47,31,68,31,68,30,156,31,156,30,156,29,54,31,54,30,150,31,150,30,85,31,30,31,30,30,4,31,69,31,122,31,184,31,249,31,113,31,113,30,113,29,220,31,57,31,57,31,13,31,16,31,121,31,59,31,82,31,86,31,102,31,33,31,252,31,212,31,212,30,245,31,93,31,93,30,244,31,195,31,60,31,165,31,116,31,37,31,37,30,37,29,203,31,24,31,55,31,39,31,134,31,246,31,96,31,244,31,21,31,48,31,195,31,195,30,217,31,105,31,59,31,77,31,24,31,224,31,50,31,50,30,118,31,139,31,139,30,45,31,182,31,208,31,166,31,148,31,164,31,223,31,222,31,24,31,24,30,24,29,217,31,241,31,110,31,42,31,133,31,152,31,9,31,98,31,118,31,97,31,90,31,72,31,92,31,149,31,146,31,146,30,99,31,59,31,59,30,59,29,30,31,76,31,76,30,73,31,146,31,143,31,143,30,29,31,243,31,168,31,168,30,131,31,115,31,115,30,147,31,12,31,157,31,189,31,221,31,93,31,161,31,100,31,100,30,179,31,179,30,179,29,202,31,97,31,166,31,164,31,194,31,194,30,32,31,101,31,101,30,189,31,218,31,82,31,13,31,120,31,11,31,189,31,247,31,239,31,41,31,122,31,192,31,16,31,47,31,108,31,82,31,130,31,252,31,252,30,54,31,86,31,162,31,3,31,58,31,223,31,80,31,155,31,194,31,29,31,29,30,248,31,82,31,73,31,49,31,94,31,94,30,94,29,64,31,21,31,120,31,120,30,123,31,1,31,1,30,128,31,186,31,186,30,186,29,206,31,178,31,142,31,38,31,122,31,90,31,102,31,102,30,114,31,122,31,45,31,67,31,40,31,30,31,30,30,29,31,132,31,241,31,135,31,173,31,173,30,18,31,82,31,38,31,95,31,91,31,29,31,186,31,186,31,186,30,224,31,225,31,112,31,223,31,173,31,219,31,247,31,190,31,34,31,24,31,205,31,218,31,51,31,99,31,99,30,99,29,45,31,32,31,169,31,166,31,217,31,10,31,76,31,24,31,121,31,44,31,44,30,168,31,221,31,244,31,216,31,73,31,73,30,77,31,73,31,204,31,114,31,221,31,185,31,102,31,102,30,221,31,45,31,121,31,121,30,4,31,9,31,111,31,128,31,217,31,60,31,57,31,74,31,92,31,15,31,15,30,198,31,31,31,46,31,46,30,140,31,112,31,141,31,101,31,27,31,250,31,227,31,233,31,239,31,238,31,198,31,198,30,165,31,225,31,248,31,81,31,126,31,186,31,76,31,55,31,203,31,149,31,216,31,90,31,163,31,220,31,237,31,185,31,77,31,158,31,85,31,177,31,167,31,190,31,223,31,129,31,167,31,13,31,160,31,135,31,52,31,64,31,64,30,211,31,63,31,223,31,48,31,48,30,48,29,79,31,82,31,96,31,235,31,109,31,227,31,137,31,158,31,107,31,108,31,48,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
