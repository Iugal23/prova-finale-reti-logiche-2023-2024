-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_821 is
end project_tb_821;

architecture project_tb_arch_821 of project_tb_821 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 463;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (98,0,182,0,194,0,0,0,62,0,255,0,85,0,0,0,239,0,0,0,0,0,150,0,248,0,194,0,0,0,0,0,207,0,0,0,138,0,119,0,194,0,0,0,241,0,102,0,123,0,188,0,159,0,60,0,59,0,118,0,85,0,95,0,0,0,105,0,138,0,240,0,28,0,71,0,248,0,0,0,0,0,244,0,126,0,0,0,220,0,225,0,0,0,63,0,117,0,18,0,109,0,82,0,165,0,200,0,16,0,248,0,177,0,168,0,157,0,0,0,215,0,50,0,221,0,236,0,220,0,238,0,80,0,134,0,117,0,178,0,144,0,0,0,42,0,7,0,106,0,185,0,62,0,221,0,0,0,27,0,230,0,0,0,0,0,0,0,124,0,121,0,0,0,82,0,193,0,251,0,120,0,121,0,229,0,128,0,198,0,19,0,147,0,0,0,128,0,25,0,96,0,0,0,29,0,0,0,155,0,72,0,0,0,65,0,26,0,152,0,106,0,60,0,0,0,98,0,247,0,173,0,0,0,108,0,25,0,84,0,182,0,0,0,69,0,175,0,140,0,58,0,3,0,0,0,45,0,61,0,177,0,0,0,28,0,104,0,0,0,0,0,48,0,93,0,249,0,253,0,150,0,0,0,119,0,114,0,115,0,107,0,164,0,247,0,162,0,94,0,9,0,133,0,246,0,0,0,2,0,197,0,0,0,190,0,68,0,220,0,194,0,133,0,104,0,0,0,126,0,25,0,6,0,133,0,175,0,12,0,152,0,221,0,0,0,0,0,140,0,250,0,207,0,0,0,22,0,41,0,144,0,25,0,23,0,23,0,0,0,66,0,10,0,94,0,27,0,247,0,192,0,0,0,62,0,0,0,31,0,191,0,172,0,0,0,102,0,155,0,63,0,174,0,137,0,228,0,0,0,239,0,179,0,170,0,40,0,151,0,69,0,172,0,58,0,10,0,116,0,0,0,109,0,143,0,25,0,52,0,24,0,162,0,215,0,80,0,0,0,43,0,65,0,0,0,141,0,154,0,186,0,152,0,82,0,13,0,0,0,142,0,0,0,186,0,0,0,242,0,64,0,0,0,210,0,28,0,0,0,139,0,154,0,62,0,245,0,0,0,0,0,112,0,72,0,5,0,105,0,97,0,0,0,89,0,136,0,0,0,88,0,0,0,11,0,229,0,250,0,0,0,201,0,34,0,98,0,235,0,213,0,115,0,0,0,151,0,58,0,114,0,123,0,0,0,0,0,222,0,253,0,128,0,241,0,240,0,0,0,27,0,100,0,175,0,0,0,0,0,0,0,112,0,193,0,72,0,180,0,171,0,0,0,191,0,52,0,116,0,161,0,5,0,29,0,216,0,178,0,159,0,191,0,0,0,19,0,16,0,237,0,77,0,180,0,62,0,91,0,0,0,207,0,242,0,186,0,89,0,141,0,121,0,91,0,255,0,121,0,68,0,23,0,252,0,198,0,11,0,226,0,72,0,148,0,201,0,51,0,60,0,45,0,204,0,0,0,43,0,185,0,231,0,0,0,87,0,63,0,232,0,250,0,120,0,204,0,237,0,195,0,113,0,0,0,114,0,60,0,0,0,161,0,145,0,126,0,84,0,103,0,232,0,0,0,1,0,0,0,0,0,91,0,99,0,25,0,137,0,174,0,135,0,100,0,244,0,34,0,89,0,204,0,123,0,210,0,250,0,55,0,113,0,48,0,249,0,126,0,205,0,169,0,0,0,0,0,201,0,77,0,88,0,0,0,39,0,219,0,139,0,250,0,227,0,0,0,0,0,209,0,173,0,197,0,239,0,187,0,5,0,104,0,72,0,0,0,150,0,182,0,56,0,154,0,0,0,246,0,81,0,114,0,9,0,97,0,20,0,222,0,43,0,60,0,25,0,151,0,187,0,34,0,0,0,143,0,39,0,28,0,0,0,104,0,140,0,185,0,162,0,239,0,131,0,223,0,77,0,23,0,0,0,172,0,58,0,4,0,54,0,177,0,7,0,32,0,217,0,0,0,231,0,132,0,104,0,193,0,84,0,164,0,176,0,23,0,0,0,75,0,33,0,0,0);
signal scenario_full  : scenario_type := (98,31,182,31,194,31,194,30,62,31,255,31,85,31,85,30,239,31,239,30,239,29,150,31,248,31,194,31,194,30,194,29,207,31,207,30,138,31,119,31,194,31,194,30,241,31,102,31,123,31,188,31,159,31,60,31,59,31,118,31,85,31,95,31,95,30,105,31,138,31,240,31,28,31,71,31,248,31,248,30,248,29,244,31,126,31,126,30,220,31,225,31,225,30,63,31,117,31,18,31,109,31,82,31,165,31,200,31,16,31,248,31,177,31,168,31,157,31,157,30,215,31,50,31,221,31,236,31,220,31,238,31,80,31,134,31,117,31,178,31,144,31,144,30,42,31,7,31,106,31,185,31,62,31,221,31,221,30,27,31,230,31,230,30,230,29,230,28,124,31,121,31,121,30,82,31,193,31,251,31,120,31,121,31,229,31,128,31,198,31,19,31,147,31,147,30,128,31,25,31,96,31,96,30,29,31,29,30,155,31,72,31,72,30,65,31,26,31,152,31,106,31,60,31,60,30,98,31,247,31,173,31,173,30,108,31,25,31,84,31,182,31,182,30,69,31,175,31,140,31,58,31,3,31,3,30,45,31,61,31,177,31,177,30,28,31,104,31,104,30,104,29,48,31,93,31,249,31,253,31,150,31,150,30,119,31,114,31,115,31,107,31,164,31,247,31,162,31,94,31,9,31,133,31,246,31,246,30,2,31,197,31,197,30,190,31,68,31,220,31,194,31,133,31,104,31,104,30,126,31,25,31,6,31,133,31,175,31,12,31,152,31,221,31,221,30,221,29,140,31,250,31,207,31,207,30,22,31,41,31,144,31,25,31,23,31,23,31,23,30,66,31,10,31,94,31,27,31,247,31,192,31,192,30,62,31,62,30,31,31,191,31,172,31,172,30,102,31,155,31,63,31,174,31,137,31,228,31,228,30,239,31,179,31,170,31,40,31,151,31,69,31,172,31,58,31,10,31,116,31,116,30,109,31,143,31,25,31,52,31,24,31,162,31,215,31,80,31,80,30,43,31,65,31,65,30,141,31,154,31,186,31,152,31,82,31,13,31,13,30,142,31,142,30,186,31,186,30,242,31,64,31,64,30,210,31,28,31,28,30,139,31,154,31,62,31,245,31,245,30,245,29,112,31,72,31,5,31,105,31,97,31,97,30,89,31,136,31,136,30,88,31,88,30,11,31,229,31,250,31,250,30,201,31,34,31,98,31,235,31,213,31,115,31,115,30,151,31,58,31,114,31,123,31,123,30,123,29,222,31,253,31,128,31,241,31,240,31,240,30,27,31,100,31,175,31,175,30,175,29,175,28,112,31,193,31,72,31,180,31,171,31,171,30,191,31,52,31,116,31,161,31,5,31,29,31,216,31,178,31,159,31,191,31,191,30,19,31,16,31,237,31,77,31,180,31,62,31,91,31,91,30,207,31,242,31,186,31,89,31,141,31,121,31,91,31,255,31,121,31,68,31,23,31,252,31,198,31,11,31,226,31,72,31,148,31,201,31,51,31,60,31,45,31,204,31,204,30,43,31,185,31,231,31,231,30,87,31,63,31,232,31,250,31,120,31,204,31,237,31,195,31,113,31,113,30,114,31,60,31,60,30,161,31,145,31,126,31,84,31,103,31,232,31,232,30,1,31,1,30,1,29,91,31,99,31,25,31,137,31,174,31,135,31,100,31,244,31,34,31,89,31,204,31,123,31,210,31,250,31,55,31,113,31,48,31,249,31,126,31,205,31,169,31,169,30,169,29,201,31,77,31,88,31,88,30,39,31,219,31,139,31,250,31,227,31,227,30,227,29,209,31,173,31,197,31,239,31,187,31,5,31,104,31,72,31,72,30,150,31,182,31,56,31,154,31,154,30,246,31,81,31,114,31,9,31,97,31,20,31,222,31,43,31,60,31,25,31,151,31,187,31,34,31,34,30,143,31,39,31,28,31,28,30,104,31,140,31,185,31,162,31,239,31,131,31,223,31,77,31,23,31,23,30,172,31,58,31,4,31,54,31,177,31,7,31,32,31,217,31,217,30,231,31,132,31,104,31,193,31,84,31,164,31,176,31,23,31,23,30,75,31,33,31,33,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
