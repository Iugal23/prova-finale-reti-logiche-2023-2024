-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_16 is
end project_tb_16;

architecture project_tb_arch_16 of project_tb_16 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 772;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (3,0,167,0,0,0,31,0,80,0,89,0,0,0,50,0,221,0,36,0,0,0,0,0,0,0,178,0,161,0,159,0,237,0,139,0,0,0,216,0,62,0,4,0,129,0,0,0,0,0,83,0,174,0,0,0,221,0,46,0,0,0,0,0,94,0,58,0,184,0,22,0,25,0,121,0,165,0,232,0,180,0,25,0,36,0,211,0,69,0,82,0,120,0,234,0,94,0,197,0,0,0,153,0,115,0,170,0,132,0,94,0,145,0,255,0,71,0,0,0,224,0,0,0,252,0,92,0,243,0,133,0,78,0,191,0,0,0,211,0,128,0,0,0,0,0,96,0,156,0,29,0,225,0,0,0,0,0,63,0,0,0,0,0,8,0,180,0,190,0,5,0,159,0,211,0,83,0,251,0,0,0,168,0,0,0,154,0,71,0,153,0,125,0,200,0,0,0,188,0,62,0,118,0,183,0,184,0,87,0,0,0,88,0,0,0,169,0,0,0,157,0,183,0,134,0,27,0,34,0,97,0,75,0,142,0,162,0,186,0,216,0,126,0,191,0,127,0,143,0,0,0,70,0,92,0,0,0,26,0,239,0,191,0,121,0,125,0,0,0,113,0,195,0,14,0,0,0,249,0,0,0,67,0,199,0,0,0,71,0,34,0,149,0,210,0,209,0,116,0,24,0,0,0,0,0,66,0,192,0,59,0,236,0,225,0,57,0,189,0,9,0,134,0,105,0,178,0,164,0,47,0,165,0,215,0,26,0,179,0,36,0,0,0,137,0,65,0,243,0,0,0,223,0,0,0,0,0,142,0,202,0,0,0,78,0,47,0,80,0,114,0,29,0,141,0,251,0,226,0,0,0,129,0,113,0,5,0,179,0,180,0,103,0,165,0,58,0,0,0,82,0,107,0,29,0,63,0,108,0,69,0,205,0,243,0,137,0,0,0,181,0,233,0,0,0,0,0,46,0,98,0,0,0,228,0,26,0,0,0,244,0,219,0,15,0,255,0,175,0,26,0,112,0,240,0,63,0,147,0,143,0,0,0,144,0,249,0,36,0,0,0,200,0,53,0,17,0,47,0,144,0,143,0,42,0,0,0,53,0,121,0,190,0,230,0,30,0,251,0,249,0,30,0,217,0,0,0,90,0,224,0,0,0,0,0,30,0,130,0,0,0,46,0,69,0,247,0,175,0,136,0,1,0,176,0,150,0,83,0,170,0,8,0,202,0,11,0,142,0,246,0,34,0,135,0,75,0,0,0,2,0,107,0,6,0,0,0,0,0,209,0,232,0,142,0,223,0,0,0,61,0,175,0,31,0,0,0,191,0,4,0,175,0,40,0,214,0,178,0,53,0,122,0,78,0,227,0,0,0,69,0,233,0,148,0,0,0,117,0,174,0,175,0,181,0,168,0,12,0,108,0,0,0,97,0,0,0,80,0,44,0,44,0,150,0,0,0,175,0,183,0,0,0,80,0,0,0,0,0,200,0,6,0,156,0,100,0,0,0,95,0,172,0,0,0,116,0,166,0,233,0,253,0,187,0,62,0,204,0,213,0,0,0,47,0,209,0,126,0,232,0,74,0,71,0,166,0,0,0,251,0,142,0,219,0,0,0,140,0,148,0,178,0,0,0,180,0,177,0,191,0,114,0,233,0,224,0,0,0,255,0,143,0,98,0,143,0,144,0,116,0,221,0,40,0,199,0,169,0,126,0,121,0,240,0,210,0,100,0,105,0,66,0,214,0,205,0,140,0,0,0,133,0,24,0,199,0,106,0,232,0,101,0,92,0,9,0,84,0,128,0,152,0,225,0,45,0,219,0,185,0,231,0,75,0,200,0,160,0,0,0,208,0,168,0,202,0,95,0,246,0,55,0,223,0,18,0,142,0,0,0,227,0,175,0,225,0,6,0,66,0,201,0,127,0,225,0,21,0,58,0,66,0,34,0,40,0,0,0,197,0,0,0,205,0,157,0,193,0,0,0,132,0,0,0,232,0,99,0,85,0,25,0,0,0,233,0,0,0,107,0,184,0,106,0,60,0,0,0,0,0,214,0,152,0,177,0,49,0,60,0,0,0,0,0,0,0,115,0,87,0,207,0,126,0,26,0,14,0,65,0,0,0,64,0,202,0,144,0,118,0,7,0,148,0,45,0,0,0,68,0,37,0,89,0,128,0,19,0,238,0,4,0,132,0,38,0,0,0,1,0,0,0,26,0,211,0,78,0,176,0,107,0,203,0,205,0,0,0,0,0,205,0,191,0,150,0,122,0,0,0,13,0,238,0,0,0,89,0,21,0,254,0,19,0,0,0,0,0,170,0,0,0,138,0,118,0,183,0,0,0,40,0,191,0,0,0,123,0,109,0,239,0,154,0,88,0,56,0,135,0,86,0,248,0,94,0,140,0,0,0,153,0,159,0,0,0,159,0,247,0,0,0,0,0,164,0,0,0,155,0,24,0,105,0,123,0,6,0,110,0,97,0,205,0,108,0,195,0,82,0,7,0,0,0,199,0,0,0,156,0,134,0,0,0,123,0,106,0,167,0,255,0,184,0,7,0,97,0,0,0,88,0,0,0,204,0,248,0,0,0,0,0,148,0,241,0,239,0,127,0,114,0,77,0,0,0,176,0,171,0,0,0,183,0,152,0,224,0,156,0,190,0,0,0,0,0,159,0,90,0,192,0,207,0,51,0,38,0,40,0,192,0,169,0,82,0,213,0,231,0,90,0,0,0,143,0,108,0,0,0,0,0,69,0,33,0,65,0,59,0,204,0,0,0,36,0,0,0,0,0,131,0,0,0,0,0,206,0,192,0,111,0,233,0,0,0,23,0,0,0,118,0,64,0,0,0,0,0,0,0,189,0,134,0,89,0,204,0,92,0,0,0,107,0,141,0,5,0,0,0,15,0,142,0,0,0,246,0,0,0,0,0,0,0,38,0,221,0,133,0,0,0,255,0,160,0,0,0,0,0,100,0,139,0,192,0,177,0,99,0,29,0,236,0,216,0,0,0,158,0,228,0,49,0,194,0,226,0,123,0,126,0,53,0,70,0,88,0,94,0,158,0,115,0,194,0,83,0,0,0,61,0,98,0,170,0,81,0,0,0,0,0,178,0,0,0,230,0,227,0,64,0,205,0,17,0,189,0,228,0,238,0,35,0,86,0,147,0,27,0,76,0,87,0,231,0,227,0,98,0,0,0,0,0,85,0,247,0,73,0,44,0,159,0,74,0,217,0,244,0,134,0,19,0,128,0,86,0,168,0,82,0,0,0,233,0,163,0,193,0,124,0,34,0,139,0,198,0,0,0,1,0,112,0,148,0,146,0,28,0,32,0,31,0,0,0,206,0,32,0,140,0,205,0,82,0,228,0,203,0,95,0,189,0,161,0,1,0,78,0,97,0,0,0,173,0,179,0,80,0,222,0,201,0,187,0,180,0,0,0,254,0,212,0,23,0,222,0,233,0,168,0);
signal scenario_full  : scenario_type := (3,31,167,31,167,30,31,31,80,31,89,31,89,30,50,31,221,31,36,31,36,30,36,29,36,28,178,31,161,31,159,31,237,31,139,31,139,30,216,31,62,31,4,31,129,31,129,30,129,29,83,31,174,31,174,30,221,31,46,31,46,30,46,29,94,31,58,31,184,31,22,31,25,31,121,31,165,31,232,31,180,31,25,31,36,31,211,31,69,31,82,31,120,31,234,31,94,31,197,31,197,30,153,31,115,31,170,31,132,31,94,31,145,31,255,31,71,31,71,30,224,31,224,30,252,31,92,31,243,31,133,31,78,31,191,31,191,30,211,31,128,31,128,30,128,29,96,31,156,31,29,31,225,31,225,30,225,29,63,31,63,30,63,29,8,31,180,31,190,31,5,31,159,31,211,31,83,31,251,31,251,30,168,31,168,30,154,31,71,31,153,31,125,31,200,31,200,30,188,31,62,31,118,31,183,31,184,31,87,31,87,30,88,31,88,30,169,31,169,30,157,31,183,31,134,31,27,31,34,31,97,31,75,31,142,31,162,31,186,31,216,31,126,31,191,31,127,31,143,31,143,30,70,31,92,31,92,30,26,31,239,31,191,31,121,31,125,31,125,30,113,31,195,31,14,31,14,30,249,31,249,30,67,31,199,31,199,30,71,31,34,31,149,31,210,31,209,31,116,31,24,31,24,30,24,29,66,31,192,31,59,31,236,31,225,31,57,31,189,31,9,31,134,31,105,31,178,31,164,31,47,31,165,31,215,31,26,31,179,31,36,31,36,30,137,31,65,31,243,31,243,30,223,31,223,30,223,29,142,31,202,31,202,30,78,31,47,31,80,31,114,31,29,31,141,31,251,31,226,31,226,30,129,31,113,31,5,31,179,31,180,31,103,31,165,31,58,31,58,30,82,31,107,31,29,31,63,31,108,31,69,31,205,31,243,31,137,31,137,30,181,31,233,31,233,30,233,29,46,31,98,31,98,30,228,31,26,31,26,30,244,31,219,31,15,31,255,31,175,31,26,31,112,31,240,31,63,31,147,31,143,31,143,30,144,31,249,31,36,31,36,30,200,31,53,31,17,31,47,31,144,31,143,31,42,31,42,30,53,31,121,31,190,31,230,31,30,31,251,31,249,31,30,31,217,31,217,30,90,31,224,31,224,30,224,29,30,31,130,31,130,30,46,31,69,31,247,31,175,31,136,31,1,31,176,31,150,31,83,31,170,31,8,31,202,31,11,31,142,31,246,31,34,31,135,31,75,31,75,30,2,31,107,31,6,31,6,30,6,29,209,31,232,31,142,31,223,31,223,30,61,31,175,31,31,31,31,30,191,31,4,31,175,31,40,31,214,31,178,31,53,31,122,31,78,31,227,31,227,30,69,31,233,31,148,31,148,30,117,31,174,31,175,31,181,31,168,31,12,31,108,31,108,30,97,31,97,30,80,31,44,31,44,31,150,31,150,30,175,31,183,31,183,30,80,31,80,30,80,29,200,31,6,31,156,31,100,31,100,30,95,31,172,31,172,30,116,31,166,31,233,31,253,31,187,31,62,31,204,31,213,31,213,30,47,31,209,31,126,31,232,31,74,31,71,31,166,31,166,30,251,31,142,31,219,31,219,30,140,31,148,31,178,31,178,30,180,31,177,31,191,31,114,31,233,31,224,31,224,30,255,31,143,31,98,31,143,31,144,31,116,31,221,31,40,31,199,31,169,31,126,31,121,31,240,31,210,31,100,31,105,31,66,31,214,31,205,31,140,31,140,30,133,31,24,31,199,31,106,31,232,31,101,31,92,31,9,31,84,31,128,31,152,31,225,31,45,31,219,31,185,31,231,31,75,31,200,31,160,31,160,30,208,31,168,31,202,31,95,31,246,31,55,31,223,31,18,31,142,31,142,30,227,31,175,31,225,31,6,31,66,31,201,31,127,31,225,31,21,31,58,31,66,31,34,31,40,31,40,30,197,31,197,30,205,31,157,31,193,31,193,30,132,31,132,30,232,31,99,31,85,31,25,31,25,30,233,31,233,30,107,31,184,31,106,31,60,31,60,30,60,29,214,31,152,31,177,31,49,31,60,31,60,30,60,29,60,28,115,31,87,31,207,31,126,31,26,31,14,31,65,31,65,30,64,31,202,31,144,31,118,31,7,31,148,31,45,31,45,30,68,31,37,31,89,31,128,31,19,31,238,31,4,31,132,31,38,31,38,30,1,31,1,30,26,31,211,31,78,31,176,31,107,31,203,31,205,31,205,30,205,29,205,31,191,31,150,31,122,31,122,30,13,31,238,31,238,30,89,31,21,31,254,31,19,31,19,30,19,29,170,31,170,30,138,31,118,31,183,31,183,30,40,31,191,31,191,30,123,31,109,31,239,31,154,31,88,31,56,31,135,31,86,31,248,31,94,31,140,31,140,30,153,31,159,31,159,30,159,31,247,31,247,30,247,29,164,31,164,30,155,31,24,31,105,31,123,31,6,31,110,31,97,31,205,31,108,31,195,31,82,31,7,31,7,30,199,31,199,30,156,31,134,31,134,30,123,31,106,31,167,31,255,31,184,31,7,31,97,31,97,30,88,31,88,30,204,31,248,31,248,30,248,29,148,31,241,31,239,31,127,31,114,31,77,31,77,30,176,31,171,31,171,30,183,31,152,31,224,31,156,31,190,31,190,30,190,29,159,31,90,31,192,31,207,31,51,31,38,31,40,31,192,31,169,31,82,31,213,31,231,31,90,31,90,30,143,31,108,31,108,30,108,29,69,31,33,31,65,31,59,31,204,31,204,30,36,31,36,30,36,29,131,31,131,30,131,29,206,31,192,31,111,31,233,31,233,30,23,31,23,30,118,31,64,31,64,30,64,29,64,28,189,31,134,31,89,31,204,31,92,31,92,30,107,31,141,31,5,31,5,30,15,31,142,31,142,30,246,31,246,30,246,29,246,28,38,31,221,31,133,31,133,30,255,31,160,31,160,30,160,29,100,31,139,31,192,31,177,31,99,31,29,31,236,31,216,31,216,30,158,31,228,31,49,31,194,31,226,31,123,31,126,31,53,31,70,31,88,31,94,31,158,31,115,31,194,31,83,31,83,30,61,31,98,31,170,31,81,31,81,30,81,29,178,31,178,30,230,31,227,31,64,31,205,31,17,31,189,31,228,31,238,31,35,31,86,31,147,31,27,31,76,31,87,31,231,31,227,31,98,31,98,30,98,29,85,31,247,31,73,31,44,31,159,31,74,31,217,31,244,31,134,31,19,31,128,31,86,31,168,31,82,31,82,30,233,31,163,31,193,31,124,31,34,31,139,31,198,31,198,30,1,31,112,31,148,31,146,31,28,31,32,31,31,31,31,30,206,31,32,31,140,31,205,31,82,31,228,31,203,31,95,31,189,31,161,31,1,31,78,31,97,31,97,30,173,31,179,31,80,31,222,31,201,31,187,31,180,31,180,30,254,31,212,31,23,31,222,31,233,31,168,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
