-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_659 is
end project_tb_659;

architecture project_tb_arch_659 of project_tb_659 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 939;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (73,0,194,0,52,0,232,0,228,0,240,0,0,0,13,0,179,0,229,0,35,0,21,0,214,0,228,0,204,0,215,0,0,0,217,0,246,0,138,0,79,0,148,0,102,0,150,0,211,0,164,0,214,0,45,0,0,0,12,0,200,0,0,0,0,0,0,0,0,0,0,0,159,0,210,0,217,0,61,0,53,0,0,0,19,0,196,0,209,0,178,0,199,0,0,0,166,0,0,0,0,0,20,0,124,0,91,0,187,0,62,0,51,0,11,0,117,0,188,0,193,0,165,0,254,0,238,0,0,0,234,0,126,0,155,0,107,0,0,0,0,0,235,0,116,0,209,0,204,0,255,0,58,0,124,0,0,0,161,0,0,0,159,0,106,0,4,0,17,0,208,0,147,0,0,0,222,0,140,0,115,0,243,0,0,0,0,0,0,0,201,0,0,0,14,0,66,0,0,0,250,0,177,0,76,0,133,0,0,0,205,0,233,0,179,0,60,0,30,0,69,0,240,0,0,0,46,0,177,0,153,0,71,0,34,0,41,0,64,0,153,0,39,0,52,0,0,0,73,0,238,0,189,0,122,0,167,0,0,0,234,0,0,0,119,0,101,0,50,0,40,0,31,0,0,0,199,0,163,0,38,0,174,0,0,0,130,0,165,0,212,0,183,0,0,0,85,0,194,0,111,0,113,0,241,0,56,0,0,0,179,0,131,0,42,0,223,0,0,0,229,0,70,0,137,0,181,0,249,0,34,0,139,0,0,0,247,0,231,0,0,0,0,0,30,0,0,0,122,0,97,0,0,0,212,0,232,0,78,0,158,0,167,0,103,0,93,0,7,0,255,0,220,0,0,0,0,0,0,0,142,0,252,0,0,0,155,0,5,0,0,0,5,0,178,0,151,0,26,0,9,0,8,0,124,0,79,0,94,0,25,0,73,0,0,0,197,0,36,0,20,0,138,0,0,0,216,0,209,0,95,0,0,0,32,0,105,0,194,0,34,0,208,0,0,0,59,0,102,0,186,0,171,0,80,0,0,0,39,0,23,0,183,0,223,0,186,0,134,0,233,0,223,0,88,0,71,0,6,0,48,0,0,0,15,0,59,0,11,0,214,0,238,0,118,0,199,0,112,0,65,0,3,0,188,0,216,0,25,0,91,0,208,0,0,0,190,0,0,0,181,0,149,0,233,0,0,0,45,0,117,0,123,0,110,0,60,0,174,0,83,0,148,0,211,0,214,0,86,0,66,0,0,0,0,0,1,0,214,0,58,0,228,0,73,0,0,0,0,0,57,0,37,0,139,0,116,0,24,0,168,0,0,0,125,0,188,0,105,0,111,0,0,0,0,0,97,0,0,0,59,0,197,0,76,0,236,0,208,0,0,0,109,0,185,0,151,0,125,0,136,0,28,0,0,0,193,0,158,0,3,0,76,0,152,0,107,0,148,0,26,0,37,0,37,0,145,0,91,0,6,0,245,0,182,0,58,0,183,0,0,0,57,0,6,0,142,0,191,0,62,0,116,0,18,0,0,0,225,0,109,0,0,0,104,0,138,0,0,0,130,0,49,0,0,0,152,0,128,0,22,0,58,0,21,0,0,0,0,0,116,0,32,0,195,0,231,0,241,0,201,0,68,0,169,0,152,0,53,0,145,0,0,0,110,0,47,0,40,0,204,0,135,0,40,0,0,0,174,0,213,0,246,0,99,0,242,0,133,0,85,0,139,0,70,0,190,0,139,0,213,0,147,0,43,0,137,0,0,0,95,0,217,0,0,0,183,0,110,0,180,0,159,0,95,0,129,0,185,0,16,0,68,0,144,0,130,0,0,0,24,0,114,0,26,0,211,0,0,0,0,0,70,0,139,0,213,0,45,0,108,0,188,0,0,0,74,0,100,0,161,0,236,0,17,0,81,0,185,0,0,0,20,0,7,0,0,0,215,0,75,0,251,0,75,0,0,0,0,0,91,0,0,0,255,0,93,0,28,0,32,0,160,0,192,0,0,0,0,0,136,0,206,0,184,0,77,0,11,0,249,0,204,0,175,0,14,0,167,0,0,0,97,0,115,0,225,0,82,0,124,0,170,0,99,0,215,0,210,0,214,0,197,0,195,0,49,0,78,0,142,0,63,0,94,0,47,0,7,0,0,0,132,0,76,0,159,0,37,0,92,0,12,0,115,0,153,0,0,0,0,0,119,0,74,0,0,0,0,0,161,0,0,0,196,0,161,0,0,0,0,0,36,0,47,0,161,0,26,0,36,0,9,0,0,0,242,0,196,0,206,0,204,0,237,0,178,0,178,0,116,0,43,0,0,0,250,0,120,0,31,0,18,0,224,0,0,0,239,0,224,0,228,0,0,0,85,0,131,0,13,0,0,0,125,0,86,0,126,0,0,0,182,0,103,0,62,0,246,0,145,0,45,0,213,0,89,0,189,0,0,0,101,0,6,0,101,0,0,0,69,0,163,0,33,0,44,0,7,0,154,0,124,0,205,0,18,0,0,0,0,0,112,0,150,0,55,0,37,0,214,0,213,0,154,0,154,0,8,0,120,0,134,0,5,0,0,0,93,0,52,0,105,0,133,0,49,0,0,0,203,0,223,0,29,0,147,0,71,0,112,0,251,0,0,0,134,0,199,0,39,0,45,0,119,0,226,0,185,0,240,0,136,0,63,0,205,0,17,0,0,0,137,0,160,0,117,0,210,0,46,0,90,0,0,0,44,0,180,0,66,0,0,0,110,0,20,0,250,0,164,0,31,0,131,0,0,0,227,0,202,0,244,0,142,0,128,0,0,0,152,0,223,0,247,0,136,0,64,0,165,0,238,0,0,0,210,0,239,0,150,0,22,0,237,0,11,0,44,0,182,0,250,0,254,0,0,0,236,0,154,0,144,0,185,0,177,0,0,0,121,0,0,0,248,0,244,0,235,0,40,0,72,0,52,0,0,0,53,0,30,0,245,0,0,0,47,0,0,0,250,0,105,0,36,0,13,0,0,0,115,0,74,0,178,0,0,0,41,0,131,0,41,0,142,0,157,0,0,0,15,0,114,0,93,0,4,0,65,0,96,0,39,0,0,0,203,0,43,0,0,0,125,0,65,0,244,0,185,0,160,0,238,0,211,0,13,0,135,0,152,0,78,0,42,0,182,0,233,0,193,0,0,0,189,0,177,0,186,0,0,0,109,0,0,0,82,0,229,0,145,0,248,0,0,0,114,0,0,0,169,0,0,0,244,0,0,0,24,0,194,0,198,0,144,0,0,0,144,0,212,0,110,0,0,0,250,0,116,0,244,0,133,0,20,0,196,0,0,0,184,0,207,0,65,0,75,0,0,0,12,0,0,0,0,0,0,0,91,0,50,0,10,0,76,0,18,0,130,0,0,0,152,0,176,0,0,0,96,0,188,0,194,0,0,0,62,0,95,0,101,0,210,0,0,0,136,0,106,0,137,0,0,0,60,0,31,0,100,0,45,0,0,0,0,0,176,0,0,0,52,0,120,0,146,0,23,0,0,0,0,0,117,0,71,0,146,0,30,0,146,0,5,0,240,0,208,0,123,0,1,0,120,0,115,0,193,0,23,0,20,0,211,0,141,0,67,0,111,0,29,0,62,0,139,0,94,0,27,0,108,0,201,0,171,0,0,0,77,0,153,0,150,0,169,0,124,0,219,0,0,0,240,0,0,0,108,0,0,0,0,0,0,0,43,0,62,0,117,0,0,0,52,0,0,0,248,0,183,0,0,0,239,0,31,0,58,0,8,0,40,0,84,0,108,0,200,0,0,0,123,0,245,0,215,0,186,0,139,0,130,0,228,0,0,0,28,0,31,0,212,0,35,0,84,0,168,0,248,0,9,0,166,0,215,0,192,0,186,0,180,0,112,0,62,0,95,0,91,0,251,0,142,0,190,0,13,0,87,0,11,0,201,0,47,0,0,0,248,0,49,0,0,0,63,0,227,0,49,0,189,0,0,0,231,0,161,0,21,0,0,0,0,0,168,0,0,0,118,0,36,0,166,0,142,0,0,0,144,0,76,0,0,0,0,0,41,0,35,0,75,0,36,0,19,0,186,0,159,0,56,0,181,0,147,0,82,0,247,0,24,0,111,0,70,0,0,0,40,0,216,0,90,0,19,0,0,0,83,0,194,0,106,0,194,0,204,0,150,0,0,0,67,0,145,0,51,0,50,0,67,0,0,0,105,0,0,0,52,0,8,0,118,0,0,0,33,0);
signal scenario_full  : scenario_type := (73,31,194,31,52,31,232,31,228,31,240,31,240,30,13,31,179,31,229,31,35,31,21,31,214,31,228,31,204,31,215,31,215,30,217,31,246,31,138,31,79,31,148,31,102,31,150,31,211,31,164,31,214,31,45,31,45,30,12,31,200,31,200,30,200,29,200,28,200,27,200,26,159,31,210,31,217,31,61,31,53,31,53,30,19,31,196,31,209,31,178,31,199,31,199,30,166,31,166,30,166,29,20,31,124,31,91,31,187,31,62,31,51,31,11,31,117,31,188,31,193,31,165,31,254,31,238,31,238,30,234,31,126,31,155,31,107,31,107,30,107,29,235,31,116,31,209,31,204,31,255,31,58,31,124,31,124,30,161,31,161,30,159,31,106,31,4,31,17,31,208,31,147,31,147,30,222,31,140,31,115,31,243,31,243,30,243,29,243,28,201,31,201,30,14,31,66,31,66,30,250,31,177,31,76,31,133,31,133,30,205,31,233,31,179,31,60,31,30,31,69,31,240,31,240,30,46,31,177,31,153,31,71,31,34,31,41,31,64,31,153,31,39,31,52,31,52,30,73,31,238,31,189,31,122,31,167,31,167,30,234,31,234,30,119,31,101,31,50,31,40,31,31,31,31,30,199,31,163,31,38,31,174,31,174,30,130,31,165,31,212,31,183,31,183,30,85,31,194,31,111,31,113,31,241,31,56,31,56,30,179,31,131,31,42,31,223,31,223,30,229,31,70,31,137,31,181,31,249,31,34,31,139,31,139,30,247,31,231,31,231,30,231,29,30,31,30,30,122,31,97,31,97,30,212,31,232,31,78,31,158,31,167,31,103,31,93,31,7,31,255,31,220,31,220,30,220,29,220,28,142,31,252,31,252,30,155,31,5,31,5,30,5,31,178,31,151,31,26,31,9,31,8,31,124,31,79,31,94,31,25,31,73,31,73,30,197,31,36,31,20,31,138,31,138,30,216,31,209,31,95,31,95,30,32,31,105,31,194,31,34,31,208,31,208,30,59,31,102,31,186,31,171,31,80,31,80,30,39,31,23,31,183,31,223,31,186,31,134,31,233,31,223,31,88,31,71,31,6,31,48,31,48,30,15,31,59,31,11,31,214,31,238,31,118,31,199,31,112,31,65,31,3,31,188,31,216,31,25,31,91,31,208,31,208,30,190,31,190,30,181,31,149,31,233,31,233,30,45,31,117,31,123,31,110,31,60,31,174,31,83,31,148,31,211,31,214,31,86,31,66,31,66,30,66,29,1,31,214,31,58,31,228,31,73,31,73,30,73,29,57,31,37,31,139,31,116,31,24,31,168,31,168,30,125,31,188,31,105,31,111,31,111,30,111,29,97,31,97,30,59,31,197,31,76,31,236,31,208,31,208,30,109,31,185,31,151,31,125,31,136,31,28,31,28,30,193,31,158,31,3,31,76,31,152,31,107,31,148,31,26,31,37,31,37,31,145,31,91,31,6,31,245,31,182,31,58,31,183,31,183,30,57,31,6,31,142,31,191,31,62,31,116,31,18,31,18,30,225,31,109,31,109,30,104,31,138,31,138,30,130,31,49,31,49,30,152,31,128,31,22,31,58,31,21,31,21,30,21,29,116,31,32,31,195,31,231,31,241,31,201,31,68,31,169,31,152,31,53,31,145,31,145,30,110,31,47,31,40,31,204,31,135,31,40,31,40,30,174,31,213,31,246,31,99,31,242,31,133,31,85,31,139,31,70,31,190,31,139,31,213,31,147,31,43,31,137,31,137,30,95,31,217,31,217,30,183,31,110,31,180,31,159,31,95,31,129,31,185,31,16,31,68,31,144,31,130,31,130,30,24,31,114,31,26,31,211,31,211,30,211,29,70,31,139,31,213,31,45,31,108,31,188,31,188,30,74,31,100,31,161,31,236,31,17,31,81,31,185,31,185,30,20,31,7,31,7,30,215,31,75,31,251,31,75,31,75,30,75,29,91,31,91,30,255,31,93,31,28,31,32,31,160,31,192,31,192,30,192,29,136,31,206,31,184,31,77,31,11,31,249,31,204,31,175,31,14,31,167,31,167,30,97,31,115,31,225,31,82,31,124,31,170,31,99,31,215,31,210,31,214,31,197,31,195,31,49,31,78,31,142,31,63,31,94,31,47,31,7,31,7,30,132,31,76,31,159,31,37,31,92,31,12,31,115,31,153,31,153,30,153,29,119,31,74,31,74,30,74,29,161,31,161,30,196,31,161,31,161,30,161,29,36,31,47,31,161,31,26,31,36,31,9,31,9,30,242,31,196,31,206,31,204,31,237,31,178,31,178,31,116,31,43,31,43,30,250,31,120,31,31,31,18,31,224,31,224,30,239,31,224,31,228,31,228,30,85,31,131,31,13,31,13,30,125,31,86,31,126,31,126,30,182,31,103,31,62,31,246,31,145,31,45,31,213,31,89,31,189,31,189,30,101,31,6,31,101,31,101,30,69,31,163,31,33,31,44,31,7,31,154,31,124,31,205,31,18,31,18,30,18,29,112,31,150,31,55,31,37,31,214,31,213,31,154,31,154,31,8,31,120,31,134,31,5,31,5,30,93,31,52,31,105,31,133,31,49,31,49,30,203,31,223,31,29,31,147,31,71,31,112,31,251,31,251,30,134,31,199,31,39,31,45,31,119,31,226,31,185,31,240,31,136,31,63,31,205,31,17,31,17,30,137,31,160,31,117,31,210,31,46,31,90,31,90,30,44,31,180,31,66,31,66,30,110,31,20,31,250,31,164,31,31,31,131,31,131,30,227,31,202,31,244,31,142,31,128,31,128,30,152,31,223,31,247,31,136,31,64,31,165,31,238,31,238,30,210,31,239,31,150,31,22,31,237,31,11,31,44,31,182,31,250,31,254,31,254,30,236,31,154,31,144,31,185,31,177,31,177,30,121,31,121,30,248,31,244,31,235,31,40,31,72,31,52,31,52,30,53,31,30,31,245,31,245,30,47,31,47,30,250,31,105,31,36,31,13,31,13,30,115,31,74,31,178,31,178,30,41,31,131,31,41,31,142,31,157,31,157,30,15,31,114,31,93,31,4,31,65,31,96,31,39,31,39,30,203,31,43,31,43,30,125,31,65,31,244,31,185,31,160,31,238,31,211,31,13,31,135,31,152,31,78,31,42,31,182,31,233,31,193,31,193,30,189,31,177,31,186,31,186,30,109,31,109,30,82,31,229,31,145,31,248,31,248,30,114,31,114,30,169,31,169,30,244,31,244,30,24,31,194,31,198,31,144,31,144,30,144,31,212,31,110,31,110,30,250,31,116,31,244,31,133,31,20,31,196,31,196,30,184,31,207,31,65,31,75,31,75,30,12,31,12,30,12,29,12,28,91,31,50,31,10,31,76,31,18,31,130,31,130,30,152,31,176,31,176,30,96,31,188,31,194,31,194,30,62,31,95,31,101,31,210,31,210,30,136,31,106,31,137,31,137,30,60,31,31,31,100,31,45,31,45,30,45,29,176,31,176,30,52,31,120,31,146,31,23,31,23,30,23,29,117,31,71,31,146,31,30,31,146,31,5,31,240,31,208,31,123,31,1,31,120,31,115,31,193,31,23,31,20,31,211,31,141,31,67,31,111,31,29,31,62,31,139,31,94,31,27,31,108,31,201,31,171,31,171,30,77,31,153,31,150,31,169,31,124,31,219,31,219,30,240,31,240,30,108,31,108,30,108,29,108,28,43,31,62,31,117,31,117,30,52,31,52,30,248,31,183,31,183,30,239,31,31,31,58,31,8,31,40,31,84,31,108,31,200,31,200,30,123,31,245,31,215,31,186,31,139,31,130,31,228,31,228,30,28,31,31,31,212,31,35,31,84,31,168,31,248,31,9,31,166,31,215,31,192,31,186,31,180,31,112,31,62,31,95,31,91,31,251,31,142,31,190,31,13,31,87,31,11,31,201,31,47,31,47,30,248,31,49,31,49,30,63,31,227,31,49,31,189,31,189,30,231,31,161,31,21,31,21,30,21,29,168,31,168,30,118,31,36,31,166,31,142,31,142,30,144,31,76,31,76,30,76,29,41,31,35,31,75,31,36,31,19,31,186,31,159,31,56,31,181,31,147,31,82,31,247,31,24,31,111,31,70,31,70,30,40,31,216,31,90,31,19,31,19,30,83,31,194,31,106,31,194,31,204,31,150,31,150,30,67,31,145,31,51,31,50,31,67,31,67,30,105,31,105,30,52,31,8,31,118,31,118,30,33,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
