-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 833;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (183,0,220,0,252,0,108,0,73,0,153,0,81,0,0,0,0,0,103,0,221,0,0,0,0,0,135,0,132,0,149,0,24,0,0,0,105,0,0,0,43,0,249,0,54,0,0,0,59,0,0,0,214,0,0,0,68,0,0,0,0,0,17,0,0,0,82,0,0,0,36,0,224,0,114,0,0,0,235,0,226,0,21,0,86,0,112,0,0,0,0,0,0,0,26,0,0,0,226,0,193,0,84,0,232,0,211,0,150,0,138,0,179,0,185,0,0,0,204,0,113,0,0,0,73,0,0,0,96,0,164,0,6,0,213,0,98,0,188,0,116,0,44,0,116,0,75,0,159,0,112,0,197,0,248,0,130,0,191,0,115,0,252,0,211,0,217,0,44,0,0,0,215,0,251,0,181,0,0,0,233,0,221,0,213,0,0,0,0,0,43,0,42,0,191,0,0,0,113,0,2,0,49,0,0,0,3,0,125,0,37,0,0,0,0,0,0,0,114,0,111,0,113,0,106,0,89,0,0,0,161,0,237,0,26,0,246,0,0,0,160,0,0,0,118,0,48,0,220,0,72,0,0,0,102,0,15,0,27,0,56,0,159,0,116,0,118,0,121,0,28,0,37,0,225,0,0,0,0,0,20,0,0,0,14,0,63,0,178,0,0,0,178,0,196,0,169,0,170,0,61,0,178,0,237,0,158,0,0,0,9,0,204,0,192,0,0,0,82,0,191,0,0,0,212,0,56,0,249,0,42,0,0,0,124,0,75,0,251,0,189,0,0,0,224,0,221,0,61,0,0,0,123,0,143,0,39,0,64,0,0,0,46,0,123,0,49,0,227,0,103,0,28,0,134,0,151,0,127,0,157,0,237,0,95,0,147,0,156,0,87,0,198,0,144,0,100,0,88,0,125,0,189,0,44,0,0,0,0,0,63,0,17,0,0,0,227,0,111,0,134,0,205,0,80,0,205,0,219,0,7,0,46,0,34,0,41,0,98,0,188,0,19,0,0,0,0,0,0,0,1,0,199,0,39,0,37,0,10,0,190,0,50,0,0,0,28,0,190,0,39,0,46,0,2,0,0,0,127,0,90,0,13,0,151,0,18,0,156,0,0,0,146,0,51,0,60,0,176,0,49,0,107,0,85,0,142,0,85,0,153,0,16,0,124,0,70,0,0,0,42,0,133,0,123,0,93,0,218,0,1,0,0,0,222,0,24,0,115,0,210,0,134,0,238,0,111,0,252,0,23,0,224,0,0,0,178,0,204,0,207,0,139,0,62,0,25,0,119,0,129,0,93,0,54,0,0,0,181,0,36,0,92,0,207,0,135,0,123,0,150,0,182,0,0,0,234,0,7,0,89,0,72,0,202,0,0,0,75,0,24,0,205,0,189,0,36,0,102,0,98,0,173,0,142,0,81,0,0,0,73,0,0,0,29,0,0,0,120,0,8,0,248,0,70,0,199,0,173,0,69,0,66,0,43,0,165,0,71,0,232,0,29,0,8,0,27,0,0,0,28,0,0,0,191,0,244,0,1,0,31,0,97,0,71,0,45,0,229,0,74,0,112,0,77,0,119,0,4,0,4,0,163,0,139,0,193,0,0,0,163,0,68,0,0,0,176,0,0,0,76,0,145,0,178,0,40,0,0,0,141,0,0,0,249,0,173,0,8,0,71,0,61,0,0,0,15,0,52,0,111,0,160,0,0,0,160,0,0,0,84,0,167,0,188,0,116,0,140,0,0,0,0,0,105,0,170,0,30,0,241,0,159,0,172,0,22,0,244,0,142,0,135,0,0,0,230,0,32,0,0,0,27,0,252,0,88,0,56,0,232,0,189,0,244,0,41,0,164,0,97,0,87,0,96,0,72,0,195,0,56,0,0,0,11,0,182,0,0,0,74,0,3,0,0,0,0,0,0,0,181,0,200,0,138,0,0,0,38,0,187,0,6,0,234,0,187,0,183,0,118,0,0,0,234,0,147,0,193,0,54,0,7,0,3,0,8,0,24,0,179,0,89,0,34,0,86,0,126,0,86,0,65,0,0,0,0,0,236,0,104,0,0,0,70,0,204,0,44,0,153,0,113,0,0,0,232,0,86,0,240,0,236,0,229,0,181,0,19,0,131,0,186,0,47,0,26,0,0,0,37,0,28,0,24,0,0,0,19,0,183,0,0,0,187,0,120,0,130,0,138,0,13,0,242,0,7,0,139,0,165,0,20,0,35,0,0,0,141,0,33,0,227,0,249,0,111,0,0,0,43,0,151,0,176,0,19,0,102,0,30,0,81,0,171,0,0,0,0,0,206,0,76,0,0,0,124,0,103,0,23,0,228,0,69,0,130,0,10,0,151,0,80,0,169,0,237,0,0,0,146,0,219,0,132,0,194,0,28,0,8,0,33,0,0,0,253,0,16,0,105,0,0,0,106,0,180,0,0,0,0,0,90,0,92,0,28,0,230,0,243,0,106,0,27,0,209,0,57,0,119,0,201,0,62,0,228,0,80,0,0,0,123,0,160,0,0,0,177,0,0,0,239,0,0,0,0,0,0,0,40,0,225,0,14,0,0,0,52,0,232,0,141,0,10,0,0,0,5,0,8,0,31,0,139,0,3,0,12,0,0,0,0,0,67,0,195,0,0,0,80,0,140,0,36,0,23,0,22,0,138,0,255,0,0,0,189,0,0,0,0,0,164,0,179,0,46,0,216,0,24,0,0,0,0,0,47,0,0,0,0,0,230,0,6,0,59,0,240,0,151,0,199,0,181,0,203,0,0,0,37,0,169,0,145,0,120,0,235,0,17,0,106,0,185,0,28,0,133,0,224,0,0,0,206,0,88,0,0,0,37,0,42,0,71,0,0,0,132,0,61,0,74,0,66,0,74,0,62,0,45,0,170,0,148,0,139,0,78,0,84,0,193,0,165,0,162,0,18,0,51,0,118,0,0,0,183,0,21,0,195,0,239,0,238,0,103,0,0,0,222,0,186,0,91,0,182,0,233,0,0,0,12,0,230,0,56,0,97,0,10,0,101,0,0,0,178,0,141,0,0,0,29,0,75,0,164,0,120,0,0,0,0,0,110,0,0,0,1,0,67,0,246,0,0,0,68,0,119,0,27,0,0,0,196,0,249,0,17,0,0,0,0,0,242,0,212,0,0,0,0,0,233,0,46,0,115,0,111,0,84,0,137,0,7,0,51,0,201,0,118,0,151,0,63,0,252,0,0,0,0,0,0,0,0,0,110,0,0,0,33,0,175,0,99,0,167,0,250,0,0,0,26,0,197,0,229,0,84,0,151,0,107,0,153,0,0,0,82,0,29,0,48,0,30,0,216,0,64,0,192,0,0,0,0,0,101,0,191,0,4,0,32,0,0,0,87,0,52,0,248,0,144,0,0,0,140,0,159,0,170,0,22,0,130,0,145,0,149,0,73,0,242,0,116,0,0,0,153,0,229,0,235,0,116,0,0,0,243,0,171,0,168,0,58,0,242,0,0,0,204,0,1,0,81,0,171,0,209,0,0,0,0,0,54,0,126,0,207,0,157,0,232,0,158,0,77,0,59,0,239,0,0,0,108,0,87,0,131,0,65,0,0,0,92,0,214,0,0,0,11,0,199,0,196,0,32,0,124,0,49,0,37,0,0,0,0,0,150,0,0,0,22,0,0,0,98,0,195,0,0,0,0,0,168,0,97,0,247,0,203,0,180,0,96,0,43,0,70,0,0,0,201,0,0,0,239,0,153,0,120,0,170,0,207,0);
signal scenario_full  : scenario_type := (183,31,220,31,252,31,108,31,73,31,153,31,81,31,81,30,81,29,103,31,221,31,221,30,221,29,135,31,132,31,149,31,24,31,24,30,105,31,105,30,43,31,249,31,54,31,54,30,59,31,59,30,214,31,214,30,68,31,68,30,68,29,17,31,17,30,82,31,82,30,36,31,224,31,114,31,114,30,235,31,226,31,21,31,86,31,112,31,112,30,112,29,112,28,26,31,26,30,226,31,193,31,84,31,232,31,211,31,150,31,138,31,179,31,185,31,185,30,204,31,113,31,113,30,73,31,73,30,96,31,164,31,6,31,213,31,98,31,188,31,116,31,44,31,116,31,75,31,159,31,112,31,197,31,248,31,130,31,191,31,115,31,252,31,211,31,217,31,44,31,44,30,215,31,251,31,181,31,181,30,233,31,221,31,213,31,213,30,213,29,43,31,42,31,191,31,191,30,113,31,2,31,49,31,49,30,3,31,125,31,37,31,37,30,37,29,37,28,114,31,111,31,113,31,106,31,89,31,89,30,161,31,237,31,26,31,246,31,246,30,160,31,160,30,118,31,48,31,220,31,72,31,72,30,102,31,15,31,27,31,56,31,159,31,116,31,118,31,121,31,28,31,37,31,225,31,225,30,225,29,20,31,20,30,14,31,63,31,178,31,178,30,178,31,196,31,169,31,170,31,61,31,178,31,237,31,158,31,158,30,9,31,204,31,192,31,192,30,82,31,191,31,191,30,212,31,56,31,249,31,42,31,42,30,124,31,75,31,251,31,189,31,189,30,224,31,221,31,61,31,61,30,123,31,143,31,39,31,64,31,64,30,46,31,123,31,49,31,227,31,103,31,28,31,134,31,151,31,127,31,157,31,237,31,95,31,147,31,156,31,87,31,198,31,144,31,100,31,88,31,125,31,189,31,44,31,44,30,44,29,63,31,17,31,17,30,227,31,111,31,134,31,205,31,80,31,205,31,219,31,7,31,46,31,34,31,41,31,98,31,188,31,19,31,19,30,19,29,19,28,1,31,199,31,39,31,37,31,10,31,190,31,50,31,50,30,28,31,190,31,39,31,46,31,2,31,2,30,127,31,90,31,13,31,151,31,18,31,156,31,156,30,146,31,51,31,60,31,176,31,49,31,107,31,85,31,142,31,85,31,153,31,16,31,124,31,70,31,70,30,42,31,133,31,123,31,93,31,218,31,1,31,1,30,222,31,24,31,115,31,210,31,134,31,238,31,111,31,252,31,23,31,224,31,224,30,178,31,204,31,207,31,139,31,62,31,25,31,119,31,129,31,93,31,54,31,54,30,181,31,36,31,92,31,207,31,135,31,123,31,150,31,182,31,182,30,234,31,7,31,89,31,72,31,202,31,202,30,75,31,24,31,205,31,189,31,36,31,102,31,98,31,173,31,142,31,81,31,81,30,73,31,73,30,29,31,29,30,120,31,8,31,248,31,70,31,199,31,173,31,69,31,66,31,43,31,165,31,71,31,232,31,29,31,8,31,27,31,27,30,28,31,28,30,191,31,244,31,1,31,31,31,97,31,71,31,45,31,229,31,74,31,112,31,77,31,119,31,4,31,4,31,163,31,139,31,193,31,193,30,163,31,68,31,68,30,176,31,176,30,76,31,145,31,178,31,40,31,40,30,141,31,141,30,249,31,173,31,8,31,71,31,61,31,61,30,15,31,52,31,111,31,160,31,160,30,160,31,160,30,84,31,167,31,188,31,116,31,140,31,140,30,140,29,105,31,170,31,30,31,241,31,159,31,172,31,22,31,244,31,142,31,135,31,135,30,230,31,32,31,32,30,27,31,252,31,88,31,56,31,232,31,189,31,244,31,41,31,164,31,97,31,87,31,96,31,72,31,195,31,56,31,56,30,11,31,182,31,182,30,74,31,3,31,3,30,3,29,3,28,181,31,200,31,138,31,138,30,38,31,187,31,6,31,234,31,187,31,183,31,118,31,118,30,234,31,147,31,193,31,54,31,7,31,3,31,8,31,24,31,179,31,89,31,34,31,86,31,126,31,86,31,65,31,65,30,65,29,236,31,104,31,104,30,70,31,204,31,44,31,153,31,113,31,113,30,232,31,86,31,240,31,236,31,229,31,181,31,19,31,131,31,186,31,47,31,26,31,26,30,37,31,28,31,24,31,24,30,19,31,183,31,183,30,187,31,120,31,130,31,138,31,13,31,242,31,7,31,139,31,165,31,20,31,35,31,35,30,141,31,33,31,227,31,249,31,111,31,111,30,43,31,151,31,176,31,19,31,102,31,30,31,81,31,171,31,171,30,171,29,206,31,76,31,76,30,124,31,103,31,23,31,228,31,69,31,130,31,10,31,151,31,80,31,169,31,237,31,237,30,146,31,219,31,132,31,194,31,28,31,8,31,33,31,33,30,253,31,16,31,105,31,105,30,106,31,180,31,180,30,180,29,90,31,92,31,28,31,230,31,243,31,106,31,27,31,209,31,57,31,119,31,201,31,62,31,228,31,80,31,80,30,123,31,160,31,160,30,177,31,177,30,239,31,239,30,239,29,239,28,40,31,225,31,14,31,14,30,52,31,232,31,141,31,10,31,10,30,5,31,8,31,31,31,139,31,3,31,12,31,12,30,12,29,67,31,195,31,195,30,80,31,140,31,36,31,23,31,22,31,138,31,255,31,255,30,189,31,189,30,189,29,164,31,179,31,46,31,216,31,24,31,24,30,24,29,47,31,47,30,47,29,230,31,6,31,59,31,240,31,151,31,199,31,181,31,203,31,203,30,37,31,169,31,145,31,120,31,235,31,17,31,106,31,185,31,28,31,133,31,224,31,224,30,206,31,88,31,88,30,37,31,42,31,71,31,71,30,132,31,61,31,74,31,66,31,74,31,62,31,45,31,170,31,148,31,139,31,78,31,84,31,193,31,165,31,162,31,18,31,51,31,118,31,118,30,183,31,21,31,195,31,239,31,238,31,103,31,103,30,222,31,186,31,91,31,182,31,233,31,233,30,12,31,230,31,56,31,97,31,10,31,101,31,101,30,178,31,141,31,141,30,29,31,75,31,164,31,120,31,120,30,120,29,110,31,110,30,1,31,67,31,246,31,246,30,68,31,119,31,27,31,27,30,196,31,249,31,17,31,17,30,17,29,242,31,212,31,212,30,212,29,233,31,46,31,115,31,111,31,84,31,137,31,7,31,51,31,201,31,118,31,151,31,63,31,252,31,252,30,252,29,252,28,252,27,110,31,110,30,33,31,175,31,99,31,167,31,250,31,250,30,26,31,197,31,229,31,84,31,151,31,107,31,153,31,153,30,82,31,29,31,48,31,30,31,216,31,64,31,192,31,192,30,192,29,101,31,191,31,4,31,32,31,32,30,87,31,52,31,248,31,144,31,144,30,140,31,159,31,170,31,22,31,130,31,145,31,149,31,73,31,242,31,116,31,116,30,153,31,229,31,235,31,116,31,116,30,243,31,171,31,168,31,58,31,242,31,242,30,204,31,1,31,81,31,171,31,209,31,209,30,209,29,54,31,126,31,207,31,157,31,232,31,158,31,77,31,59,31,239,31,239,30,108,31,87,31,131,31,65,31,65,30,92,31,214,31,214,30,11,31,199,31,196,31,32,31,124,31,49,31,37,31,37,30,37,29,150,31,150,30,22,31,22,30,98,31,195,31,195,30,195,29,168,31,97,31,247,31,203,31,180,31,96,31,43,31,70,31,70,30,201,31,201,30,239,31,153,31,120,31,170,31,207,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
