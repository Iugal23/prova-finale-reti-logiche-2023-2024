-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1014;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (156,0,0,0,24,0,111,0,239,0,0,0,159,0,140,0,153,0,122,0,149,0,223,0,0,0,0,0,217,0,0,0,165,0,12,0,0,0,59,0,198,0,0,0,0,0,140,0,0,0,133,0,25,0,0,0,205,0,136,0,140,0,24,0,61,0,200,0,52,0,191,0,114,0,231,0,37,0,59,0,15,0,58,0,13,0,78,0,56,0,0,0,45,0,191,0,164,0,253,0,0,0,150,0,69,0,247,0,0,0,36,0,171,0,0,0,0,0,47,0,0,0,182,0,144,0,4,0,19,0,112,0,11,0,211,0,32,0,124,0,100,0,200,0,52,0,23,0,182,0,209,0,211,0,136,0,0,0,242,0,252,0,223,0,0,0,0,0,250,0,218,0,133,0,165,0,61,0,254,0,88,0,153,0,0,0,128,0,66,0,28,0,0,0,0,0,127,0,235,0,109,0,147,0,46,0,164,0,132,0,242,0,52,0,69,0,148,0,245,0,149,0,105,0,88,0,179,0,108,0,0,0,0,0,198,0,4,0,118,0,0,0,160,0,249,0,127,0,230,0,0,0,0,0,18,0,121,0,143,0,115,0,22,0,166,0,0,0,111,0,0,0,155,0,0,0,0,0,226,0,0,0,68,0,93,0,36,0,176,0,0,0,115,0,184,0,169,0,187,0,0,0,0,0,119,0,0,0,155,0,228,0,158,0,231,0,12,0,250,0,165,0,0,0,19,0,206,0,175,0,0,0,166,0,134,0,0,0,0,0,188,0,67,0,133,0,40,0,99,0,84,0,0,0,35,0,249,0,244,0,22,0,71,0,0,0,32,0,255,0,39,0,99,0,64,0,93,0,91,0,227,0,0,0,54,0,15,0,78,0,99,0,119,0,146,0,174,0,0,0,49,0,165,0,222,0,222,0,207,0,213,0,162,0,44,0,46,0,163,0,0,0,207,0,101,0,12,0,218,0,68,0,111,0,156,0,18,0,153,0,254,0,132,0,213,0,76,0,96,0,66,0,153,0,0,0,216,0,161,0,206,0,101,0,82,0,0,0,108,0,141,0,244,0,136,0,124,0,59,0,0,0,80,0,216,0,158,0,93,0,205,0,0,0,188,0,113,0,0,0,251,0,40,0,59,0,247,0,144,0,243,0,132,0,0,0,90,0,0,0,200,0,92,0,105,0,252,0,154,0,166,0,20,0,62,0,160,0,249,0,170,0,74,0,243,0,99,0,67,0,211,0,222,0,0,0,150,0,115,0,106,0,213,0,0,0,98,0,66,0,93,0,177,0,214,0,240,0,115,0,0,0,157,0,47,0,234,0,44,0,20,0,165,0,217,0,181,0,187,0,248,0,82,0,0,0,68,0,240,0,0,0,0,0,0,0,173,0,0,0,0,0,241,0,52,0,173,0,138,0,213,0,0,0,44,0,0,0,0,0,137,0,184,0,0,0,191,0,170,0,75,0,58,0,196,0,156,0,138,0,0,0,80,0,0,0,203,0,0,0,75,0,25,0,202,0,17,0,101,0,26,0,15,0,20,0,0,0,120,0,147,0,80,0,161,0,169,0,244,0,88,0,255,0,121,0,0,0,139,0,109,0,20,0,11,0,215,0,0,0,0,0,167,0,135,0,99,0,135,0,168,0,134,0,254,0,227,0,252,0,118,0,0,0,91,0,222,0,0,0,239,0,65,0,0,0,244,0,215,0,165,0,207,0,152,0,49,0,128,0,63,0,192,0,255,0,153,0,176,0,43,0,139,0,179,0,86,0,0,0,14,0,233,0,186,0,43,0,190,0,228,0,31,0,0,0,109,0,175,0,239,0,100,0,150,0,186,0,131,0,144,0,205,0,0,0,163,0,0,0,125,0,235,0,153,0,0,0,34,0,0,0,20,0,20,0,90,0,246,0,62,0,253,0,0,0,158,0,160,0,137,0,240,0,13,0,28,0,100,0,163,0,4,0,166,0,0,0,206,0,183,0,113,0,25,0,119,0,117,0,0,0,0,0,27,0,184,0,203,0,143,0,109,0,95,0,8,0,183,0,103,0,224,0,71,0,5,0,217,0,24,0,237,0,0,0,247,0,0,0,0,0,113,0,215,0,237,0,33,0,180,0,59,0,115,0,7,0,209,0,35,0,210,0,0,0,0,0,52,0,0,0,0,0,39,0,31,0,89,0,0,0,191,0,213,0,51,0,130,0,2,0,142,0,226,0,192,0,73,0,133,0,5,0,28,0,39,0,35,0,0,0,45,0,66,0,111,0,102,0,0,0,145,0,177,0,39,0,254,0,0,0,184,0,122,0,168,0,80,0,147,0,29,0,168,0,0,0,27,0,0,0,221,0,195,0,0,0,198,0,83,0,211,0,161,0,141,0,75,0,136,0,0,0,156,0,130,0,0,0,154,0,232,0,100,0,43,0,158,0,172,0,10,0,0,0,36,0,124,0,229,0,0,0,40,0,113,0,2,0,0,0,172,0,30,0,100,0,186,0,81,0,196,0,181,0,180,0,164,0,87,0,65,0,136,0,0,0,148,0,175,0,7,0,0,0,194,0,1,0,0,0,164,0,241,0,212,0,58,0,147,0,0,0,118,0,0,0,134,0,90,0,102,0,87,0,0,0,0,0,0,0,0,0,135,0,77,0,81,0,0,0,6,0,224,0,31,0,0,0,75,0,179,0,0,0,180,0,160,0,48,0,46,0,0,0,160,0,0,0,144,0,60,0,104,0,0,0,0,0,0,0,150,0,0,0,204,0,163,0,175,0,0,0,0,0,0,0,79,0,134,0,75,0,0,0,145,0,239,0,56,0,153,0,0,0,0,0,121,0,210,0,155,0,203,0,168,0,21,0,190,0,217,0,46,0,0,0,0,0,9,0,189,0,0,0,32,0,231,0,149,0,2,0,53,0,68,0,130,0,3,0,231,0,74,0,200,0,0,0,137,0,182,0,0,0,48,0,3,0,247,0,62,0,134,0,220,0,32,0,0,0,132,0,2,0,0,0,21,0,98,0,44,0,0,0,0,0,42,0,90,0,117,0,252,0,137,0,0,0,0,0,131,0,21,0,0,0,0,0,0,0,0,0,0,0,218,0,215,0,230,0,134,0,252,0,211,0,131,0,159,0,0,0,0,0,194,0,97,0,33,0,85,0,48,0,244,0,57,0,143,0,0,0,0,0,150,0,58,0,0,0,0,0,0,0,62,0,42,0,179,0,219,0,0,0,207,0,29,0,0,0,192,0,0,0,0,0,33,0,0,0,106,0,118,0,37,0,98,0,180,0,0,0,0,0,173,0,87,0,159,0,75,0,9,0,158,0,0,0,92,0,61,0,37,0,0,0,0,0,0,0,0,0,89,0,209,0,216,0,141,0,89,0,85,0,0,0,0,0,185,0,178,0,39,0,228,0,116,0,0,0,80,0,98,0,214,0,178,0,0,0,228,0,99,0,227,0,219,0,186,0,132,0,0,0,62,0,0,0,0,0,190,0,0,0,11,0,78,0,102,0,144,0,78,0,250,0,76,0,49,0,182,0,0,0,76,0,145,0,195,0,242,0,180,0,0,0,0,0,113,0,28,0,115,0,32,0,202,0,47,0,193,0,0,0,123,0,199,0,49,0,11,0,94,0,247,0,217,0,53,0,6,0,0,0,193,0,84,0,73,0,0,0,227,0,191,0,202,0,0,0,204,0,39,0,2,0,95,0,142,0,79,0,158,0,240,0,130,0,0,0,57,0,38,0,157,0,23,0,130,0,60,0,128,0,0,0,201,0,3,0,142,0,0,0,247,0,222,0,68,0,0,0,0,0,58,0,27,0,187,0,229,0,165,0,184,0,199,0,242,0,41,0,146,0,40,0,79,0,0,0,35,0,253,0,212,0,33,0,53,0,187,0,119,0,218,0,114,0,92,0,2,0,97,0,0,0,0,0,163,0,0,0,97,0,248,0,0,0,57,0,208,0,51,0,184,0,153,0,97,0,56,0,8,0,240,0,201,0,0,0,247,0,0,0,215,0,103,0,16,0,61,0,196,0,98,0,0,0,191,0,145,0,202,0,73,0,203,0,130,0,155,0,138,0,0,0,0,0,183,0,134,0,142,0,23,0,99,0,123,0,0,0,0,0,242,0,173,0,19,0,126,0,215,0,84,0,70,0,159,0,26,0,58,0,54,0,37,0,105,0,231,0,183,0,117,0,159,0,163,0,163,0,217,0,0,0,196,0,139,0,0,0,15,0,227,0,232,0,217,0,0,0,56,0,134,0,219,0,239,0,221,0,150,0,53,0,100,0,98,0,0,0,68,0,144,0,133,0,88,0,100,0,0,0,38,0,108,0,194,0,0,0,16,0,250,0,0,0,16,0,176,0,235,0,105,0,109,0,0,0,232,0,77,0,2,0,121,0,52,0,64,0,0,0,180,0,0,0,204,0,160,0,0,0,92,0,107,0,81,0,0,0,193,0,88,0,0,0,48,0,98,0,37,0,189,0,245,0,0,0,53,0,28,0,0,0,35,0,179,0,157,0,0,0,179,0,181,0,109,0,97,0,141,0,189,0);
signal scenario_full  : scenario_type := (156,31,156,30,24,31,111,31,239,31,239,30,159,31,140,31,153,31,122,31,149,31,223,31,223,30,223,29,217,31,217,30,165,31,12,31,12,30,59,31,198,31,198,30,198,29,140,31,140,30,133,31,25,31,25,30,205,31,136,31,140,31,24,31,61,31,200,31,52,31,191,31,114,31,231,31,37,31,59,31,15,31,58,31,13,31,78,31,56,31,56,30,45,31,191,31,164,31,253,31,253,30,150,31,69,31,247,31,247,30,36,31,171,31,171,30,171,29,47,31,47,30,182,31,144,31,4,31,19,31,112,31,11,31,211,31,32,31,124,31,100,31,200,31,52,31,23,31,182,31,209,31,211,31,136,31,136,30,242,31,252,31,223,31,223,30,223,29,250,31,218,31,133,31,165,31,61,31,254,31,88,31,153,31,153,30,128,31,66,31,28,31,28,30,28,29,127,31,235,31,109,31,147,31,46,31,164,31,132,31,242,31,52,31,69,31,148,31,245,31,149,31,105,31,88,31,179,31,108,31,108,30,108,29,198,31,4,31,118,31,118,30,160,31,249,31,127,31,230,31,230,30,230,29,18,31,121,31,143,31,115,31,22,31,166,31,166,30,111,31,111,30,155,31,155,30,155,29,226,31,226,30,68,31,93,31,36,31,176,31,176,30,115,31,184,31,169,31,187,31,187,30,187,29,119,31,119,30,155,31,228,31,158,31,231,31,12,31,250,31,165,31,165,30,19,31,206,31,175,31,175,30,166,31,134,31,134,30,134,29,188,31,67,31,133,31,40,31,99,31,84,31,84,30,35,31,249,31,244,31,22,31,71,31,71,30,32,31,255,31,39,31,99,31,64,31,93,31,91,31,227,31,227,30,54,31,15,31,78,31,99,31,119,31,146,31,174,31,174,30,49,31,165,31,222,31,222,31,207,31,213,31,162,31,44,31,46,31,163,31,163,30,207,31,101,31,12,31,218,31,68,31,111,31,156,31,18,31,153,31,254,31,132,31,213,31,76,31,96,31,66,31,153,31,153,30,216,31,161,31,206,31,101,31,82,31,82,30,108,31,141,31,244,31,136,31,124,31,59,31,59,30,80,31,216,31,158,31,93,31,205,31,205,30,188,31,113,31,113,30,251,31,40,31,59,31,247,31,144,31,243,31,132,31,132,30,90,31,90,30,200,31,92,31,105,31,252,31,154,31,166,31,20,31,62,31,160,31,249,31,170,31,74,31,243,31,99,31,67,31,211,31,222,31,222,30,150,31,115,31,106,31,213,31,213,30,98,31,66,31,93,31,177,31,214,31,240,31,115,31,115,30,157,31,47,31,234,31,44,31,20,31,165,31,217,31,181,31,187,31,248,31,82,31,82,30,68,31,240,31,240,30,240,29,240,28,173,31,173,30,173,29,241,31,52,31,173,31,138,31,213,31,213,30,44,31,44,30,44,29,137,31,184,31,184,30,191,31,170,31,75,31,58,31,196,31,156,31,138,31,138,30,80,31,80,30,203,31,203,30,75,31,25,31,202,31,17,31,101,31,26,31,15,31,20,31,20,30,120,31,147,31,80,31,161,31,169,31,244,31,88,31,255,31,121,31,121,30,139,31,109,31,20,31,11,31,215,31,215,30,215,29,167,31,135,31,99,31,135,31,168,31,134,31,254,31,227,31,252,31,118,31,118,30,91,31,222,31,222,30,239,31,65,31,65,30,244,31,215,31,165,31,207,31,152,31,49,31,128,31,63,31,192,31,255,31,153,31,176,31,43,31,139,31,179,31,86,31,86,30,14,31,233,31,186,31,43,31,190,31,228,31,31,31,31,30,109,31,175,31,239,31,100,31,150,31,186,31,131,31,144,31,205,31,205,30,163,31,163,30,125,31,235,31,153,31,153,30,34,31,34,30,20,31,20,31,90,31,246,31,62,31,253,31,253,30,158,31,160,31,137,31,240,31,13,31,28,31,100,31,163,31,4,31,166,31,166,30,206,31,183,31,113,31,25,31,119,31,117,31,117,30,117,29,27,31,184,31,203,31,143,31,109,31,95,31,8,31,183,31,103,31,224,31,71,31,5,31,217,31,24,31,237,31,237,30,247,31,247,30,247,29,113,31,215,31,237,31,33,31,180,31,59,31,115,31,7,31,209,31,35,31,210,31,210,30,210,29,52,31,52,30,52,29,39,31,31,31,89,31,89,30,191,31,213,31,51,31,130,31,2,31,142,31,226,31,192,31,73,31,133,31,5,31,28,31,39,31,35,31,35,30,45,31,66,31,111,31,102,31,102,30,145,31,177,31,39,31,254,31,254,30,184,31,122,31,168,31,80,31,147,31,29,31,168,31,168,30,27,31,27,30,221,31,195,31,195,30,198,31,83,31,211,31,161,31,141,31,75,31,136,31,136,30,156,31,130,31,130,30,154,31,232,31,100,31,43,31,158,31,172,31,10,31,10,30,36,31,124,31,229,31,229,30,40,31,113,31,2,31,2,30,172,31,30,31,100,31,186,31,81,31,196,31,181,31,180,31,164,31,87,31,65,31,136,31,136,30,148,31,175,31,7,31,7,30,194,31,1,31,1,30,164,31,241,31,212,31,58,31,147,31,147,30,118,31,118,30,134,31,90,31,102,31,87,31,87,30,87,29,87,28,87,27,135,31,77,31,81,31,81,30,6,31,224,31,31,31,31,30,75,31,179,31,179,30,180,31,160,31,48,31,46,31,46,30,160,31,160,30,144,31,60,31,104,31,104,30,104,29,104,28,150,31,150,30,204,31,163,31,175,31,175,30,175,29,175,28,79,31,134,31,75,31,75,30,145,31,239,31,56,31,153,31,153,30,153,29,121,31,210,31,155,31,203,31,168,31,21,31,190,31,217,31,46,31,46,30,46,29,9,31,189,31,189,30,32,31,231,31,149,31,2,31,53,31,68,31,130,31,3,31,231,31,74,31,200,31,200,30,137,31,182,31,182,30,48,31,3,31,247,31,62,31,134,31,220,31,32,31,32,30,132,31,2,31,2,30,21,31,98,31,44,31,44,30,44,29,42,31,90,31,117,31,252,31,137,31,137,30,137,29,131,31,21,31,21,30,21,29,21,28,21,27,21,26,218,31,215,31,230,31,134,31,252,31,211,31,131,31,159,31,159,30,159,29,194,31,97,31,33,31,85,31,48,31,244,31,57,31,143,31,143,30,143,29,150,31,58,31,58,30,58,29,58,28,62,31,42,31,179,31,219,31,219,30,207,31,29,31,29,30,192,31,192,30,192,29,33,31,33,30,106,31,118,31,37,31,98,31,180,31,180,30,180,29,173,31,87,31,159,31,75,31,9,31,158,31,158,30,92,31,61,31,37,31,37,30,37,29,37,28,37,27,89,31,209,31,216,31,141,31,89,31,85,31,85,30,85,29,185,31,178,31,39,31,228,31,116,31,116,30,80,31,98,31,214,31,178,31,178,30,228,31,99,31,227,31,219,31,186,31,132,31,132,30,62,31,62,30,62,29,190,31,190,30,11,31,78,31,102,31,144,31,78,31,250,31,76,31,49,31,182,31,182,30,76,31,145,31,195,31,242,31,180,31,180,30,180,29,113,31,28,31,115,31,32,31,202,31,47,31,193,31,193,30,123,31,199,31,49,31,11,31,94,31,247,31,217,31,53,31,6,31,6,30,193,31,84,31,73,31,73,30,227,31,191,31,202,31,202,30,204,31,39,31,2,31,95,31,142,31,79,31,158,31,240,31,130,31,130,30,57,31,38,31,157,31,23,31,130,31,60,31,128,31,128,30,201,31,3,31,142,31,142,30,247,31,222,31,68,31,68,30,68,29,58,31,27,31,187,31,229,31,165,31,184,31,199,31,242,31,41,31,146,31,40,31,79,31,79,30,35,31,253,31,212,31,33,31,53,31,187,31,119,31,218,31,114,31,92,31,2,31,97,31,97,30,97,29,163,31,163,30,97,31,248,31,248,30,57,31,208,31,51,31,184,31,153,31,97,31,56,31,8,31,240,31,201,31,201,30,247,31,247,30,215,31,103,31,16,31,61,31,196,31,98,31,98,30,191,31,145,31,202,31,73,31,203,31,130,31,155,31,138,31,138,30,138,29,183,31,134,31,142,31,23,31,99,31,123,31,123,30,123,29,242,31,173,31,19,31,126,31,215,31,84,31,70,31,159,31,26,31,58,31,54,31,37,31,105,31,231,31,183,31,117,31,159,31,163,31,163,31,217,31,217,30,196,31,139,31,139,30,15,31,227,31,232,31,217,31,217,30,56,31,134,31,219,31,239,31,221,31,150,31,53,31,100,31,98,31,98,30,68,31,144,31,133,31,88,31,100,31,100,30,38,31,108,31,194,31,194,30,16,31,250,31,250,30,16,31,176,31,235,31,105,31,109,31,109,30,232,31,77,31,2,31,121,31,52,31,64,31,64,30,180,31,180,30,204,31,160,31,160,30,92,31,107,31,81,31,81,30,193,31,88,31,88,30,48,31,98,31,37,31,189,31,245,31,245,30,53,31,28,31,28,30,35,31,179,31,157,31,157,30,179,31,181,31,109,31,97,31,141,31,189,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
