-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 392;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (160,0,168,0,0,0,174,0,0,0,130,0,36,0,79,0,110,0,82,0,0,0,46,0,133,0,133,0,236,0,166,0,150,0,0,0,87,0,68,0,56,0,97,0,208,0,133,0,132,0,17,0,0,0,255,0,103,0,252,0,219,0,0,0,10,0,102,0,0,0,14,0,200,0,5,0,41,0,204,0,0,0,0,0,123,0,185,0,85,0,190,0,194,0,0,0,37,0,101,0,229,0,0,0,0,0,83,0,196,0,0,0,19,0,241,0,193,0,125,0,0,0,0,0,98,0,0,0,99,0,228,0,94,0,186,0,85,0,0,0,4,0,0,0,167,0,67,0,92,0,0,0,176,0,238,0,206,0,86,0,198,0,151,0,240,0,250,0,38,0,144,0,51,0,113,0,0,0,65,0,70,0,11,0,191,0,204,0,107,0,89,0,253,0,185,0,161,0,62,0,84,0,0,0,10,0,78,0,0,0,0,0,146,0,60,0,37,0,39,0,0,0,0,0,27,0,146,0,100,0,0,0,23,0,0,0,64,0,0,0,27,0,73,0,0,0,57,0,165,0,139,0,66,0,148,0,51,0,0,0,196,0,79,0,72,0,188,0,194,0,238,0,186,0,218,0,201,0,9,0,0,0,241,0,73,0,205,0,244,0,0,0,178,0,0,0,93,0,0,0,0,0,0,0,0,0,60,0,100,0,0,0,138,0,164,0,162,0,141,0,127,0,125,0,131,0,22,0,80,0,245,0,224,0,65,0,0,0,56,0,6,0,115,0,75,0,134,0,0,0,248,0,207,0,91,0,28,0,237,0,214,0,128,0,110,0,80,0,237,0,0,0,160,0,0,0,155,0,84,0,55,0,198,0,208,0,0,0,206,0,185,0,0,0,85,0,183,0,0,0,248,0,16,0,41,0,101,0,80,0,224,0,71,0,156,0,229,0,52,0,165,0,184,0,102,0,227,0,193,0,162,0,128,0,130,0,189,0,26,0,207,0,4,0,235,0,20,0,0,0,99,0,106,0,226,0,33,0,0,0,213,0,133,0,0,0,0,0,0,0,5,0,61,0,219,0,238,0,80,0,0,0,0,0,212,0,16,0,145,0,86,0,0,0,27,0,1,0,206,0,17,0,163,0,179,0,0,0,139,0,204,0,0,0,0,0,95,0,128,0,231,0,51,0,215,0,71,0,0,0,201,0,185,0,215,0,19,0,42,0,58,0,0,0,81,0,81,0,0,0,17,0,71,0,18,0,146,0,190,0,0,0,0,0,0,0,0,0,15,0,45,0,213,0,254,0,238,0,52,0,192,0,0,0,202,0,0,0,105,0,32,0,0,0,230,0,0,0,141,0,189,0,246,0,189,0,198,0,35,0,44,0,0,0,0,0,153,0,0,0,0,0,77,0,103,0,221,0,130,0,0,0,227,0,246,0,0,0,163,0,50,0,101,0,20,0,213,0,122,0,89,0,245,0,9,0,181,0,101,0,59,0,171,0,0,0,119,0,89,0,0,0,0,0,212,0,198,0,187,0,0,0,0,0,159,0,97,0,0,0,0,0,47,0,165,0,202,0,76,0,165,0,131,0,187,0,71,0,0,0,46,0,141,0,189,0,209,0,163,0,0,0,0,0,169,0,129,0,231,0,88,0,221,0,0,0,233,0,92,0,0,0,183,0,0,0,20,0,252,0,175,0,195,0,241,0,133,0,47,0,59,0,0,0,144,0,238,0,87,0,0,0,0,0,107,0,38,0,148,0,0,0,182,0);
signal scenario_full  : scenario_type := (160,31,168,31,168,30,174,31,174,30,130,31,36,31,79,31,110,31,82,31,82,30,46,31,133,31,133,31,236,31,166,31,150,31,150,30,87,31,68,31,56,31,97,31,208,31,133,31,132,31,17,31,17,30,255,31,103,31,252,31,219,31,219,30,10,31,102,31,102,30,14,31,200,31,5,31,41,31,204,31,204,30,204,29,123,31,185,31,85,31,190,31,194,31,194,30,37,31,101,31,229,31,229,30,229,29,83,31,196,31,196,30,19,31,241,31,193,31,125,31,125,30,125,29,98,31,98,30,99,31,228,31,94,31,186,31,85,31,85,30,4,31,4,30,167,31,67,31,92,31,92,30,176,31,238,31,206,31,86,31,198,31,151,31,240,31,250,31,38,31,144,31,51,31,113,31,113,30,65,31,70,31,11,31,191,31,204,31,107,31,89,31,253,31,185,31,161,31,62,31,84,31,84,30,10,31,78,31,78,30,78,29,146,31,60,31,37,31,39,31,39,30,39,29,27,31,146,31,100,31,100,30,23,31,23,30,64,31,64,30,27,31,73,31,73,30,57,31,165,31,139,31,66,31,148,31,51,31,51,30,196,31,79,31,72,31,188,31,194,31,238,31,186,31,218,31,201,31,9,31,9,30,241,31,73,31,205,31,244,31,244,30,178,31,178,30,93,31,93,30,93,29,93,28,93,27,60,31,100,31,100,30,138,31,164,31,162,31,141,31,127,31,125,31,131,31,22,31,80,31,245,31,224,31,65,31,65,30,56,31,6,31,115,31,75,31,134,31,134,30,248,31,207,31,91,31,28,31,237,31,214,31,128,31,110,31,80,31,237,31,237,30,160,31,160,30,155,31,84,31,55,31,198,31,208,31,208,30,206,31,185,31,185,30,85,31,183,31,183,30,248,31,16,31,41,31,101,31,80,31,224,31,71,31,156,31,229,31,52,31,165,31,184,31,102,31,227,31,193,31,162,31,128,31,130,31,189,31,26,31,207,31,4,31,235,31,20,31,20,30,99,31,106,31,226,31,33,31,33,30,213,31,133,31,133,30,133,29,133,28,5,31,61,31,219,31,238,31,80,31,80,30,80,29,212,31,16,31,145,31,86,31,86,30,27,31,1,31,206,31,17,31,163,31,179,31,179,30,139,31,204,31,204,30,204,29,95,31,128,31,231,31,51,31,215,31,71,31,71,30,201,31,185,31,215,31,19,31,42,31,58,31,58,30,81,31,81,31,81,30,17,31,71,31,18,31,146,31,190,31,190,30,190,29,190,28,190,27,15,31,45,31,213,31,254,31,238,31,52,31,192,31,192,30,202,31,202,30,105,31,32,31,32,30,230,31,230,30,141,31,189,31,246,31,189,31,198,31,35,31,44,31,44,30,44,29,153,31,153,30,153,29,77,31,103,31,221,31,130,31,130,30,227,31,246,31,246,30,163,31,50,31,101,31,20,31,213,31,122,31,89,31,245,31,9,31,181,31,101,31,59,31,171,31,171,30,119,31,89,31,89,30,89,29,212,31,198,31,187,31,187,30,187,29,159,31,97,31,97,30,97,29,47,31,165,31,202,31,76,31,165,31,131,31,187,31,71,31,71,30,46,31,141,31,189,31,209,31,163,31,163,30,163,29,169,31,129,31,231,31,88,31,221,31,221,30,233,31,92,31,92,30,183,31,183,30,20,31,252,31,175,31,195,31,241,31,133,31,47,31,59,31,59,30,144,31,238,31,87,31,87,30,87,29,107,31,38,31,148,31,148,30,182,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
