-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 676;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (181,0,0,0,76,0,42,0,44,0,42,0,42,0,228,0,0,0,96,0,7,0,69,0,234,0,0,0,54,0,212,0,200,0,134,0,67,0,138,0,0,0,26,0,0,0,236,0,48,0,150,0,0,0,90,0,0,0,203,0,205,0,220,0,56,0,0,0,127,0,0,0,0,0,214,0,0,0,53,0,28,0,33,0,37,0,216,0,14,0,193,0,81,0,31,0,142,0,66,0,0,0,123,0,192,0,21,0,39,0,230,0,17,0,219,0,3,0,0,0,180,0,83,0,44,0,128,0,103,0,181,0,201,0,116,0,157,0,191,0,0,0,91,0,217,0,248,0,146,0,126,0,237,0,188,0,47,0,179,0,250,0,36,0,0,0,92,0,27,0,0,0,225,0,150,0,144,0,0,0,66,0,32,0,158,0,0,0,15,0,151,0,0,0,47,0,153,0,25,0,96,0,255,0,0,0,110,0,94,0,157,0,69,0,0,0,32,0,120,0,143,0,248,0,24,0,90,0,144,0,165,0,55,0,20,0,114,0,201,0,37,0,51,0,194,0,32,0,199,0,0,0,21,0,1,0,49,0,145,0,0,0,108,0,13,0,124,0,3,0,44,0,0,0,52,0,78,0,61,0,0,0,123,0,150,0,127,0,236,0,76,0,13,0,104,0,214,0,243,0,158,0,250,0,12,0,171,0,112,0,61,0,193,0,117,0,154,0,0,0,144,0,0,0,26,0,163,0,190,0,27,0,16,0,244,0,0,0,108,0,35,0,176,0,0,0,245,0,17,0,82,0,159,0,0,0,0,0,0,0,0,0,114,0,0,0,0,0,219,0,6,0,184,0,0,0,13,0,52,0,195,0,48,0,82,0,0,0,232,0,245,0,76,0,64,0,239,0,210,0,201,0,0,0,245,0,11,0,102,0,0,0,127,0,254,0,237,0,16,0,0,0,50,0,50,0,232,0,0,0,21,0,140,0,0,0,205,0,94,0,209,0,139,0,94,0,245,0,11,0,0,0,0,0,32,0,202,0,146,0,172,0,35,0,214,0,137,0,74,0,0,0,169,0,242,0,65,0,249,0,55,0,218,0,0,0,60,0,100,0,196,0,169,0,0,0,118,0,195,0,76,0,217,0,189,0,243,0,218,0,248,0,152,0,255,0,212,0,0,0,2,0,63,0,145,0,64,0,0,0,208,0,13,0,76,0,26,0,83,0,0,0,0,0,8,0,46,0,58,0,181,0,31,0,10,0,73,0,37,0,0,0,18,0,15,0,27,0,22,0,206,0,66,0,110,0,0,0,0,0,0,0,241,0,0,0,16,0,144,0,0,0,224,0,212,0,0,0,174,0,184,0,0,0,77,0,29,0,96,0,0,0,0,0,0,0,147,0,156,0,182,0,217,0,230,0,235,0,120,0,91,0,198,0,141,0,0,0,43,0,137,0,4,0,148,0,119,0,0,0,57,0,9,0,127,0,222,0,40,0,212,0,150,0,233,0,13,0,0,0,137,0,88,0,176,0,128,0,0,0,0,0,0,0,233,0,123,0,28,0,176,0,0,0,67,0,0,0,0,0,16,0,37,0,246,0,0,0,182,0,117,0,11,0,251,0,187,0,83,0,104,0,4,0,174,0,143,0,112,0,10,0,235,0,53,0,0,0,159,0,0,0,183,0,0,0,0,0,55,0,0,0,0,0,25,0,63,0,162,0,68,0,191,0,45,0,0,0,148,0,34,0,0,0,238,0,101,0,159,0,0,0,152,0,29,0,58,0,148,0,0,0,153,0,95,0,0,0,102,0,0,0,0,0,168,0,19,0,0,0,242,0,71,0,231,0,151,0,0,0,129,0,216,0,181,0,149,0,76,0,4,0,82,0,52,0,7,0,179,0,194,0,108,0,0,0,125,0,0,0,69,0,6,0,0,0,105,0,123,0,253,0,57,0,175,0,176,0,0,0,172,0,254,0,47,0,137,0,16,0,217,0,0,0,0,0,0,0,0,0,31,0,111,0,244,0,134,0,221,0,0,0,83,0,250,0,70,0,140,0,0,0,21,0,182,0,135,0,112,0,156,0,57,0,255,0,175,0,0,0,237,0,28,0,162,0,208,0,175,0,193,0,0,0,208,0,0,0,75,0,204,0,80,0,227,0,0,0,21,0,76,0,83,0,74,0,20,0,147,0,0,0,0,0,126,0,0,0,185,0,13,0,25,0,179,0,131,0,19,0,0,0,0,0,107,0,0,0,234,0,125,0,5,0,51,0,0,0,0,0,0,0,84,0,125,0,247,0,0,0,200,0,144,0,64,0,207,0,168,0,0,0,25,0,100,0,0,0,229,0,88,0,232,0,0,0,0,0,239,0,68,0,82,0,75,0,95,0,213,0,0,0,99,0,74,0,4,0,128,0,117,0,57,0,217,0,147,0,0,0,247,0,108,0,244,0,208,0,12,0,242,0,242,0,144,0,191,0,107,0,7,0,248,0,250,0,216,0,43,0,114,0,0,0,156,0,66,0,16,0,94,0,211,0,114,0,211,0,144,0,249,0,212,0,228,0,72,0,173,0,0,0,4,0,188,0,0,0,157,0,121,0,178,0,122,0,0,0,252,0,2,0,212,0,176,0,0,0,17,0,155,0,0,0,130,0,242,0,57,0,83,0,157,0,127,0,77,0,234,0,108,0,16,0,28,0,206,0,0,0,0,0,145,0,183,0,0,0,98,0,0,0,0,0,0,0,0,0,122,0,166,0,213,0,239,0,222,0,244,0,63,0,120,0,231,0,196,0,54,0,0,0,70,0,239,0,236,0,147,0,63,0,0,0,0,0,0,0,110,0,104,0,180,0,228,0,154,0,7,0,183,0,105,0,114,0,0,0,142,0,247,0,0,0,134,0,243,0,182,0,74,0,80,0,60,0,32,0,137,0,0,0,250,0,207,0,0,0,186,0,242,0,196,0,0,0,0,0,81,0,171,0,0,0,157,0,177,0,15,0,122,0,49,0,0,0,36,0,36,0,168,0,109,0,221,0,92,0,184,0,228,0);
signal scenario_full  : scenario_type := (181,31,181,30,76,31,42,31,44,31,42,31,42,31,228,31,228,30,96,31,7,31,69,31,234,31,234,30,54,31,212,31,200,31,134,31,67,31,138,31,138,30,26,31,26,30,236,31,48,31,150,31,150,30,90,31,90,30,203,31,205,31,220,31,56,31,56,30,127,31,127,30,127,29,214,31,214,30,53,31,28,31,33,31,37,31,216,31,14,31,193,31,81,31,31,31,142,31,66,31,66,30,123,31,192,31,21,31,39,31,230,31,17,31,219,31,3,31,3,30,180,31,83,31,44,31,128,31,103,31,181,31,201,31,116,31,157,31,191,31,191,30,91,31,217,31,248,31,146,31,126,31,237,31,188,31,47,31,179,31,250,31,36,31,36,30,92,31,27,31,27,30,225,31,150,31,144,31,144,30,66,31,32,31,158,31,158,30,15,31,151,31,151,30,47,31,153,31,25,31,96,31,255,31,255,30,110,31,94,31,157,31,69,31,69,30,32,31,120,31,143,31,248,31,24,31,90,31,144,31,165,31,55,31,20,31,114,31,201,31,37,31,51,31,194,31,32,31,199,31,199,30,21,31,1,31,49,31,145,31,145,30,108,31,13,31,124,31,3,31,44,31,44,30,52,31,78,31,61,31,61,30,123,31,150,31,127,31,236,31,76,31,13,31,104,31,214,31,243,31,158,31,250,31,12,31,171,31,112,31,61,31,193,31,117,31,154,31,154,30,144,31,144,30,26,31,163,31,190,31,27,31,16,31,244,31,244,30,108,31,35,31,176,31,176,30,245,31,17,31,82,31,159,31,159,30,159,29,159,28,159,27,114,31,114,30,114,29,219,31,6,31,184,31,184,30,13,31,52,31,195,31,48,31,82,31,82,30,232,31,245,31,76,31,64,31,239,31,210,31,201,31,201,30,245,31,11,31,102,31,102,30,127,31,254,31,237,31,16,31,16,30,50,31,50,31,232,31,232,30,21,31,140,31,140,30,205,31,94,31,209,31,139,31,94,31,245,31,11,31,11,30,11,29,32,31,202,31,146,31,172,31,35,31,214,31,137,31,74,31,74,30,169,31,242,31,65,31,249,31,55,31,218,31,218,30,60,31,100,31,196,31,169,31,169,30,118,31,195,31,76,31,217,31,189,31,243,31,218,31,248,31,152,31,255,31,212,31,212,30,2,31,63,31,145,31,64,31,64,30,208,31,13,31,76,31,26,31,83,31,83,30,83,29,8,31,46,31,58,31,181,31,31,31,10,31,73,31,37,31,37,30,18,31,15,31,27,31,22,31,206,31,66,31,110,31,110,30,110,29,110,28,241,31,241,30,16,31,144,31,144,30,224,31,212,31,212,30,174,31,184,31,184,30,77,31,29,31,96,31,96,30,96,29,96,28,147,31,156,31,182,31,217,31,230,31,235,31,120,31,91,31,198,31,141,31,141,30,43,31,137,31,4,31,148,31,119,31,119,30,57,31,9,31,127,31,222,31,40,31,212,31,150,31,233,31,13,31,13,30,137,31,88,31,176,31,128,31,128,30,128,29,128,28,233,31,123,31,28,31,176,31,176,30,67,31,67,30,67,29,16,31,37,31,246,31,246,30,182,31,117,31,11,31,251,31,187,31,83,31,104,31,4,31,174,31,143,31,112,31,10,31,235,31,53,31,53,30,159,31,159,30,183,31,183,30,183,29,55,31,55,30,55,29,25,31,63,31,162,31,68,31,191,31,45,31,45,30,148,31,34,31,34,30,238,31,101,31,159,31,159,30,152,31,29,31,58,31,148,31,148,30,153,31,95,31,95,30,102,31,102,30,102,29,168,31,19,31,19,30,242,31,71,31,231,31,151,31,151,30,129,31,216,31,181,31,149,31,76,31,4,31,82,31,52,31,7,31,179,31,194,31,108,31,108,30,125,31,125,30,69,31,6,31,6,30,105,31,123,31,253,31,57,31,175,31,176,31,176,30,172,31,254,31,47,31,137,31,16,31,217,31,217,30,217,29,217,28,217,27,31,31,111,31,244,31,134,31,221,31,221,30,83,31,250,31,70,31,140,31,140,30,21,31,182,31,135,31,112,31,156,31,57,31,255,31,175,31,175,30,237,31,28,31,162,31,208,31,175,31,193,31,193,30,208,31,208,30,75,31,204,31,80,31,227,31,227,30,21,31,76,31,83,31,74,31,20,31,147,31,147,30,147,29,126,31,126,30,185,31,13,31,25,31,179,31,131,31,19,31,19,30,19,29,107,31,107,30,234,31,125,31,5,31,51,31,51,30,51,29,51,28,84,31,125,31,247,31,247,30,200,31,144,31,64,31,207,31,168,31,168,30,25,31,100,31,100,30,229,31,88,31,232,31,232,30,232,29,239,31,68,31,82,31,75,31,95,31,213,31,213,30,99,31,74,31,4,31,128,31,117,31,57,31,217,31,147,31,147,30,247,31,108,31,244,31,208,31,12,31,242,31,242,31,144,31,191,31,107,31,7,31,248,31,250,31,216,31,43,31,114,31,114,30,156,31,66,31,16,31,94,31,211,31,114,31,211,31,144,31,249,31,212,31,228,31,72,31,173,31,173,30,4,31,188,31,188,30,157,31,121,31,178,31,122,31,122,30,252,31,2,31,212,31,176,31,176,30,17,31,155,31,155,30,130,31,242,31,57,31,83,31,157,31,127,31,77,31,234,31,108,31,16,31,28,31,206,31,206,30,206,29,145,31,183,31,183,30,98,31,98,30,98,29,98,28,98,27,122,31,166,31,213,31,239,31,222,31,244,31,63,31,120,31,231,31,196,31,54,31,54,30,70,31,239,31,236,31,147,31,63,31,63,30,63,29,63,28,110,31,104,31,180,31,228,31,154,31,7,31,183,31,105,31,114,31,114,30,142,31,247,31,247,30,134,31,243,31,182,31,74,31,80,31,60,31,32,31,137,31,137,30,250,31,207,31,207,30,186,31,242,31,196,31,196,30,196,29,81,31,171,31,171,30,157,31,177,31,15,31,122,31,49,31,49,30,36,31,36,31,168,31,109,31,221,31,92,31,184,31,228,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
