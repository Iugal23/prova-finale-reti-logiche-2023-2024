-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 347;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (200,0,127,0,0,0,34,0,1,0,222,0,32,0,76,0,97,0,24,0,20,0,122,0,95,0,0,0,98,0,0,0,41,0,218,0,113,0,81,0,0,0,116,0,0,0,0,0,204,0,39,0,0,0,0,0,126,0,26,0,163,0,158,0,86,0,0,0,193,0,60,0,0,0,0,0,15,0,7,0,27,0,25,0,177,0,67,0,0,0,0,0,0,0,132,0,132,0,210,0,149,0,0,0,203,0,143,0,187,0,86,0,195,0,226,0,27,0,84,0,142,0,63,0,221,0,0,0,127,0,39,0,195,0,29,0,150,0,0,0,184,0,0,0,104,0,0,0,91,0,232,0,159,0,161,0,0,0,71,0,9,0,40,0,36,0,67,0,118,0,0,0,174,0,126,0,253,0,163,0,249,0,19,0,218,0,33,0,247,0,68,0,248,0,205,0,137,0,202,0,0,0,171,0,74,0,105,0,102,0,235,0,253,0,0,0,209,0,189,0,121,0,185,0,232,0,0,0,78,0,20,0,34,0,175,0,139,0,245,0,0,0,191,0,29,0,84,0,0,0,96,0,49,0,84,0,131,0,137,0,62,0,32,0,54,0,238,0,0,0,0,0,171,0,0,0,65,0,86,0,128,0,25,0,154,0,0,0,110,0,143,0,67,0,114,0,22,0,191,0,54,0,194,0,207,0,183,0,168,0,230,0,95,0,0,0,211,0,0,0,0,0,213,0,0,0,142,0,75,0,0,0,122,0,162,0,203,0,27,0,253,0,1,0,19,0,57,0,0,0,0,0,40,0,0,0,239,0,155,0,49,0,0,0,121,0,81,0,34,0,43,0,113,0,73,0,0,0,7,0,40,0,220,0,156,0,197,0,0,0,129,0,212,0,26,0,245,0,228,0,0,0,133,0,186,0,0,0,0,0,169,0,182,0,0,0,200,0,81,0,0,0,133,0,39,0,186,0,212,0,85,0,17,0,0,0,82,0,57,0,84,0,160,0,166,0,146,0,0,0,139,0,114,0,0,0,0,0,45,0,32,0,197,0,0,0,0,0,54,0,56,0,98,0,11,0,68,0,64,0,0,0,0,0,240,0,0,0,34,0,148,0,45,0,17,0,0,0,79,0,199,0,228,0,0,0,236,0,216,0,108,0,243,0,166,0,0,0,193,0,221,0,114,0,136,0,0,0,160,0,0,0,239,0,0,0,81,0,223,0,0,0,249,0,213,0,113,0,227,0,73,0,0,0,65,0,12,0,0,0,134,0,152,0,249,0,181,0,212,0,0,0,6,0,153,0,88,0,0,0,35,0,208,0,0,0,58,0,68,0,0,0,42,0,0,0,6,0,0,0,248,0,139,0,73,0,125,0,80,0,0,0,87,0,71,0,147,0,16,0,172,0,220,0,23,0,107,0,119,0,25,0,86,0,238,0,164,0,41,0,0,0,252,0,145,0,179,0,0,0,0,0,86,0,30,0,87,0,174,0,186,0,243,0,97,0,114,0,0,0,239,0,0,0,199,0,64,0,184,0,118,0,188,0,225,0,41,0,135,0,161,0,178,0);
signal scenario_full  : scenario_type := (200,31,127,31,127,30,34,31,1,31,222,31,32,31,76,31,97,31,24,31,20,31,122,31,95,31,95,30,98,31,98,30,41,31,218,31,113,31,81,31,81,30,116,31,116,30,116,29,204,31,39,31,39,30,39,29,126,31,26,31,163,31,158,31,86,31,86,30,193,31,60,31,60,30,60,29,15,31,7,31,27,31,25,31,177,31,67,31,67,30,67,29,67,28,132,31,132,31,210,31,149,31,149,30,203,31,143,31,187,31,86,31,195,31,226,31,27,31,84,31,142,31,63,31,221,31,221,30,127,31,39,31,195,31,29,31,150,31,150,30,184,31,184,30,104,31,104,30,91,31,232,31,159,31,161,31,161,30,71,31,9,31,40,31,36,31,67,31,118,31,118,30,174,31,126,31,253,31,163,31,249,31,19,31,218,31,33,31,247,31,68,31,248,31,205,31,137,31,202,31,202,30,171,31,74,31,105,31,102,31,235,31,253,31,253,30,209,31,189,31,121,31,185,31,232,31,232,30,78,31,20,31,34,31,175,31,139,31,245,31,245,30,191,31,29,31,84,31,84,30,96,31,49,31,84,31,131,31,137,31,62,31,32,31,54,31,238,31,238,30,238,29,171,31,171,30,65,31,86,31,128,31,25,31,154,31,154,30,110,31,143,31,67,31,114,31,22,31,191,31,54,31,194,31,207,31,183,31,168,31,230,31,95,31,95,30,211,31,211,30,211,29,213,31,213,30,142,31,75,31,75,30,122,31,162,31,203,31,27,31,253,31,1,31,19,31,57,31,57,30,57,29,40,31,40,30,239,31,155,31,49,31,49,30,121,31,81,31,34,31,43,31,113,31,73,31,73,30,7,31,40,31,220,31,156,31,197,31,197,30,129,31,212,31,26,31,245,31,228,31,228,30,133,31,186,31,186,30,186,29,169,31,182,31,182,30,200,31,81,31,81,30,133,31,39,31,186,31,212,31,85,31,17,31,17,30,82,31,57,31,84,31,160,31,166,31,146,31,146,30,139,31,114,31,114,30,114,29,45,31,32,31,197,31,197,30,197,29,54,31,56,31,98,31,11,31,68,31,64,31,64,30,64,29,240,31,240,30,34,31,148,31,45,31,17,31,17,30,79,31,199,31,228,31,228,30,236,31,216,31,108,31,243,31,166,31,166,30,193,31,221,31,114,31,136,31,136,30,160,31,160,30,239,31,239,30,81,31,223,31,223,30,249,31,213,31,113,31,227,31,73,31,73,30,65,31,12,31,12,30,134,31,152,31,249,31,181,31,212,31,212,30,6,31,153,31,88,31,88,30,35,31,208,31,208,30,58,31,68,31,68,30,42,31,42,30,6,31,6,30,248,31,139,31,73,31,125,31,80,31,80,30,87,31,71,31,147,31,16,31,172,31,220,31,23,31,107,31,119,31,25,31,86,31,238,31,164,31,41,31,41,30,252,31,145,31,179,31,179,30,179,29,86,31,30,31,87,31,174,31,186,31,243,31,97,31,114,31,114,30,239,31,239,30,199,31,64,31,184,31,118,31,188,31,225,31,41,31,135,31,161,31,178,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
