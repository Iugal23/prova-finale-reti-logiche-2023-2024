-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_227 is
end project_tb_227;

architecture project_tb_arch_227 of project_tb_227 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 681;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (159,0,98,0,144,0,248,0,203,0,0,0,255,0,208,0,248,0,201,0,7,0,0,0,0,0,204,0,136,0,0,0,235,0,229,0,9,0,39,0,182,0,0,0,26,0,0,0,0,0,0,0,65,0,0,0,97,0,4,0,51,0,81,0,86,0,0,0,200,0,250,0,252,0,33,0,161,0,25,0,149,0,199,0,43,0,0,0,0,0,171,0,78,0,0,0,0,0,0,0,109,0,120,0,0,0,151,0,34,0,0,0,230,0,0,0,0,0,0,0,102,0,16,0,0,0,100,0,165,0,40,0,0,0,0,0,0,0,112,0,103,0,165,0,69,0,142,0,192,0,203,0,187,0,168,0,191,0,1,0,50,0,129,0,0,0,12,0,168,0,0,0,55,0,0,0,135,0,3,0,132,0,54,0,81,0,0,0,203,0,247,0,80,0,202,0,86,0,83,0,225,0,0,0,78,0,215,0,182,0,51,0,0,0,54,0,96,0,0,0,149,0,0,0,99,0,39,0,0,0,134,0,91,0,0,0,166,0,244,0,234,0,0,0,0,0,239,0,252,0,19,0,0,0,177,0,198,0,107,0,61,0,0,0,211,0,180,0,31,0,72,0,97,0,0,0,83,0,125,0,124,0,199,0,18,0,76,0,0,0,0,0,80,0,15,0,151,0,120,0,0,0,146,0,0,0,105,0,48,0,0,0,134,0,231,0,0,0,70,0,0,0,129,0,77,0,142,0,29,0,38,0,18,0,40,0,7,0,0,0,0,0,214,0,94,0,0,0,90,0,0,0,0,0,0,0,161,0,111,0,0,0,194,0,169,0,37,0,34,0,54,0,158,0,195,0,10,0,0,0,191,0,0,0,52,0,153,0,33,0,0,0,21,0,161,0,19,0,168,0,43,0,180,0,221,0,12,0,175,0,0,0,147,0,95,0,0,0,92,0,115,0,0,0,136,0,176,0,122,0,160,0,51,0,38,0,140,0,159,0,255,0,40,0,170,0,70,0,82,0,0,0,69,0,52,0,99,0,197,0,18,0,33,0,0,0,2,0,196,0,0,0,0,0,117,0,0,0,103,0,98,0,29,0,123,0,246,0,168,0,140,0,44,0,218,0,144,0,0,0,174,0,208,0,22,0,222,0,14,0,205,0,175,0,20,0,72,0,88,0,211,0,101,0,243,0,180,0,249,0,23,0,35,0,42,0,42,0,6,0,178,0,155,0,109,0,144,0,222,0,129,0,7,0,95,0,41,0,80,0,58,0,16,0,0,0,71,0,251,0,0,0,101,0,132,0,149,0,127,0,20,0,247,0,6,0,85,0,159,0,128,0,186,0,55,0,62,0,179,0,86,0,188,0,42,0,132,0,56,0,208,0,146,0,158,0,172,0,245,0,115,0,26,0,38,0,248,0,229,0,15,0,101,0,12,0,30,0,133,0,249,0,0,0,24,0,22,0,14,0,180,0,41,0,177,0,240,0,138,0,197,0,249,0,215,0,151,0,158,0,106,0,118,0,155,0,129,0,0,0,87,0,133,0,0,0,46,0,246,0,35,0,171,0,0,0,246,0,170,0,209,0,115,0,114,0,91,0,153,0,90,0,102,0,220,0,0,0,101,0,0,0,23,0,91,0,212,0,0,0,206,0,251,0,0,0,190,0,129,0,196,0,0,0,106,0,0,0,29,0,0,0,0,0,65,0,87,0,185,0,0,0,145,0,152,0,0,0,230,0,70,0,141,0,98,0,154,0,135,0,212,0,37,0,164,0,62,0,145,0,237,0,212,0,0,0,0,0,92,0,0,0,82,0,85,0,69,0,153,0,114,0,107,0,0,0,232,0,111,0,248,0,233,0,136,0,19,0,222,0,44,0,141,0,187,0,0,0,0,0,132,0,11,0,88,0,0,0,16,0,136,0,146,0,0,0,255,0,19,0,134,0,195,0,30,0,193,0,77,0,247,0,140,0,78,0,0,0,170,0,122,0,201,0,170,0,30,0,253,0,91,0,97,0,196,0,61,0,143,0,176,0,58,0,187,0,184,0,180,0,183,0,16,0,70,0,0,0,204,0,100,0,26,0,40,0,38,0,0,0,159,0,236,0,66,0,38,0,100,0,39,0,188,0,202,0,212,0,129,0,59,0,193,0,79,0,130,0,31,0,4,0,85,0,16,0,244,0,244,0,204,0,66,0,198,0,101,0,0,0,0,0,0,0,0,0,38,0,229,0,89,0,0,0,238,0,228,0,0,0,16,0,147,0,134,0,166,0,0,0,160,0,0,0,8,0,153,0,248,0,87,0,235,0,0,0,149,0,1,0,224,0,101,0,224,0,200,0,0,0,0,0,247,0,59,0,162,0,0,0,255,0,249,0,50,0,20,0,171,0,0,0,247,0,217,0,0,0,222,0,212,0,0,0,206,0,138,0,205,0,60,0,0,0,103,0,6,0,66,0,156,0,45,0,54,0,68,0,144,0,0,0,58,0,67,0,240,0,9,0,76,0,57,0,189,0,82,0,141,0,0,0,39,0,106,0,192,0,193,0,248,0,0,0,0,0,111,0,72,0,0,0,0,0,122,0,50,0,0,0,0,0,238,0,21,0,0,0,0,0,174,0,147,0,131,0,0,0,100,0,244,0,94,0,27,0,142,0,122,0,253,0,223,0,242,0,96,0,212,0,0,0,195,0,222,0,2,0,1,0,138,0,0,0,125,0,142,0,0,0,242,0,187,0,68,0,49,0,58,0,0,0,85,0,0,0,105,0,63,0,254,0,235,0,99,0,36,0,156,0,181,0,117,0,49,0,79,0,176,0,94,0,0,0,194,0,0,0,234,0,26,0,215,0,0,0,28,0,0,0,232,0,211,0,0,0,167,0,0,0,41,0,206,0,245,0,129,0,121,0,168,0,251,0,115,0,0,0,210,0,115,0,12,0,255,0,148,0,155,0,142,0,35,0,133,0,166,0,0,0,221,0,0,0,12,0,77,0,236,0,0,0,94,0,112,0,161,0,217,0,79,0,186,0,23,0,0,0,200,0,213,0,154,0,18,0,143,0,254,0,77,0);
signal scenario_full  : scenario_type := (159,31,98,31,144,31,248,31,203,31,203,30,255,31,208,31,248,31,201,31,7,31,7,30,7,29,204,31,136,31,136,30,235,31,229,31,9,31,39,31,182,31,182,30,26,31,26,30,26,29,26,28,65,31,65,30,97,31,4,31,51,31,81,31,86,31,86,30,200,31,250,31,252,31,33,31,161,31,25,31,149,31,199,31,43,31,43,30,43,29,171,31,78,31,78,30,78,29,78,28,109,31,120,31,120,30,151,31,34,31,34,30,230,31,230,30,230,29,230,28,102,31,16,31,16,30,100,31,165,31,40,31,40,30,40,29,40,28,112,31,103,31,165,31,69,31,142,31,192,31,203,31,187,31,168,31,191,31,1,31,50,31,129,31,129,30,12,31,168,31,168,30,55,31,55,30,135,31,3,31,132,31,54,31,81,31,81,30,203,31,247,31,80,31,202,31,86,31,83,31,225,31,225,30,78,31,215,31,182,31,51,31,51,30,54,31,96,31,96,30,149,31,149,30,99,31,39,31,39,30,134,31,91,31,91,30,166,31,244,31,234,31,234,30,234,29,239,31,252,31,19,31,19,30,177,31,198,31,107,31,61,31,61,30,211,31,180,31,31,31,72,31,97,31,97,30,83,31,125,31,124,31,199,31,18,31,76,31,76,30,76,29,80,31,15,31,151,31,120,31,120,30,146,31,146,30,105,31,48,31,48,30,134,31,231,31,231,30,70,31,70,30,129,31,77,31,142,31,29,31,38,31,18,31,40,31,7,31,7,30,7,29,214,31,94,31,94,30,90,31,90,30,90,29,90,28,161,31,111,31,111,30,194,31,169,31,37,31,34,31,54,31,158,31,195,31,10,31,10,30,191,31,191,30,52,31,153,31,33,31,33,30,21,31,161,31,19,31,168,31,43,31,180,31,221,31,12,31,175,31,175,30,147,31,95,31,95,30,92,31,115,31,115,30,136,31,176,31,122,31,160,31,51,31,38,31,140,31,159,31,255,31,40,31,170,31,70,31,82,31,82,30,69,31,52,31,99,31,197,31,18,31,33,31,33,30,2,31,196,31,196,30,196,29,117,31,117,30,103,31,98,31,29,31,123,31,246,31,168,31,140,31,44,31,218,31,144,31,144,30,174,31,208,31,22,31,222,31,14,31,205,31,175,31,20,31,72,31,88,31,211,31,101,31,243,31,180,31,249,31,23,31,35,31,42,31,42,31,6,31,178,31,155,31,109,31,144,31,222,31,129,31,7,31,95,31,41,31,80,31,58,31,16,31,16,30,71,31,251,31,251,30,101,31,132,31,149,31,127,31,20,31,247,31,6,31,85,31,159,31,128,31,186,31,55,31,62,31,179,31,86,31,188,31,42,31,132,31,56,31,208,31,146,31,158,31,172,31,245,31,115,31,26,31,38,31,248,31,229,31,15,31,101,31,12,31,30,31,133,31,249,31,249,30,24,31,22,31,14,31,180,31,41,31,177,31,240,31,138,31,197,31,249,31,215,31,151,31,158,31,106,31,118,31,155,31,129,31,129,30,87,31,133,31,133,30,46,31,246,31,35,31,171,31,171,30,246,31,170,31,209,31,115,31,114,31,91,31,153,31,90,31,102,31,220,31,220,30,101,31,101,30,23,31,91,31,212,31,212,30,206,31,251,31,251,30,190,31,129,31,196,31,196,30,106,31,106,30,29,31,29,30,29,29,65,31,87,31,185,31,185,30,145,31,152,31,152,30,230,31,70,31,141,31,98,31,154,31,135,31,212,31,37,31,164,31,62,31,145,31,237,31,212,31,212,30,212,29,92,31,92,30,82,31,85,31,69,31,153,31,114,31,107,31,107,30,232,31,111,31,248,31,233,31,136,31,19,31,222,31,44,31,141,31,187,31,187,30,187,29,132,31,11,31,88,31,88,30,16,31,136,31,146,31,146,30,255,31,19,31,134,31,195,31,30,31,193,31,77,31,247,31,140,31,78,31,78,30,170,31,122,31,201,31,170,31,30,31,253,31,91,31,97,31,196,31,61,31,143,31,176,31,58,31,187,31,184,31,180,31,183,31,16,31,70,31,70,30,204,31,100,31,26,31,40,31,38,31,38,30,159,31,236,31,66,31,38,31,100,31,39,31,188,31,202,31,212,31,129,31,59,31,193,31,79,31,130,31,31,31,4,31,85,31,16,31,244,31,244,31,204,31,66,31,198,31,101,31,101,30,101,29,101,28,101,27,38,31,229,31,89,31,89,30,238,31,228,31,228,30,16,31,147,31,134,31,166,31,166,30,160,31,160,30,8,31,153,31,248,31,87,31,235,31,235,30,149,31,1,31,224,31,101,31,224,31,200,31,200,30,200,29,247,31,59,31,162,31,162,30,255,31,249,31,50,31,20,31,171,31,171,30,247,31,217,31,217,30,222,31,212,31,212,30,206,31,138,31,205,31,60,31,60,30,103,31,6,31,66,31,156,31,45,31,54,31,68,31,144,31,144,30,58,31,67,31,240,31,9,31,76,31,57,31,189,31,82,31,141,31,141,30,39,31,106,31,192,31,193,31,248,31,248,30,248,29,111,31,72,31,72,30,72,29,122,31,50,31,50,30,50,29,238,31,21,31,21,30,21,29,174,31,147,31,131,31,131,30,100,31,244,31,94,31,27,31,142,31,122,31,253,31,223,31,242,31,96,31,212,31,212,30,195,31,222,31,2,31,1,31,138,31,138,30,125,31,142,31,142,30,242,31,187,31,68,31,49,31,58,31,58,30,85,31,85,30,105,31,63,31,254,31,235,31,99,31,36,31,156,31,181,31,117,31,49,31,79,31,176,31,94,31,94,30,194,31,194,30,234,31,26,31,215,31,215,30,28,31,28,30,232,31,211,31,211,30,167,31,167,30,41,31,206,31,245,31,129,31,121,31,168,31,251,31,115,31,115,30,210,31,115,31,12,31,255,31,148,31,155,31,142,31,35,31,133,31,166,31,166,30,221,31,221,30,12,31,77,31,236,31,236,30,94,31,112,31,161,31,217,31,79,31,186,31,23,31,23,30,200,31,213,31,154,31,18,31,143,31,254,31,77,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
