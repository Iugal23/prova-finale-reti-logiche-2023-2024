-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_923 is
end project_tb_923;

architecture project_tb_arch_923 of project_tb_923 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 804;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,205,0,34,0,66,0,153,0,171,0,114,0,103,0,209,0,91,0,199,0,243,0,0,0,103,0,107,0,231,0,49,0,26,0,207,0,93,0,0,0,152,0,0,0,170,0,203,0,0,0,143,0,223,0,0,0,99,0,128,0,68,0,21,0,151,0,135,0,27,0,215,0,94,0,137,0,181,0,0,0,229,0,82,0,237,0,35,0,21,0,17,0,191,0,70,0,27,0,59,0,67,0,0,0,0,0,154,0,0,0,39,0,170,0,47,0,121,0,184,0,10,0,34,0,0,0,120,0,20,0,0,0,85,0,39,0,155,0,194,0,87,0,157,0,249,0,0,0,85,0,248,0,99,0,14,0,0,0,135,0,35,0,0,0,4,0,226,0,0,0,149,0,46,0,0,0,161,0,21,0,189,0,152,0,184,0,232,0,233,0,141,0,110,0,245,0,114,0,0,0,202,0,19,0,103,0,255,0,60,0,0,0,207,0,215,0,24,0,108,0,208,0,22,0,0,0,255,0,0,0,143,0,195,0,0,0,81,0,0,0,204,0,143,0,6,0,192,0,209,0,86,0,176,0,230,0,153,0,133,0,232,0,20,0,68,0,36,0,0,0,110,0,224,0,119,0,186,0,189,0,64,0,153,0,0,0,0,0,0,0,0,0,27,0,86,0,118,0,70,0,81,0,44,0,65,0,0,0,197,0,41,0,201,0,187,0,0,0,181,0,150,0,0,0,217,0,0,0,50,0,125,0,47,0,186,0,26,0,0,0,74,0,160,0,237,0,130,0,15,0,214,0,4,0,0,0,100,0,45,0,103,0,86,0,0,0,77,0,116,0,13,0,36,0,144,0,0,0,190,0,110,0,99,0,0,0,0,0,224,0,4,0,188,0,147,0,0,0,235,0,238,0,94,0,131,0,227,0,40,0,49,0,150,0,0,0,223,0,0,0,29,0,105,0,27,0,57,0,60,0,213,0,0,0,0,0,6,0,81,0,76,0,204,0,38,0,71,0,30,0,25,0,0,0,212,0,241,0,80,0,185,0,108,0,89,0,0,0,0,0,65,0,0,0,221,0,96,0,36,0,132,0,159,0,33,0,49,0,167,0,0,0,35,0,13,0,63,0,80,0,240,0,196,0,208,0,22,0,251,0,170,0,0,0,198,0,100,0,153,0,185,0,153,0,71,0,209,0,158,0,6,0,44,0,28,0,131,0,0,0,173,0,90,0,46,0,169,0,27,0,0,0,241,0,50,0,55,0,67,0,63,0,0,0,96,0,113,0,0,0,0,0,126,0,0,0,0,0,16,0,249,0,39,0,147,0,167,0,31,0,81,0,171,0,0,0,166,0,106,0,0,0,98,0,0,0,111,0,4,0,117,0,112,0,185,0,184,0,52,0,233,0,221,0,45,0,159,0,90,0,209,0,234,0,45,0,0,0,119,0,226,0,0,0,227,0,191,0,56,0,191,0,0,0,240,0,151,0,223,0,103,0,66,0,66,0,106,0,84,0,160,0,133,0,29,0,0,0,108,0,199,0,170,0,108,0,250,0,85,0,0,0,206,0,199,0,84,0,90,0,140,0,194,0,0,0,149,0,0,0,197,0,218,0,36,0,139,0,35,0,192,0,130,0,200,0,246,0,58,0,247,0,253,0,0,0,118,0,160,0,0,0,123,0,60,0,206,0,149,0,78,0,78,0,1,0,0,0,244,0,199,0,117,0,176,0,105,0,128,0,230,0,36,0,125,0,212,0,127,0,13,0,0,0,133,0,54,0,234,0,18,0,0,0,71,0,157,0,18,0,16,0,153,0,205,0,43,0,75,0,78,0,0,0,137,0,0,0,52,0,110,0,119,0,98,0,72,0,202,0,202,0,0,0,16,0,127,0,227,0,252,0,53,0,129,0,179,0,0,0,245,0,0,0,0,0,174,0,0,0,178,0,194,0,45,0,63,0,118,0,165,0,233,0,71,0,80,0,209,0,0,0,0,0,222,0,111,0,119,0,37,0,92,0,34,0,174,0,38,0,45,0,197,0,205,0,122,0,231,0,34,0,124,0,120,0,0,0,135,0,97,0,72,0,0,0,4,0,159,0,0,0,96,0,163,0,28,0,0,0,243,0,114,0,83,0,0,0,204,0,255,0,0,0,183,0,218,0,247,0,229,0,47,0,1,0,0,0,130,0,180,0,219,0,221,0,72,0,4,0,0,0,141,0,101,0,0,0,169,0,101,0,77,0,103,0,67,0,0,0,147,0,0,0,151,0,162,0,2,0,153,0,34,0,61,0,162,0,89,0,36,0,10,0,0,0,188,0,57,0,120,0,47,0,200,0,0,0,103,0,0,0,101,0,50,0,0,0,0,0,0,0,107,0,0,0,0,0,102,0,164,0,239,0,0,0,55,0,166,0,121,0,114,0,255,0,213,0,215,0,23,0,0,0,0,0,62,0,0,0,0,0,216,0,152,0,199,0,0,0,178,0,194,0,91,0,106,0,74,0,67,0,37,0,0,0,102,0,100,0,98,0,54,0,81,0,110,0,141,0,247,0,136,0,245,0,126,0,31,0,158,0,223,0,0,0,60,0,136,0,0,0,0,0,49,0,75,0,25,0,92,0,138,0,208,0,97,0,164,0,43,0,75,0,84,0,133,0,146,0,60,0,36,0,32,0,43,0,247,0,189,0,0,0,0,0,13,0,220,0,225,0,0,0,138,0,165,0,175,0,246,0,36,0,62,0,208,0,104,0,193,0,0,0,243,0,116,0,35,0,0,0,32,0,244,0,204,0,0,0,0,0,178,0,0,0,100,0,7,0,153,0,0,0,135,0,227,0,0,0,53,0,0,0,146,0,159,0,246,0,219,0,238,0,211,0,123,0,79,0,13,0,179,0,1,0,77,0,0,0,36,0,88,0,0,0,0,0,0,0,239,0,58,0,148,0,185,0,0,0,203,0,66,0,50,0,121,0,111,0,0,0,0,0,0,0,199,0,118,0,198,0,0,0,204,0,0,0,133,0,65,0,121,0,35,0,111,0,236,0,26,0,236,0,0,0,0,0,10,0,14,0,0,0,0,0,106,0,0,0,208,0,181,0,221,0,249,0,0,0,142,0,87,0,0,0,0,0,140,0,101,0,0,0,103,0,180,0,0,0,118,0,244,0,238,0,0,0,78,0,108,0,143,0,105,0,161,0,234,0,155,0,130,0,249,0,85,0,0,0,16,0,198,0,18,0,138,0,36,0,152,0,216,0,0,0,12,0,85,0,105,0,139,0,210,0,0,0,0,0,215,0,184,0,18,0,0,0,196,0,0,0,232,0,176,0,207,0,234,0,0,0,0,0,2,0,44,0,167,0,95,0,192,0,130,0,92,0,3,0,80,0,0,0,0,0,8,0,19,0,103,0,155,0,108,0,44,0,203,0,242,0,103,0,245,0,0,0,0,0,21,0,75,0,155,0,148,0,0,0,225,0,186,0,0,0,93,0,100,0,228,0,250,0,216,0,194,0,151,0,187,0,0,0,189,0,0,0,156,0,186,0,152,0,3,0,93,0,25,0,0,0,99,0,79,0,191,0,108,0,243,0,75,0,230,0,127,0,66,0,5,0,68,0,64,0);
signal scenario_full  : scenario_type := (0,0,205,31,34,31,66,31,153,31,171,31,114,31,103,31,209,31,91,31,199,31,243,31,243,30,103,31,107,31,231,31,49,31,26,31,207,31,93,31,93,30,152,31,152,30,170,31,203,31,203,30,143,31,223,31,223,30,99,31,128,31,68,31,21,31,151,31,135,31,27,31,215,31,94,31,137,31,181,31,181,30,229,31,82,31,237,31,35,31,21,31,17,31,191,31,70,31,27,31,59,31,67,31,67,30,67,29,154,31,154,30,39,31,170,31,47,31,121,31,184,31,10,31,34,31,34,30,120,31,20,31,20,30,85,31,39,31,155,31,194,31,87,31,157,31,249,31,249,30,85,31,248,31,99,31,14,31,14,30,135,31,35,31,35,30,4,31,226,31,226,30,149,31,46,31,46,30,161,31,21,31,189,31,152,31,184,31,232,31,233,31,141,31,110,31,245,31,114,31,114,30,202,31,19,31,103,31,255,31,60,31,60,30,207,31,215,31,24,31,108,31,208,31,22,31,22,30,255,31,255,30,143,31,195,31,195,30,81,31,81,30,204,31,143,31,6,31,192,31,209,31,86,31,176,31,230,31,153,31,133,31,232,31,20,31,68,31,36,31,36,30,110,31,224,31,119,31,186,31,189,31,64,31,153,31,153,30,153,29,153,28,153,27,27,31,86,31,118,31,70,31,81,31,44,31,65,31,65,30,197,31,41,31,201,31,187,31,187,30,181,31,150,31,150,30,217,31,217,30,50,31,125,31,47,31,186,31,26,31,26,30,74,31,160,31,237,31,130,31,15,31,214,31,4,31,4,30,100,31,45,31,103,31,86,31,86,30,77,31,116,31,13,31,36,31,144,31,144,30,190,31,110,31,99,31,99,30,99,29,224,31,4,31,188,31,147,31,147,30,235,31,238,31,94,31,131,31,227,31,40,31,49,31,150,31,150,30,223,31,223,30,29,31,105,31,27,31,57,31,60,31,213,31,213,30,213,29,6,31,81,31,76,31,204,31,38,31,71,31,30,31,25,31,25,30,212,31,241,31,80,31,185,31,108,31,89,31,89,30,89,29,65,31,65,30,221,31,96,31,36,31,132,31,159,31,33,31,49,31,167,31,167,30,35,31,13,31,63,31,80,31,240,31,196,31,208,31,22,31,251,31,170,31,170,30,198,31,100,31,153,31,185,31,153,31,71,31,209,31,158,31,6,31,44,31,28,31,131,31,131,30,173,31,90,31,46,31,169,31,27,31,27,30,241,31,50,31,55,31,67,31,63,31,63,30,96,31,113,31,113,30,113,29,126,31,126,30,126,29,16,31,249,31,39,31,147,31,167,31,31,31,81,31,171,31,171,30,166,31,106,31,106,30,98,31,98,30,111,31,4,31,117,31,112,31,185,31,184,31,52,31,233,31,221,31,45,31,159,31,90,31,209,31,234,31,45,31,45,30,119,31,226,31,226,30,227,31,191,31,56,31,191,31,191,30,240,31,151,31,223,31,103,31,66,31,66,31,106,31,84,31,160,31,133,31,29,31,29,30,108,31,199,31,170,31,108,31,250,31,85,31,85,30,206,31,199,31,84,31,90,31,140,31,194,31,194,30,149,31,149,30,197,31,218,31,36,31,139,31,35,31,192,31,130,31,200,31,246,31,58,31,247,31,253,31,253,30,118,31,160,31,160,30,123,31,60,31,206,31,149,31,78,31,78,31,1,31,1,30,244,31,199,31,117,31,176,31,105,31,128,31,230,31,36,31,125,31,212,31,127,31,13,31,13,30,133,31,54,31,234,31,18,31,18,30,71,31,157,31,18,31,16,31,153,31,205,31,43,31,75,31,78,31,78,30,137,31,137,30,52,31,110,31,119,31,98,31,72,31,202,31,202,31,202,30,16,31,127,31,227,31,252,31,53,31,129,31,179,31,179,30,245,31,245,30,245,29,174,31,174,30,178,31,194,31,45,31,63,31,118,31,165,31,233,31,71,31,80,31,209,31,209,30,209,29,222,31,111,31,119,31,37,31,92,31,34,31,174,31,38,31,45,31,197,31,205,31,122,31,231,31,34,31,124,31,120,31,120,30,135,31,97,31,72,31,72,30,4,31,159,31,159,30,96,31,163,31,28,31,28,30,243,31,114,31,83,31,83,30,204,31,255,31,255,30,183,31,218,31,247,31,229,31,47,31,1,31,1,30,130,31,180,31,219,31,221,31,72,31,4,31,4,30,141,31,101,31,101,30,169,31,101,31,77,31,103,31,67,31,67,30,147,31,147,30,151,31,162,31,2,31,153,31,34,31,61,31,162,31,89,31,36,31,10,31,10,30,188,31,57,31,120,31,47,31,200,31,200,30,103,31,103,30,101,31,50,31,50,30,50,29,50,28,107,31,107,30,107,29,102,31,164,31,239,31,239,30,55,31,166,31,121,31,114,31,255,31,213,31,215,31,23,31,23,30,23,29,62,31,62,30,62,29,216,31,152,31,199,31,199,30,178,31,194,31,91,31,106,31,74,31,67,31,37,31,37,30,102,31,100,31,98,31,54,31,81,31,110,31,141,31,247,31,136,31,245,31,126,31,31,31,158,31,223,31,223,30,60,31,136,31,136,30,136,29,49,31,75,31,25,31,92,31,138,31,208,31,97,31,164,31,43,31,75,31,84,31,133,31,146,31,60,31,36,31,32,31,43,31,247,31,189,31,189,30,189,29,13,31,220,31,225,31,225,30,138,31,165,31,175,31,246,31,36,31,62,31,208,31,104,31,193,31,193,30,243,31,116,31,35,31,35,30,32,31,244,31,204,31,204,30,204,29,178,31,178,30,100,31,7,31,153,31,153,30,135,31,227,31,227,30,53,31,53,30,146,31,159,31,246,31,219,31,238,31,211,31,123,31,79,31,13,31,179,31,1,31,77,31,77,30,36,31,88,31,88,30,88,29,88,28,239,31,58,31,148,31,185,31,185,30,203,31,66,31,50,31,121,31,111,31,111,30,111,29,111,28,199,31,118,31,198,31,198,30,204,31,204,30,133,31,65,31,121,31,35,31,111,31,236,31,26,31,236,31,236,30,236,29,10,31,14,31,14,30,14,29,106,31,106,30,208,31,181,31,221,31,249,31,249,30,142,31,87,31,87,30,87,29,140,31,101,31,101,30,103,31,180,31,180,30,118,31,244,31,238,31,238,30,78,31,108,31,143,31,105,31,161,31,234,31,155,31,130,31,249,31,85,31,85,30,16,31,198,31,18,31,138,31,36,31,152,31,216,31,216,30,12,31,85,31,105,31,139,31,210,31,210,30,210,29,215,31,184,31,18,31,18,30,196,31,196,30,232,31,176,31,207,31,234,31,234,30,234,29,2,31,44,31,167,31,95,31,192,31,130,31,92,31,3,31,80,31,80,30,80,29,8,31,19,31,103,31,155,31,108,31,44,31,203,31,242,31,103,31,245,31,245,30,245,29,21,31,75,31,155,31,148,31,148,30,225,31,186,31,186,30,93,31,100,31,228,31,250,31,216,31,194,31,151,31,187,31,187,30,189,31,189,30,156,31,186,31,152,31,3,31,93,31,25,31,25,30,99,31,79,31,191,31,108,31,243,31,75,31,230,31,127,31,66,31,5,31,68,31,64,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
