-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 432;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,79,0,240,0,114,0,0,0,45,0,216,0,157,0,142,0,58,0,0,0,214,0,226,0,122,0,104,0,94,0,31,0,31,0,30,0,0,0,96,0,175,0,177,0,105,0,0,0,46,0,26,0,185,0,0,0,209,0,26,0,2,0,229,0,47,0,0,0,36,0,239,0,209,0,162,0,79,0,23,0,79,0,205,0,0,0,74,0,0,0,176,0,79,0,242,0,239,0,173,0,155,0,0,0,61,0,173,0,133,0,24,0,165,0,217,0,0,0,173,0,42,0,160,0,36,0,0,0,232,0,29,0,244,0,115,0,174,0,238,0,198,0,22,0,247,0,28,0,0,0,88,0,43,0,254,0,32,0,232,0,156,0,181,0,0,0,85,0,149,0,86,0,17,0,219,0,97,0,252,0,103,0,0,0,183,0,227,0,42,0,117,0,0,0,76,0,39,0,99,0,20,0,0,0,0,0,26,0,160,0,0,0,0,0,0,0,0,0,0,0,134,0,239,0,213,0,90,0,136,0,0,0,41,0,135,0,247,0,0,0,32,0,133,0,252,0,0,0,217,0,190,0,42,0,0,0,0,0,236,0,91,0,175,0,175,0,81,0,95,0,108,0,85,0,51,0,69,0,85,0,0,0,15,0,67,0,164,0,252,0,164,0,112,0,61,0,57,0,8,0,118,0,114,0,250,0,194,0,207,0,208,0,0,0,62,0,10,0,129,0,237,0,0,0,44,0,164,0,97,0,35,0,226,0,8,0,104,0,205,0,150,0,139,0,128,0,192,0,0,0,42,0,0,0,183,0,51,0,0,0,30,0,218,0,144,0,127,0,184,0,230,0,190,0,111,0,0,0,238,0,20,0,10,0,176,0,239,0,154,0,180,0,195,0,169,0,65,0,234,0,0,0,231,0,0,0,121,0,197,0,253,0,18,0,117,0,154,0,133,0,0,0,181,0,201,0,0,0,178,0,137,0,0,0,26,0,49,0,66,0,229,0,17,0,0,0,78,0,0,0,151,0,0,0,179,0,0,0,11,0,56,0,126,0,137,0,84,0,0,0,231,0,123,0,0,0,138,0,140,0,177,0,89,0,19,0,151,0,134,0,0,0,121,0,2,0,181,0,98,0,0,0,130,0,110,0,16,0,0,0,244,0,0,0,113,0,0,0,227,0,170,0,150,0,0,0,239,0,246,0,0,0,160,0,110,0,63,0,46,0,36,0,176,0,133,0,58,0,0,0,163,0,180,0,122,0,157,0,156,0,127,0,241,0,168,0,150,0,157,0,114,0,75,0,167,0,219,0,117,0,191,0,181,0,232,0,191,0,180,0,233,0,127,0,0,0,165,0,0,0,43,0,138,0,246,0,214,0,0,0,62,0,228,0,160,0,92,0,144,0,9,0,0,0,52,0,111,0,236,0,0,0,249,0,60,0,92,0,128,0,157,0,0,0,112,0,193,0,0,0,246,0,59,0,25,0,160,0,0,0,128,0,240,0,0,0,0,0,0,0,0,0,223,0,52,0,47,0,70,0,0,0,0,0,62,0,106,0,140,0,149,0,145,0,0,0,252,0,52,0,0,0,0,0,228,0,162,0,150,0,0,0,253,0,248,0,0,0,0,0,0,0,37,0,241,0,42,0,63,0,226,0,129,0,54,0,232,0,113,0,0,0,190,0,224,0,29,0,0,0,5,0,0,0,226,0,211,0,70,0,174,0,71,0,235,0,178,0,0,0,171,0,225,0,0,0,101,0,72,0,165,0,48,0,91,0,31,0,255,0,197,0,0,0,142,0,43,0,0,0,166,0,70,0,147,0,63,0,165,0,228,0,187,0,159,0,29,0,181,0,0,0,224,0,154,0,159,0,87,0,168,0,187,0,0,0,0,0,100,0,0,0,191,0,253,0,70,0,0,0,61,0,0,0,26,0,0,0,0,0,29,0);
signal scenario_full  : scenario_type := (0,0,79,31,240,31,114,31,114,30,45,31,216,31,157,31,142,31,58,31,58,30,214,31,226,31,122,31,104,31,94,31,31,31,31,31,30,31,30,30,96,31,175,31,177,31,105,31,105,30,46,31,26,31,185,31,185,30,209,31,26,31,2,31,229,31,47,31,47,30,36,31,239,31,209,31,162,31,79,31,23,31,79,31,205,31,205,30,74,31,74,30,176,31,79,31,242,31,239,31,173,31,155,31,155,30,61,31,173,31,133,31,24,31,165,31,217,31,217,30,173,31,42,31,160,31,36,31,36,30,232,31,29,31,244,31,115,31,174,31,238,31,198,31,22,31,247,31,28,31,28,30,88,31,43,31,254,31,32,31,232,31,156,31,181,31,181,30,85,31,149,31,86,31,17,31,219,31,97,31,252,31,103,31,103,30,183,31,227,31,42,31,117,31,117,30,76,31,39,31,99,31,20,31,20,30,20,29,26,31,160,31,160,30,160,29,160,28,160,27,160,26,134,31,239,31,213,31,90,31,136,31,136,30,41,31,135,31,247,31,247,30,32,31,133,31,252,31,252,30,217,31,190,31,42,31,42,30,42,29,236,31,91,31,175,31,175,31,81,31,95,31,108,31,85,31,51,31,69,31,85,31,85,30,15,31,67,31,164,31,252,31,164,31,112,31,61,31,57,31,8,31,118,31,114,31,250,31,194,31,207,31,208,31,208,30,62,31,10,31,129,31,237,31,237,30,44,31,164,31,97,31,35,31,226,31,8,31,104,31,205,31,150,31,139,31,128,31,192,31,192,30,42,31,42,30,183,31,51,31,51,30,30,31,218,31,144,31,127,31,184,31,230,31,190,31,111,31,111,30,238,31,20,31,10,31,176,31,239,31,154,31,180,31,195,31,169,31,65,31,234,31,234,30,231,31,231,30,121,31,197,31,253,31,18,31,117,31,154,31,133,31,133,30,181,31,201,31,201,30,178,31,137,31,137,30,26,31,49,31,66,31,229,31,17,31,17,30,78,31,78,30,151,31,151,30,179,31,179,30,11,31,56,31,126,31,137,31,84,31,84,30,231,31,123,31,123,30,138,31,140,31,177,31,89,31,19,31,151,31,134,31,134,30,121,31,2,31,181,31,98,31,98,30,130,31,110,31,16,31,16,30,244,31,244,30,113,31,113,30,227,31,170,31,150,31,150,30,239,31,246,31,246,30,160,31,110,31,63,31,46,31,36,31,176,31,133,31,58,31,58,30,163,31,180,31,122,31,157,31,156,31,127,31,241,31,168,31,150,31,157,31,114,31,75,31,167,31,219,31,117,31,191,31,181,31,232,31,191,31,180,31,233,31,127,31,127,30,165,31,165,30,43,31,138,31,246,31,214,31,214,30,62,31,228,31,160,31,92,31,144,31,9,31,9,30,52,31,111,31,236,31,236,30,249,31,60,31,92,31,128,31,157,31,157,30,112,31,193,31,193,30,246,31,59,31,25,31,160,31,160,30,128,31,240,31,240,30,240,29,240,28,240,27,223,31,52,31,47,31,70,31,70,30,70,29,62,31,106,31,140,31,149,31,145,31,145,30,252,31,52,31,52,30,52,29,228,31,162,31,150,31,150,30,253,31,248,31,248,30,248,29,248,28,37,31,241,31,42,31,63,31,226,31,129,31,54,31,232,31,113,31,113,30,190,31,224,31,29,31,29,30,5,31,5,30,226,31,211,31,70,31,174,31,71,31,235,31,178,31,178,30,171,31,225,31,225,30,101,31,72,31,165,31,48,31,91,31,31,31,255,31,197,31,197,30,142,31,43,31,43,30,166,31,70,31,147,31,63,31,165,31,228,31,187,31,159,31,29,31,181,31,181,30,224,31,154,31,159,31,87,31,168,31,187,31,187,30,187,29,100,31,100,30,191,31,253,31,70,31,70,30,61,31,61,30,26,31,26,30,26,29,29,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
