-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_788 is
end project_tb_788;

architecture project_tb_arch_788 of project_tb_788 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 841;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,7,0,146,0,240,0,205,0,79,0,227,0,213,0,209,0,253,0,0,0,10,0,0,0,0,0,0,0,2,0,0,0,212,0,184,0,237,0,77,0,202,0,88,0,12,0,52,0,67,0,141,0,0,0,224,0,241,0,109,0,95,0,224,0,158,0,5,0,0,0,214,0,38,0,191,0,0,0,177,0,74,0,192,0,111,0,206,0,230,0,21,0,128,0,63,0,173,0,197,0,15,0,0,0,191,0,219,0,0,0,83,0,117,0,214,0,11,0,177,0,0,0,233,0,29,0,73,0,0,0,38,0,88,0,96,0,131,0,0,0,0,0,182,0,84,0,0,0,0,0,108,0,225,0,13,0,120,0,122,0,0,0,124,0,60,0,34,0,0,0,216,0,4,0,132,0,0,0,193,0,0,0,29,0,0,0,95,0,65,0,41,0,113,0,108,0,75,0,195,0,0,0,173,0,61,0,213,0,196,0,22,0,184,0,204,0,207,0,55,0,0,0,73,0,0,0,0,0,33,0,190,0,0,0,175,0,159,0,0,0,0,0,1,0,0,0,0,0,0,0,101,0,105,0,107,0,4,0,121,0,75,0,208,0,0,0,8,0,92,0,0,0,7,0,196,0,0,0,55,0,0,0,58,0,73,0,206,0,123,0,7,0,247,0,208,0,57,0,251,0,0,0,117,0,0,0,131,0,0,0,171,0,192,0,0,0,166,0,196,0,169,0,209,0,244,0,195,0,17,0,0,0,68,0,0,0,2,0,47,0,218,0,188,0,0,0,64,0,206,0,35,0,103,0,0,0,72,0,186,0,162,0,204,0,147,0,131,0,12,0,0,0,3,0,0,0,226,0,131,0,141,0,203,0,134,0,226,0,31,0,0,0,196,0,254,0,190,0,121,0,130,0,144,0,0,0,95,0,27,0,172,0,0,0,247,0,0,0,224,0,237,0,0,0,36,0,54,0,202,0,77,0,169,0,97,0,0,0,0,0,227,0,208,0,188,0,211,0,178,0,152,0,243,0,0,0,34,0,231,0,22,0,0,0,105,0,50,0,0,0,72,0,254,0,96,0,132,0,225,0,122,0,222,0,67,0,0,0,0,0,0,0,104,0,127,0,97,0,121,0,134,0,0,0,0,0,202,0,189,0,159,0,209,0,212,0,145,0,25,0,0,0,0,0,55,0,93,0,0,0,36,0,247,0,100,0,0,0,103,0,233,0,101,0,235,0,0,0,60,0,0,0,68,0,94,0,0,0,164,0,109,0,63,0,209,0,87,0,59,0,226,0,87,0,0,0,240,0,0,0,140,0,152,0,111,0,6,0,169,0,0,0,169,0,209,0,91,0,249,0,0,0,132,0,169,0,160,0,81,0,0,0,88,0,85,0,114,0,88,0,0,0,230,0,193,0,55,0,0,0,186,0,114,0,246,0,128,0,165,0,220,0,47,0,227,0,39,0,149,0,0,0,0,0,83,0,0,0,41,0,214,0,215,0,0,0,208,0,170,0,171,0,23,0,94,0,0,0,203,0,173,0,181,0,239,0,0,0,231,0,212,0,103,0,72,0,122,0,2,0,0,0,0,0,67,0,141,0,0,0,74,0,241,0,63,0,70,0,9,0,8,0,0,0,251,0,63,0,0,0,235,0,0,0,2,0,0,0,6,0,78,0,102,0,75,0,0,0,0,0,230,0,24,0,251,0,177,0,41,0,163,0,44,0,56,0,211,0,0,0,204,0,248,0,159,0,0,0,0,0,121,0,157,0,141,0,193,0,147,0,221,0,0,0,149,0,183,0,143,0,233,0,19,0,18,0,16,0,29,0,64,0,51,0,240,0,185,0,85,0,50,0,0,0,0,0,236,0,0,0,85,0,113,0,199,0,0,0,38,0,251,0,0,0,175,0,0,0,115,0,45,0,41,0,176,0,0,0,43,0,120,0,150,0,0,0,192,0,46,0,152,0,103,0,30,0,7,0,187,0,11,0,144,0,0,0,0,0,157,0,148,0,21,0,139,0,1,0,0,0,0,0,175,0,0,0,89,0,163,0,173,0,0,0,224,0,243,0,36,0,0,0,153,0,51,0,244,0,86,0,37,0,141,0,18,0,99,0,87,0,119,0,64,0,102,0,22,0,182,0,61,0,245,0,0,0,129,0,0,0,186,0,20,0,5,0,58,0,104,0,43,0,251,0,123,0,127,0,82,0,104,0,22,0,27,0,160,0,223,0,224,0,251,0,87,0,59,0,205,0,224,0,7,0,113,0,207,0,193,0,46,0,0,0,119,0,170,0,206,0,119,0,59,0,25,0,0,0,250,0,235,0,78,0,0,0,2,0,134,0,119,0,11,0,49,0,142,0,0,0,8,0,105,0,3,0,0,0,24,0,200,0,0,0,24,0,2,0,117,0,47,0,0,0,211,0,0,0,0,0,62,0,107,0,241,0,107,0,201,0,138,0,152,0,248,0,22,0,132,0,232,0,0,0,183,0,229,0,0,0,190,0,0,0,186,0,58,0,172,0,0,0,0,0,30,0,135,0,37,0,170,0,28,0,0,0,64,0,238,0,73,0,67,0,46,0,37,0,105,0,0,0,73,0,118,0,238,0,212,0,88,0,184,0,114,0,249,0,121,0,176,0,213,0,2,0,0,0,155,0,244,0,198,0,0,0,94,0,104,0,226,0,26,0,74,0,66,0,120,0,0,0,110,0,87,0,0,0,217,0,196,0,27,0,170,0,210,0,0,0,86,0,0,0,46,0,0,0,60,0,93,0,66,0,225,0,66,0,0,0,130,0,161,0,27,0,0,0,0,0,94,0,0,0,130,0,147,0,14,0,18,0,205,0,117,0,0,0,113,0,206,0,13,0,132,0,29,0,82,0,0,0,56,0,133,0,147,0,0,0,231,0,112,0,194,0,7,0,169,0,159,0,236,0,29,0,0,0,222,0,217,0,152,0,105,0,173,0,188,0,0,0,43,0,0,0,249,0,102,0,45,0,240,0,213,0,205,0,16,0,0,0,178,0,116,0,0,0,241,0,0,0,102,0,0,0,159,0,188,0,100,0,158,0,9,0,147,0,128,0,68,0,33,0,133,0,192,0,177,0,0,0,62,0,16,0,0,0,119,0,46,0,98,0,0,0,244,0,48,0,169,0,28,0,0,0,208,0,240,0,0,0,190,0,0,0,194,0,0,0,81,0,202,0,0,0,250,0,0,0,226,0,20,0,100,0,207,0,205,0,153,0,0,0,0,0,0,0,43,0,0,0,235,0,0,0,0,0,64,0,175,0,245,0,134,0,53,0,114,0,141,0,100,0,0,0,154,0,237,0,123,0,149,0,42,0,204,0,54,0,0,0,107,0,68,0,180,0,94,0,227,0,45,0,145,0,180,0,190,0,31,0,198,0,0,0,75,0,0,0,0,0,127,0,77,0,204,0,90,0,61,0,179,0,122,0,238,0,252,0,0,0,105,0,57,0,153,0,59,0,214,0,17,0,50,0,0,0,48,0,154,0,202,0,46,0,177,0,199,0,168,0,252,0,38,0,91,0,218,0,188,0,0,0,131,0,109,0,140,0,216,0,147,0,226,0,214,0,148,0,194,0,255,0,0,0,248,0,161,0,88,0,145,0,203,0,131,0,0,0,0,0,0,0,176,0,32,0,128,0,0,0,0,0,172,0,0,0,0,0,1,0,126,0,222,0,0,0,0,0,235,0,139,0,0,0,47,0,75,0,0,0,98,0,83,0,0,0,255,0,208,0,0,0,154,0,39,0,0,0);
signal scenario_full  : scenario_type := (0,0,7,31,146,31,240,31,205,31,79,31,227,31,213,31,209,31,253,31,253,30,10,31,10,30,10,29,10,28,2,31,2,30,212,31,184,31,237,31,77,31,202,31,88,31,12,31,52,31,67,31,141,31,141,30,224,31,241,31,109,31,95,31,224,31,158,31,5,31,5,30,214,31,38,31,191,31,191,30,177,31,74,31,192,31,111,31,206,31,230,31,21,31,128,31,63,31,173,31,197,31,15,31,15,30,191,31,219,31,219,30,83,31,117,31,214,31,11,31,177,31,177,30,233,31,29,31,73,31,73,30,38,31,88,31,96,31,131,31,131,30,131,29,182,31,84,31,84,30,84,29,108,31,225,31,13,31,120,31,122,31,122,30,124,31,60,31,34,31,34,30,216,31,4,31,132,31,132,30,193,31,193,30,29,31,29,30,95,31,65,31,41,31,113,31,108,31,75,31,195,31,195,30,173,31,61,31,213,31,196,31,22,31,184,31,204,31,207,31,55,31,55,30,73,31,73,30,73,29,33,31,190,31,190,30,175,31,159,31,159,30,159,29,1,31,1,30,1,29,1,28,101,31,105,31,107,31,4,31,121,31,75,31,208,31,208,30,8,31,92,31,92,30,7,31,196,31,196,30,55,31,55,30,58,31,73,31,206,31,123,31,7,31,247,31,208,31,57,31,251,31,251,30,117,31,117,30,131,31,131,30,171,31,192,31,192,30,166,31,196,31,169,31,209,31,244,31,195,31,17,31,17,30,68,31,68,30,2,31,47,31,218,31,188,31,188,30,64,31,206,31,35,31,103,31,103,30,72,31,186,31,162,31,204,31,147,31,131,31,12,31,12,30,3,31,3,30,226,31,131,31,141,31,203,31,134,31,226,31,31,31,31,30,196,31,254,31,190,31,121,31,130,31,144,31,144,30,95,31,27,31,172,31,172,30,247,31,247,30,224,31,237,31,237,30,36,31,54,31,202,31,77,31,169,31,97,31,97,30,97,29,227,31,208,31,188,31,211,31,178,31,152,31,243,31,243,30,34,31,231,31,22,31,22,30,105,31,50,31,50,30,72,31,254,31,96,31,132,31,225,31,122,31,222,31,67,31,67,30,67,29,67,28,104,31,127,31,97,31,121,31,134,31,134,30,134,29,202,31,189,31,159,31,209,31,212,31,145,31,25,31,25,30,25,29,55,31,93,31,93,30,36,31,247,31,100,31,100,30,103,31,233,31,101,31,235,31,235,30,60,31,60,30,68,31,94,31,94,30,164,31,109,31,63,31,209,31,87,31,59,31,226,31,87,31,87,30,240,31,240,30,140,31,152,31,111,31,6,31,169,31,169,30,169,31,209,31,91,31,249,31,249,30,132,31,169,31,160,31,81,31,81,30,88,31,85,31,114,31,88,31,88,30,230,31,193,31,55,31,55,30,186,31,114,31,246,31,128,31,165,31,220,31,47,31,227,31,39,31,149,31,149,30,149,29,83,31,83,30,41,31,214,31,215,31,215,30,208,31,170,31,171,31,23,31,94,31,94,30,203,31,173,31,181,31,239,31,239,30,231,31,212,31,103,31,72,31,122,31,2,31,2,30,2,29,67,31,141,31,141,30,74,31,241,31,63,31,70,31,9,31,8,31,8,30,251,31,63,31,63,30,235,31,235,30,2,31,2,30,6,31,78,31,102,31,75,31,75,30,75,29,230,31,24,31,251,31,177,31,41,31,163,31,44,31,56,31,211,31,211,30,204,31,248,31,159,31,159,30,159,29,121,31,157,31,141,31,193,31,147,31,221,31,221,30,149,31,183,31,143,31,233,31,19,31,18,31,16,31,29,31,64,31,51,31,240,31,185,31,85,31,50,31,50,30,50,29,236,31,236,30,85,31,113,31,199,31,199,30,38,31,251,31,251,30,175,31,175,30,115,31,45,31,41,31,176,31,176,30,43,31,120,31,150,31,150,30,192,31,46,31,152,31,103,31,30,31,7,31,187,31,11,31,144,31,144,30,144,29,157,31,148,31,21,31,139,31,1,31,1,30,1,29,175,31,175,30,89,31,163,31,173,31,173,30,224,31,243,31,36,31,36,30,153,31,51,31,244,31,86,31,37,31,141,31,18,31,99,31,87,31,119,31,64,31,102,31,22,31,182,31,61,31,245,31,245,30,129,31,129,30,186,31,20,31,5,31,58,31,104,31,43,31,251,31,123,31,127,31,82,31,104,31,22,31,27,31,160,31,223,31,224,31,251,31,87,31,59,31,205,31,224,31,7,31,113,31,207,31,193,31,46,31,46,30,119,31,170,31,206,31,119,31,59,31,25,31,25,30,250,31,235,31,78,31,78,30,2,31,134,31,119,31,11,31,49,31,142,31,142,30,8,31,105,31,3,31,3,30,24,31,200,31,200,30,24,31,2,31,117,31,47,31,47,30,211,31,211,30,211,29,62,31,107,31,241,31,107,31,201,31,138,31,152,31,248,31,22,31,132,31,232,31,232,30,183,31,229,31,229,30,190,31,190,30,186,31,58,31,172,31,172,30,172,29,30,31,135,31,37,31,170,31,28,31,28,30,64,31,238,31,73,31,67,31,46,31,37,31,105,31,105,30,73,31,118,31,238,31,212,31,88,31,184,31,114,31,249,31,121,31,176,31,213,31,2,31,2,30,155,31,244,31,198,31,198,30,94,31,104,31,226,31,26,31,74,31,66,31,120,31,120,30,110,31,87,31,87,30,217,31,196,31,27,31,170,31,210,31,210,30,86,31,86,30,46,31,46,30,60,31,93,31,66,31,225,31,66,31,66,30,130,31,161,31,27,31,27,30,27,29,94,31,94,30,130,31,147,31,14,31,18,31,205,31,117,31,117,30,113,31,206,31,13,31,132,31,29,31,82,31,82,30,56,31,133,31,147,31,147,30,231,31,112,31,194,31,7,31,169,31,159,31,236,31,29,31,29,30,222,31,217,31,152,31,105,31,173,31,188,31,188,30,43,31,43,30,249,31,102,31,45,31,240,31,213,31,205,31,16,31,16,30,178,31,116,31,116,30,241,31,241,30,102,31,102,30,159,31,188,31,100,31,158,31,9,31,147,31,128,31,68,31,33,31,133,31,192,31,177,31,177,30,62,31,16,31,16,30,119,31,46,31,98,31,98,30,244,31,48,31,169,31,28,31,28,30,208,31,240,31,240,30,190,31,190,30,194,31,194,30,81,31,202,31,202,30,250,31,250,30,226,31,20,31,100,31,207,31,205,31,153,31,153,30,153,29,153,28,43,31,43,30,235,31,235,30,235,29,64,31,175,31,245,31,134,31,53,31,114,31,141,31,100,31,100,30,154,31,237,31,123,31,149,31,42,31,204,31,54,31,54,30,107,31,68,31,180,31,94,31,227,31,45,31,145,31,180,31,190,31,31,31,198,31,198,30,75,31,75,30,75,29,127,31,77,31,204,31,90,31,61,31,179,31,122,31,238,31,252,31,252,30,105,31,57,31,153,31,59,31,214,31,17,31,50,31,50,30,48,31,154,31,202,31,46,31,177,31,199,31,168,31,252,31,38,31,91,31,218,31,188,31,188,30,131,31,109,31,140,31,216,31,147,31,226,31,214,31,148,31,194,31,255,31,255,30,248,31,161,31,88,31,145,31,203,31,131,31,131,30,131,29,131,28,176,31,32,31,128,31,128,30,128,29,172,31,172,30,172,29,1,31,126,31,222,31,222,30,222,29,235,31,139,31,139,30,47,31,75,31,75,30,98,31,83,31,83,30,255,31,208,31,208,30,154,31,39,31,39,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
