-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 190;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (248,0,113,0,141,0,0,0,174,0,88,0,0,0,108,0,208,0,46,0,44,0,213,0,210,0,194,0,69,0,24,0,235,0,0,0,28,0,0,0,92,0,57,0,59,0,49,0,49,0,215,0,240,0,44,0,102,0,106,0,0,0,246,0,159,0,49,0,0,0,167,0,160,0,0,0,46,0,3,0,192,0,0,0,179,0,196,0,233,0,85,0,244,0,0,0,55,0,118,0,74,0,164,0,199,0,80,0,29,0,12,0,155,0,182,0,13,0,114,0,183,0,30,0,190,0,0,0,17,0,47,0,113,0,70,0,78,0,65,0,231,0,155,0,17,0,57,0,94,0,185,0,0,0,0,0,196,0,192,0,41,0,46,0,86,0,80,0,211,0,19,0,202,0,158,0,102,0,3,0,43,0,242,0,151,0,0,0,63,0,138,0,248,0,135,0,0,0,0,0,221,0,0,0,0,0,70,0,139,0,202,0,245,0,0,0,134,0,219,0,123,0,125,0,250,0,13,0,121,0,179,0,214,0,0,0,12,0,64,0,0,0,130,0,144,0,81,0,250,0,218,0,110,0,80,0,175,0,188,0,48,0,4,0,152,0,225,0,59,0,223,0,234,0,159,0,0,0,32,0,36,0,173,0,111,0,156,0,131,0,230,0,102,0,0,0,43,0,99,0,0,0,15,0,58,0,0,0,150,0,71,0,21,0,0,0,137,0,117,0,148,0,0,0,89,0,40,0,0,0,172,0,0,0,33,0,199,0,164,0,179,0,41,0,0,0,126,0,0,0,0,0,68,0,0,0,181,0,87,0,33,0,199,0,88,0,246,0,155,0,0,0,128,0,0,0,104,0,0,0);
signal scenario_full  : scenario_type := (248,31,113,31,141,31,141,30,174,31,88,31,88,30,108,31,208,31,46,31,44,31,213,31,210,31,194,31,69,31,24,31,235,31,235,30,28,31,28,30,92,31,57,31,59,31,49,31,49,31,215,31,240,31,44,31,102,31,106,31,106,30,246,31,159,31,49,31,49,30,167,31,160,31,160,30,46,31,3,31,192,31,192,30,179,31,196,31,233,31,85,31,244,31,244,30,55,31,118,31,74,31,164,31,199,31,80,31,29,31,12,31,155,31,182,31,13,31,114,31,183,31,30,31,190,31,190,30,17,31,47,31,113,31,70,31,78,31,65,31,231,31,155,31,17,31,57,31,94,31,185,31,185,30,185,29,196,31,192,31,41,31,46,31,86,31,80,31,211,31,19,31,202,31,158,31,102,31,3,31,43,31,242,31,151,31,151,30,63,31,138,31,248,31,135,31,135,30,135,29,221,31,221,30,221,29,70,31,139,31,202,31,245,31,245,30,134,31,219,31,123,31,125,31,250,31,13,31,121,31,179,31,214,31,214,30,12,31,64,31,64,30,130,31,144,31,81,31,250,31,218,31,110,31,80,31,175,31,188,31,48,31,4,31,152,31,225,31,59,31,223,31,234,31,159,31,159,30,32,31,36,31,173,31,111,31,156,31,131,31,230,31,102,31,102,30,43,31,99,31,99,30,15,31,58,31,58,30,150,31,71,31,21,31,21,30,137,31,117,31,148,31,148,30,89,31,40,31,40,30,172,31,172,30,33,31,199,31,164,31,179,31,41,31,41,30,126,31,126,30,126,29,68,31,68,30,181,31,87,31,33,31,199,31,88,31,246,31,155,31,155,30,128,31,128,30,104,31,104,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
