-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_811 is
end project_tb_811;

architecture project_tb_arch_811 of project_tb_811 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 203;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (238,0,0,0,166,0,153,0,225,0,63,0,52,0,111,0,0,0,0,0,226,0,141,0,68,0,164,0,158,0,0,0,48,0,180,0,181,0,120,0,33,0,232,0,169,0,0,0,85,0,189,0,77,0,3,0,50,0,145,0,53,0,102,0,185,0,120,0,41,0,226,0,232,0,0,0,177,0,85,0,231,0,0,0,145,0,235,0,0,0,114,0,68,0,58,0,204,0,109,0,0,0,105,0,181,0,77,0,254,0,0,0,1,0,180,0,18,0,76,0,78,0,241,0,0,0,59,0,255,0,101,0,48,0,124,0,0,0,130,0,208,0,221,0,220,0,132,0,0,0,32,0,227,0,152,0,0,0,161,0,173,0,175,0,160,0,177,0,143,0,135,0,0,0,111,0,0,0,246,0,252,0,0,0,147,0,0,0,47,0,194,0,220,0,12,0,87,0,178,0,197,0,43,0,60,0,163,0,220,0,173,0,183,0,146,0,244,0,198,0,76,0,106,0,184,0,0,0,179,0,24,0,167,0,7,0,0,0,234,0,43,0,241,0,95,0,180,0,71,0,49,0,138,0,119,0,137,0,27,0,180,0,0,0,0,0,88,0,0,0,68,0,79,0,0,0,245,0,119,0,95,0,0,0,177,0,11,0,9,0,95,0,178,0,183,0,89,0,136,0,139,0,222,0,128,0,95,0,127,0,118,0,213,0,147,0,135,0,15,0,35,0,240,0,28,0,74,0,164,0,24,0,81,0,157,0,0,0,12,0,0,0,67,0,243,0,44,0,136,0,130,0,155,0,69,0,52,0,10,0,24,0,48,0,75,0,0,0,110,0,117,0,135,0,148,0,0,0,171,0,43,0,209,0,128,0,28,0,0,0,170,0,194,0,36,0,227,0,126,0,247,0,0,0,21,0);
signal scenario_full  : scenario_type := (238,31,238,30,166,31,153,31,225,31,63,31,52,31,111,31,111,30,111,29,226,31,141,31,68,31,164,31,158,31,158,30,48,31,180,31,181,31,120,31,33,31,232,31,169,31,169,30,85,31,189,31,77,31,3,31,50,31,145,31,53,31,102,31,185,31,120,31,41,31,226,31,232,31,232,30,177,31,85,31,231,31,231,30,145,31,235,31,235,30,114,31,68,31,58,31,204,31,109,31,109,30,105,31,181,31,77,31,254,31,254,30,1,31,180,31,18,31,76,31,78,31,241,31,241,30,59,31,255,31,101,31,48,31,124,31,124,30,130,31,208,31,221,31,220,31,132,31,132,30,32,31,227,31,152,31,152,30,161,31,173,31,175,31,160,31,177,31,143,31,135,31,135,30,111,31,111,30,246,31,252,31,252,30,147,31,147,30,47,31,194,31,220,31,12,31,87,31,178,31,197,31,43,31,60,31,163,31,220,31,173,31,183,31,146,31,244,31,198,31,76,31,106,31,184,31,184,30,179,31,24,31,167,31,7,31,7,30,234,31,43,31,241,31,95,31,180,31,71,31,49,31,138,31,119,31,137,31,27,31,180,31,180,30,180,29,88,31,88,30,68,31,79,31,79,30,245,31,119,31,95,31,95,30,177,31,11,31,9,31,95,31,178,31,183,31,89,31,136,31,139,31,222,31,128,31,95,31,127,31,118,31,213,31,147,31,135,31,15,31,35,31,240,31,28,31,74,31,164,31,24,31,81,31,157,31,157,30,12,31,12,30,67,31,243,31,44,31,136,31,130,31,155,31,69,31,52,31,10,31,24,31,48,31,75,31,75,30,110,31,117,31,135,31,148,31,148,30,171,31,43,31,209,31,128,31,28,31,28,30,170,31,194,31,36,31,227,31,126,31,247,31,247,30,21,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
