-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_498 is
end project_tb_498;

architecture project_tb_arch_498 of project_tb_498 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 898;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (36,0,159,0,97,0,100,0,0,0,54,0,239,0,128,0,151,0,128,0,100,0,115,0,131,0,225,0,59,0,207,0,10,0,41,0,179,0,227,0,7,0,39,0,252,0,248,0,54,0,150,0,115,0,173,0,139,0,255,0,73,0,56,0,31,0,229,0,179,0,155,0,141,0,19,0,194,0,44,0,137,0,2,0,102,0,220,0,173,0,16,0,0,0,191,0,0,0,115,0,40,0,115,0,165,0,173,0,241,0,218,0,218,0,219,0,232,0,16,0,204,0,0,0,115,0,92,0,31,0,0,0,82,0,52,0,81,0,0,0,140,0,19,0,161,0,0,0,227,0,27,0,112,0,110,0,254,0,0,0,5,0,56,0,68,0,145,0,78,0,0,0,33,0,218,0,0,0,54,0,76,0,210,0,233,0,12,0,99,0,0,0,19,0,0,0,36,0,0,0,0,0,194,0,0,0,21,0,95,0,152,0,7,0,175,0,194,0,233,0,174,0,117,0,41,0,155,0,20,0,0,0,0,0,125,0,162,0,56,0,73,0,210,0,106,0,27,0,39,0,216,0,237,0,3,0,253,0,19,0,6,0,245,0,19,0,47,0,88,0,137,0,120,0,0,0,63,0,0,0,177,0,0,0,0,0,124,0,0,0,0,0,207,0,0,0,222,0,0,0,83,0,87,0,173,0,176,0,106,0,220,0,30,0,181,0,247,0,234,0,198,0,0,0,108,0,238,0,34,0,0,0,214,0,133,0,3,0,187,0,227,0,3,0,64,0,0,0,0,0,0,0,0,0,106,0,174,0,139,0,86,0,209,0,82,0,154,0,0,0,66,0,155,0,191,0,162,0,0,0,194,0,0,0,0,0,70,0,127,0,107,0,59,0,239,0,236,0,45,0,167,0,178,0,164,0,0,0,191,0,239,0,41,0,31,0,150,0,53,0,0,0,115,0,144,0,190,0,24,0,50,0,247,0,126,0,30,0,0,0,0,0,119,0,0,0,246,0,0,0,87,0,195,0,218,0,0,0,218,0,178,0,0,0,123,0,104,0,0,0,112,0,125,0,82,0,0,0,129,0,0,0,112,0,144,0,30,0,234,0,0,0,64,0,249,0,189,0,103,0,112,0,188,0,199,0,0,0,182,0,0,0,0,0,246,0,211,0,119,0,228,0,172,0,182,0,242,0,168,0,0,0,168,0,24,0,0,0,247,0,177,0,62,0,12,0,0,0,0,0,155,0,79,0,96,0,103,0,201,0,83,0,126,0,178,0,109,0,131,0,38,0,153,0,34,0,0,0,15,0,168,0,105,0,144,0,78,0,34,0,0,0,0,0,156,0,0,0,64,0,250,0,7,0,0,0,61,0,0,0,143,0,168,0,0,0,68,0,92,0,62,0,138,0,18,0,38,0,66,0,0,0,0,0,0,0,150,0,0,0,1,0,0,0,221,0,169,0,211,0,0,0,203,0,0,0,130,0,0,0,2,0,55,0,102,0,232,0,26,0,0,0,0,0,30,0,166,0,37,0,244,0,166,0,0,0,107,0,216,0,0,0,218,0,209,0,0,0,0,0,0,0,192,0,88,0,104,0,0,0,0,0,50,0,80,0,25,0,5,0,245,0,174,0,7,0,72,0,27,0,0,0,0,0,52,0,0,0,33,0,6,0,210,0,0,0,202,0,244,0,34,0,0,0,79,0,0,0,0,0,145,0,0,0,0,0,94,0,97,0,211,0,70,0,174,0,43,0,121,0,79,0,177,0,179,0,0,0,0,0,126,0,123,0,173,0,150,0,0,0,251,0,0,0,43,0,242,0,148,0,202,0,15,0,211,0,250,0,66,0,57,0,229,0,222,0,68,0,60,0,112,0,187,0,159,0,125,0,193,0,123,0,0,0,196,0,184,0,138,0,0,0,39,0,129,0,168,0,0,0,54,0,102,0,254,0,0,0,123,0,0,0,236,0,151,0,199,0,41,0,252,0,50,0,82,0,230,0,168,0,100,0,125,0,0,0,0,0,234,0,84,0,237,0,149,0,94,0,0,0,0,0,116,0,54,0,224,0,140,0,254,0,13,0,173,0,76,0,18,0,73,0,0,0,110,0,57,0,132,0,207,0,0,0,144,0,153,0,114,0,55,0,0,0,252,0,0,0,200,0,38,0,238,0,0,0,181,0,211,0,113,0,163,0,25,0,200,0,251,0,209,0,16,0,37,0,0,0,164,0,16,0,96,0,72,0,157,0,119,0,0,0,0,0,0,0,33,0,22,0,142,0,156,0,252,0,83,0,224,0,241,0,166,0,169,0,143,0,97,0,215,0,90,0,221,0,115,0,14,0,74,0,0,0,0,0,66,0,22,0,221,0,233,0,205,0,184,0,3,0,0,0,0,0,132,0,0,0,180,0,165,0,18,0,87,0,0,0,101,0,100,0,217,0,0,0,142,0,32,0,229,0,250,0,131,0,73,0,112,0,233,0,14,0,24,0,0,0,0,0,0,0,84,0,142,0,127,0,123,0,4,0,65,0,0,0,86,0,112,0,222,0,173,0,32,0,248,0,58,0,253,0,10,0,0,0,226,0,0,0,0,0,0,0,82,0,64,0,82,0,0,0,231,0,0,0,53,0,102,0,104,0,137,0,14,0,143,0,171,0,200,0,55,0,0,0,2,0,84,0,244,0,223,0,237,0,105,0,0,0,2,0,46,0,72,0,101,0,90,0,0,0,0,0,44,0,232,0,219,0,155,0,41,0,0,0,25,0,170,0,20,0,182,0,53,0,176,0,154,0,74,0,0,0,0,0,223,0,0,0,0,0,232,0,129,0,39,0,49,0,161,0,8,0,168,0,204,0,200,0,125,0,251,0,0,0,0,0,90,0,21,0,185,0,248,0,149,0,166,0,205,0,0,0,0,0,154,0,81,0,239,0,51,0,78,0,12,0,164,0,99,0,215,0,135,0,0,0,188,0,41,0,24,0,220,0,18,0,252,0,23,0,199,0,199,0,0,0,146,0,68,0,0,0,84,0,175,0,171,0,192,0,51,0,102,0,33,0,200,0,3,0,0,0,193,0,57,0,110,0,0,0,0,0,129,0,0,0,0,0,18,0,127,0,246,0,231,0,153,0,1,0,236,0,0,0,248,0,2,0,48,0,41,0,0,0,164,0,108,0,8,0,0,0,200,0,240,0,189,0,226,0,104,0,111,0,226,0,246,0,0,0,18,0,128,0,0,0,112,0,162,0,12,0,122,0,40,0,14,0,63,0,32,0,219,0,84,0,178,0,0,0,0,0,53,0,146,0,125,0,122,0,51,0,0,0,0,0,183,0,97,0,109,0,0,0,146,0,46,0,225,0,106,0,185,0,130,0,247,0,184,0,0,0,204,0,60,0,0,0,128,0,159,0,121,0,134,0,128,0,188,0,20,0,111,0,0,0,199,0,82,0,191,0,0,0,17,0,20,0,97,0,198,0,128,0,110,0,124,0,102,0,82,0,241,0,21,0,130,0,129,0,6,0,184,0,128,0,102,0,4,0,217,0,43,0,163,0,131,0,17,0,0,0,81,0,239,0,242,0,253,0,219,0,42,0,201,0,142,0,156,0,235,0,176,0,211,0,156,0,137,0,107,0,212,0,0,0,40,0,0,0,130,0,200,0,195,0,0,0,0,0,251,0,233,0,126,0,0,0,32,0,0,0,219,0,54,0,253,0,45,0,0,0,0,0,190,0,99,0,226,0,221,0,98,0,202,0,162,0,137,0,149,0,0,0,230,0,205,0,139,0,0,0,0,0,162,0,78,0,173,0,31,0,160,0,0,0,183,0,102,0,156,0,230,0,66,0,71,0,120,0,250,0,12,0,134,0,112,0,153,0,211,0,39,0,76,0,0,0,221,0,35,0,27,0,139,0,2,0,187,0,0,0,0,0,132,0,0,0,244,0,57,0,35,0,92,0,165,0,0,0,212,0,31,0,0,0,97,0,98,0,0,0,0,0,33,0,87,0,127,0,107,0,2,0,221,0,192,0,246,0,35,0,0,0);
signal scenario_full  : scenario_type := (36,31,159,31,97,31,100,31,100,30,54,31,239,31,128,31,151,31,128,31,100,31,115,31,131,31,225,31,59,31,207,31,10,31,41,31,179,31,227,31,7,31,39,31,252,31,248,31,54,31,150,31,115,31,173,31,139,31,255,31,73,31,56,31,31,31,229,31,179,31,155,31,141,31,19,31,194,31,44,31,137,31,2,31,102,31,220,31,173,31,16,31,16,30,191,31,191,30,115,31,40,31,115,31,165,31,173,31,241,31,218,31,218,31,219,31,232,31,16,31,204,31,204,30,115,31,92,31,31,31,31,30,82,31,52,31,81,31,81,30,140,31,19,31,161,31,161,30,227,31,27,31,112,31,110,31,254,31,254,30,5,31,56,31,68,31,145,31,78,31,78,30,33,31,218,31,218,30,54,31,76,31,210,31,233,31,12,31,99,31,99,30,19,31,19,30,36,31,36,30,36,29,194,31,194,30,21,31,95,31,152,31,7,31,175,31,194,31,233,31,174,31,117,31,41,31,155,31,20,31,20,30,20,29,125,31,162,31,56,31,73,31,210,31,106,31,27,31,39,31,216,31,237,31,3,31,253,31,19,31,6,31,245,31,19,31,47,31,88,31,137,31,120,31,120,30,63,31,63,30,177,31,177,30,177,29,124,31,124,30,124,29,207,31,207,30,222,31,222,30,83,31,87,31,173,31,176,31,106,31,220,31,30,31,181,31,247,31,234,31,198,31,198,30,108,31,238,31,34,31,34,30,214,31,133,31,3,31,187,31,227,31,3,31,64,31,64,30,64,29,64,28,64,27,106,31,174,31,139,31,86,31,209,31,82,31,154,31,154,30,66,31,155,31,191,31,162,31,162,30,194,31,194,30,194,29,70,31,127,31,107,31,59,31,239,31,236,31,45,31,167,31,178,31,164,31,164,30,191,31,239,31,41,31,31,31,150,31,53,31,53,30,115,31,144,31,190,31,24,31,50,31,247,31,126,31,30,31,30,30,30,29,119,31,119,30,246,31,246,30,87,31,195,31,218,31,218,30,218,31,178,31,178,30,123,31,104,31,104,30,112,31,125,31,82,31,82,30,129,31,129,30,112,31,144,31,30,31,234,31,234,30,64,31,249,31,189,31,103,31,112,31,188,31,199,31,199,30,182,31,182,30,182,29,246,31,211,31,119,31,228,31,172,31,182,31,242,31,168,31,168,30,168,31,24,31,24,30,247,31,177,31,62,31,12,31,12,30,12,29,155,31,79,31,96,31,103,31,201,31,83,31,126,31,178,31,109,31,131,31,38,31,153,31,34,31,34,30,15,31,168,31,105,31,144,31,78,31,34,31,34,30,34,29,156,31,156,30,64,31,250,31,7,31,7,30,61,31,61,30,143,31,168,31,168,30,68,31,92,31,62,31,138,31,18,31,38,31,66,31,66,30,66,29,66,28,150,31,150,30,1,31,1,30,221,31,169,31,211,31,211,30,203,31,203,30,130,31,130,30,2,31,55,31,102,31,232,31,26,31,26,30,26,29,30,31,166,31,37,31,244,31,166,31,166,30,107,31,216,31,216,30,218,31,209,31,209,30,209,29,209,28,192,31,88,31,104,31,104,30,104,29,50,31,80,31,25,31,5,31,245,31,174,31,7,31,72,31,27,31,27,30,27,29,52,31,52,30,33,31,6,31,210,31,210,30,202,31,244,31,34,31,34,30,79,31,79,30,79,29,145,31,145,30,145,29,94,31,97,31,211,31,70,31,174,31,43,31,121,31,79,31,177,31,179,31,179,30,179,29,126,31,123,31,173,31,150,31,150,30,251,31,251,30,43,31,242,31,148,31,202,31,15,31,211,31,250,31,66,31,57,31,229,31,222,31,68,31,60,31,112,31,187,31,159,31,125,31,193,31,123,31,123,30,196,31,184,31,138,31,138,30,39,31,129,31,168,31,168,30,54,31,102,31,254,31,254,30,123,31,123,30,236,31,151,31,199,31,41,31,252,31,50,31,82,31,230,31,168,31,100,31,125,31,125,30,125,29,234,31,84,31,237,31,149,31,94,31,94,30,94,29,116,31,54,31,224,31,140,31,254,31,13,31,173,31,76,31,18,31,73,31,73,30,110,31,57,31,132,31,207,31,207,30,144,31,153,31,114,31,55,31,55,30,252,31,252,30,200,31,38,31,238,31,238,30,181,31,211,31,113,31,163,31,25,31,200,31,251,31,209,31,16,31,37,31,37,30,164,31,16,31,96,31,72,31,157,31,119,31,119,30,119,29,119,28,33,31,22,31,142,31,156,31,252,31,83,31,224,31,241,31,166,31,169,31,143,31,97,31,215,31,90,31,221,31,115,31,14,31,74,31,74,30,74,29,66,31,22,31,221,31,233,31,205,31,184,31,3,31,3,30,3,29,132,31,132,30,180,31,165,31,18,31,87,31,87,30,101,31,100,31,217,31,217,30,142,31,32,31,229,31,250,31,131,31,73,31,112,31,233,31,14,31,24,31,24,30,24,29,24,28,84,31,142,31,127,31,123,31,4,31,65,31,65,30,86,31,112,31,222,31,173,31,32,31,248,31,58,31,253,31,10,31,10,30,226,31,226,30,226,29,226,28,82,31,64,31,82,31,82,30,231,31,231,30,53,31,102,31,104,31,137,31,14,31,143,31,171,31,200,31,55,31,55,30,2,31,84,31,244,31,223,31,237,31,105,31,105,30,2,31,46,31,72,31,101,31,90,31,90,30,90,29,44,31,232,31,219,31,155,31,41,31,41,30,25,31,170,31,20,31,182,31,53,31,176,31,154,31,74,31,74,30,74,29,223,31,223,30,223,29,232,31,129,31,39,31,49,31,161,31,8,31,168,31,204,31,200,31,125,31,251,31,251,30,251,29,90,31,21,31,185,31,248,31,149,31,166,31,205,31,205,30,205,29,154,31,81,31,239,31,51,31,78,31,12,31,164,31,99,31,215,31,135,31,135,30,188,31,41,31,24,31,220,31,18,31,252,31,23,31,199,31,199,31,199,30,146,31,68,31,68,30,84,31,175,31,171,31,192,31,51,31,102,31,33,31,200,31,3,31,3,30,193,31,57,31,110,31,110,30,110,29,129,31,129,30,129,29,18,31,127,31,246,31,231,31,153,31,1,31,236,31,236,30,248,31,2,31,48,31,41,31,41,30,164,31,108,31,8,31,8,30,200,31,240,31,189,31,226,31,104,31,111,31,226,31,246,31,246,30,18,31,128,31,128,30,112,31,162,31,12,31,122,31,40,31,14,31,63,31,32,31,219,31,84,31,178,31,178,30,178,29,53,31,146,31,125,31,122,31,51,31,51,30,51,29,183,31,97,31,109,31,109,30,146,31,46,31,225,31,106,31,185,31,130,31,247,31,184,31,184,30,204,31,60,31,60,30,128,31,159,31,121,31,134,31,128,31,188,31,20,31,111,31,111,30,199,31,82,31,191,31,191,30,17,31,20,31,97,31,198,31,128,31,110,31,124,31,102,31,82,31,241,31,21,31,130,31,129,31,6,31,184,31,128,31,102,31,4,31,217,31,43,31,163,31,131,31,17,31,17,30,81,31,239,31,242,31,253,31,219,31,42,31,201,31,142,31,156,31,235,31,176,31,211,31,156,31,137,31,107,31,212,31,212,30,40,31,40,30,130,31,200,31,195,31,195,30,195,29,251,31,233,31,126,31,126,30,32,31,32,30,219,31,54,31,253,31,45,31,45,30,45,29,190,31,99,31,226,31,221,31,98,31,202,31,162,31,137,31,149,31,149,30,230,31,205,31,139,31,139,30,139,29,162,31,78,31,173,31,31,31,160,31,160,30,183,31,102,31,156,31,230,31,66,31,71,31,120,31,250,31,12,31,134,31,112,31,153,31,211,31,39,31,76,31,76,30,221,31,35,31,27,31,139,31,2,31,187,31,187,30,187,29,132,31,132,30,244,31,57,31,35,31,92,31,165,31,165,30,212,31,31,31,31,30,97,31,98,31,98,30,98,29,33,31,87,31,127,31,107,31,2,31,221,31,192,31,246,31,35,31,35,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
