-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_424 is
end project_tb_424;

architecture project_tb_arch_424 of project_tb_424 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 800;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (125,0,184,0,194,0,164,0,8,0,139,0,204,0,165,0,98,0,128,0,78,0,0,0,78,0,0,0,195,0,172,0,249,0,234,0,0,0,227,0,0,0,111,0,19,0,191,0,57,0,0,0,45,0,251,0,238,0,110,0,72,0,129,0,226,0,0,0,252,0,162,0,21,0,214,0,46,0,65,0,201,0,127,0,0,0,82,0,0,0,200,0,25,0,0,0,121,0,31,0,236,0,163,0,0,0,136,0,0,0,1,0,63,0,0,0,241,0,247,0,147,0,1,0,192,0,230,0,141,0,0,0,41,0,163,0,4,0,99,0,34,0,29,0,249,0,168,0,5,0,7,0,0,0,206,0,45,0,142,0,75,0,0,0,17,0,32,0,0,0,166,0,0,0,55,0,0,0,91,0,0,0,81,0,0,0,253,0,243,0,181,0,124,0,139,0,23,0,173,0,138,0,177,0,197,0,130,0,0,0,168,0,6,0,17,0,130,0,145,0,104,0,42,0,34,0,196,0,238,0,0,0,84,0,53,0,78,0,146,0,132,0,222,0,123,0,40,0,127,0,251,0,42,0,64,0,201,0,96,0,6,0,141,0,244,0,129,0,145,0,243,0,48,0,54,0,54,0,33,0,137,0,139,0,0,0,0,0,0,0,79,0,24,0,36,0,0,0,208,0,222,0,131,0,159,0,0,0,16,0,251,0,134,0,232,0,75,0,163,0,125,0,90,0,0,0,146,0,143,0,6,0,241,0,0,0,64,0,244,0,199,0,32,0,186,0,224,0,154,0,251,0,36,0,42,0,59,0,202,0,107,0,162,0,122,0,0,0,229,0,0,0,61,0,57,0,131,0,65,0,26,0,31,0,0,0,2,0,28,0,92,0,140,0,62,0,0,0,238,0,188,0,246,0,0,0,162,0,0,0,29,0,137,0,128,0,22,0,176,0,144,0,197,0,172,0,41,0,107,0,222,0,83,0,44,0,188,0,152,0,13,0,33,0,88,0,46,0,166,0,107,0,128,0,199,0,160,0,235,0,0,0,103,0,246,0,121,0,114,0,130,0,172,0,22,0,23,0,0,0,31,0,16,0,247,0,0,0,18,0,177,0,161,0,202,0,35,0,35,0,83,0,0,0,0,0,80,0,103,0,175,0,0,0,129,0,0,0,129,0,110,0,249,0,45,0,51,0,12,0,105,0,227,0,1,0,0,0,151,0,252,0,127,0,0,0,95,0,0,0,0,0,13,0,123,0,184,0,0,0,22,0,25,0,190,0,160,0,87,0,37,0,54,0,205,0,153,0,4,0,38,0,245,0,42,0,103,0,121,0,161,0,123,0,211,0,37,0,99,0,64,0,30,0,46,0,226,0,160,0,206,0,219,0,247,0,22,0,239,0,42,0,0,0,0,0,36,0,0,0,195,0,171,0,237,0,99,0,136,0,27,0,114,0,240,0,27,0,0,0,160,0,68,0,0,0,207,0,0,0,0,0,67,0,0,0,186,0,102,0,233,0,228,0,146,0,200,0,203,0,26,0,190,0,132,0,17,0,137,0,38,0,0,0,7,0,230,0,146,0,0,0,157,0,76,0,252,0,10,0,60,0,128,0,215,0,0,0,79,0,0,0,0,0,0,0,0,0,135,0,169,0,61,0,115,0,183,0,0,0,232,0,0,0,0,0,123,0,124,0,0,0,77,0,105,0,120,0,0,0,0,0,77,0,170,0,239,0,52,0,236,0,160,0,71,0,0,0,86,0,0,0,204,0,226,0,114,0,43,0,106,0,68,0,22,0,211,0,206,0,15,0,31,0,206,0,0,0,34,0,0,0,12,0,161,0,214,0,114,0,0,0,60,0,117,0,133,0,208,0,242,0,236,0,252,0,204,0,172,0,118,0,148,0,0,0,178,0,0,0,72,0,195,0,209,0,111,0,151,0,81,0,206,0,210,0,30,0,0,0,0,0,29,0,86,0,167,0,103,0,172,0,0,0,75,0,0,0,133,0,254,0,0,0,220,0,158,0,230,0,255,0,92,0,3,0,27,0,0,0,157,0,0,0,0,0,198,0,79,0,0,0,196,0,11,0,149,0,0,0,4,0,144,0,0,0,88,0,233,0,188,0,252,0,0,0,145,0,0,0,138,0,176,0,68,0,9,0,0,0,229,0,34,0,19,0,25,0,51,0,46,0,144,0,0,0,214,0,208,0,151,0,203,0,145,0,0,0,203,0,198,0,195,0,129,0,148,0,0,0,206,0,65,0,33,0,218,0,196,0,209,0,123,0,227,0,16,0,0,0,188,0,160,0,5,0,30,0,27,0,39,0,225,0,130,0,49,0,28,0,222,0,74,0,132,0,162,0,72,0,164,0,185,0,173,0,99,0,59,0,0,0,173,0,85,0,63,0,69,0,60,0,32,0,69,0,7,0,246,0,183,0,0,0,0,0,0,0,0,0,0,0,199,0,6,0,241,0,235,0,38,0,244,0,220,0,0,0,241,0,40,0,4,0,0,0,157,0,0,0,99,0,179,0,197,0,98,0,196,0,0,0,208,0,0,0,54,0,0,0,0,0,74,0,0,0,8,0,214,0,37,0,0,0,241,0,0,0,247,0,44,0,210,0,158,0,0,0,173,0,172,0,70,0,11,0,76,0,8,0,121,0,251,0,156,0,0,0,34,0,89,0,107,0,203,0,0,0,149,0,98,0,207,0,0,0,98,0,206,0,145,0,20,0,146,0,0,0,9,0,12,0,140,0,218,0,134,0,233,0,183,0,0,0,40,0,82,0,122,0,64,0,111,0,130,0,45,0,142,0,78,0,145,0,143,0,247,0,195,0,233,0,226,0,233,0,95,0,195,0,201,0,193,0,39,0,0,0,0,0,0,0,103,0,245,0,135,0,176,0,0,0,138,0,223,0,221,0,203,0,80,0,54,0,129,0,163,0,183,0,3,0,59,0,150,0,116,0,134,0,58,0,207,0,76,0,90,0,0,0,125,0,29,0,147,0,185,0,0,0,183,0,5,0,94,0,228,0,244,0,146,0,15,0,73,0,10,0,100,0,31,0,210,0,0,0,0,0,0,0,136,0,37,0,168,0,227,0,73,0,230,0,55,0,14,0,189,0,46,0,97,0,0,0,0,0,133,0,0,0,64,0,236,0,0,0,0,0,211,0,0,0,163,0,193,0,0,0,203,0,217,0,13,0,234,0,70,0,90,0,0,0,13,0,144,0,0,0,223,0,0,0,204,0,249,0,165,0,237,0,65,0,66,0,113,0,108,0,0,0,247,0,177,0,228,0,146,0,136,0,46,0,251,0,17,0,0,0,65,0,95,0,210,0,50,0,228,0,196,0,0,0,0,0,45,0,0,0,42,0,0,0,222,0,43,0,244,0,90,0,222,0,22,0,17,0,225,0,216,0,187,0,0,0,39,0,230,0,40,0,123,0,0,0,246,0,118,0,149,0,151,0,0,0,181,0,0,0,178,0,251,0,0,0,157,0,108,0,0,0,0,0,215,0,183,0,232,0,245,0,0,0,22,0,0,0,179,0,0,0,61,0,5,0,167,0,218,0,183,0,69,0,74,0,119,0,0,0,134,0);
signal scenario_full  : scenario_type := (125,31,184,31,194,31,164,31,8,31,139,31,204,31,165,31,98,31,128,31,78,31,78,30,78,31,78,30,195,31,172,31,249,31,234,31,234,30,227,31,227,30,111,31,19,31,191,31,57,31,57,30,45,31,251,31,238,31,110,31,72,31,129,31,226,31,226,30,252,31,162,31,21,31,214,31,46,31,65,31,201,31,127,31,127,30,82,31,82,30,200,31,25,31,25,30,121,31,31,31,236,31,163,31,163,30,136,31,136,30,1,31,63,31,63,30,241,31,247,31,147,31,1,31,192,31,230,31,141,31,141,30,41,31,163,31,4,31,99,31,34,31,29,31,249,31,168,31,5,31,7,31,7,30,206,31,45,31,142,31,75,31,75,30,17,31,32,31,32,30,166,31,166,30,55,31,55,30,91,31,91,30,81,31,81,30,253,31,243,31,181,31,124,31,139,31,23,31,173,31,138,31,177,31,197,31,130,31,130,30,168,31,6,31,17,31,130,31,145,31,104,31,42,31,34,31,196,31,238,31,238,30,84,31,53,31,78,31,146,31,132,31,222,31,123,31,40,31,127,31,251,31,42,31,64,31,201,31,96,31,6,31,141,31,244,31,129,31,145,31,243,31,48,31,54,31,54,31,33,31,137,31,139,31,139,30,139,29,139,28,79,31,24,31,36,31,36,30,208,31,222,31,131,31,159,31,159,30,16,31,251,31,134,31,232,31,75,31,163,31,125,31,90,31,90,30,146,31,143,31,6,31,241,31,241,30,64,31,244,31,199,31,32,31,186,31,224,31,154,31,251,31,36,31,42,31,59,31,202,31,107,31,162,31,122,31,122,30,229,31,229,30,61,31,57,31,131,31,65,31,26,31,31,31,31,30,2,31,28,31,92,31,140,31,62,31,62,30,238,31,188,31,246,31,246,30,162,31,162,30,29,31,137,31,128,31,22,31,176,31,144,31,197,31,172,31,41,31,107,31,222,31,83,31,44,31,188,31,152,31,13,31,33,31,88,31,46,31,166,31,107,31,128,31,199,31,160,31,235,31,235,30,103,31,246,31,121,31,114,31,130,31,172,31,22,31,23,31,23,30,31,31,16,31,247,31,247,30,18,31,177,31,161,31,202,31,35,31,35,31,83,31,83,30,83,29,80,31,103,31,175,31,175,30,129,31,129,30,129,31,110,31,249,31,45,31,51,31,12,31,105,31,227,31,1,31,1,30,151,31,252,31,127,31,127,30,95,31,95,30,95,29,13,31,123,31,184,31,184,30,22,31,25,31,190,31,160,31,87,31,37,31,54,31,205,31,153,31,4,31,38,31,245,31,42,31,103,31,121,31,161,31,123,31,211,31,37,31,99,31,64,31,30,31,46,31,226,31,160,31,206,31,219,31,247,31,22,31,239,31,42,31,42,30,42,29,36,31,36,30,195,31,171,31,237,31,99,31,136,31,27,31,114,31,240,31,27,31,27,30,160,31,68,31,68,30,207,31,207,30,207,29,67,31,67,30,186,31,102,31,233,31,228,31,146,31,200,31,203,31,26,31,190,31,132,31,17,31,137,31,38,31,38,30,7,31,230,31,146,31,146,30,157,31,76,31,252,31,10,31,60,31,128,31,215,31,215,30,79,31,79,30,79,29,79,28,79,27,135,31,169,31,61,31,115,31,183,31,183,30,232,31,232,30,232,29,123,31,124,31,124,30,77,31,105,31,120,31,120,30,120,29,77,31,170,31,239,31,52,31,236,31,160,31,71,31,71,30,86,31,86,30,204,31,226,31,114,31,43,31,106,31,68,31,22,31,211,31,206,31,15,31,31,31,206,31,206,30,34,31,34,30,12,31,161,31,214,31,114,31,114,30,60,31,117,31,133,31,208,31,242,31,236,31,252,31,204,31,172,31,118,31,148,31,148,30,178,31,178,30,72,31,195,31,209,31,111,31,151,31,81,31,206,31,210,31,30,31,30,30,30,29,29,31,86,31,167,31,103,31,172,31,172,30,75,31,75,30,133,31,254,31,254,30,220,31,158,31,230,31,255,31,92,31,3,31,27,31,27,30,157,31,157,30,157,29,198,31,79,31,79,30,196,31,11,31,149,31,149,30,4,31,144,31,144,30,88,31,233,31,188,31,252,31,252,30,145,31,145,30,138,31,176,31,68,31,9,31,9,30,229,31,34,31,19,31,25,31,51,31,46,31,144,31,144,30,214,31,208,31,151,31,203,31,145,31,145,30,203,31,198,31,195,31,129,31,148,31,148,30,206,31,65,31,33,31,218,31,196,31,209,31,123,31,227,31,16,31,16,30,188,31,160,31,5,31,30,31,27,31,39,31,225,31,130,31,49,31,28,31,222,31,74,31,132,31,162,31,72,31,164,31,185,31,173,31,99,31,59,31,59,30,173,31,85,31,63,31,69,31,60,31,32,31,69,31,7,31,246,31,183,31,183,30,183,29,183,28,183,27,183,26,199,31,6,31,241,31,235,31,38,31,244,31,220,31,220,30,241,31,40,31,4,31,4,30,157,31,157,30,99,31,179,31,197,31,98,31,196,31,196,30,208,31,208,30,54,31,54,30,54,29,74,31,74,30,8,31,214,31,37,31,37,30,241,31,241,30,247,31,44,31,210,31,158,31,158,30,173,31,172,31,70,31,11,31,76,31,8,31,121,31,251,31,156,31,156,30,34,31,89,31,107,31,203,31,203,30,149,31,98,31,207,31,207,30,98,31,206,31,145,31,20,31,146,31,146,30,9,31,12,31,140,31,218,31,134,31,233,31,183,31,183,30,40,31,82,31,122,31,64,31,111,31,130,31,45,31,142,31,78,31,145,31,143,31,247,31,195,31,233,31,226,31,233,31,95,31,195,31,201,31,193,31,39,31,39,30,39,29,39,28,103,31,245,31,135,31,176,31,176,30,138,31,223,31,221,31,203,31,80,31,54,31,129,31,163,31,183,31,3,31,59,31,150,31,116,31,134,31,58,31,207,31,76,31,90,31,90,30,125,31,29,31,147,31,185,31,185,30,183,31,5,31,94,31,228,31,244,31,146,31,15,31,73,31,10,31,100,31,31,31,210,31,210,30,210,29,210,28,136,31,37,31,168,31,227,31,73,31,230,31,55,31,14,31,189,31,46,31,97,31,97,30,97,29,133,31,133,30,64,31,236,31,236,30,236,29,211,31,211,30,163,31,193,31,193,30,203,31,217,31,13,31,234,31,70,31,90,31,90,30,13,31,144,31,144,30,223,31,223,30,204,31,249,31,165,31,237,31,65,31,66,31,113,31,108,31,108,30,247,31,177,31,228,31,146,31,136,31,46,31,251,31,17,31,17,30,65,31,95,31,210,31,50,31,228,31,196,31,196,30,196,29,45,31,45,30,42,31,42,30,222,31,43,31,244,31,90,31,222,31,22,31,17,31,225,31,216,31,187,31,187,30,39,31,230,31,40,31,123,31,123,30,246,31,118,31,149,31,151,31,151,30,181,31,181,30,178,31,251,31,251,30,157,31,108,31,108,30,108,29,215,31,183,31,232,31,245,31,245,30,22,31,22,30,179,31,179,30,61,31,5,31,167,31,218,31,183,31,69,31,74,31,119,31,119,30,134,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
