-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_671 is
end project_tb_671;

architecture project_tb_arch_671 of project_tb_671 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 652;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,56,0,52,0,0,0,249,0,0,0,44,0,166,0,0,0,239,0,173,0,34,0,252,0,0,0,136,0,0,0,168,0,37,0,34,0,128,0,33,0,48,0,8,0,190,0,110,0,48,0,56,0,188,0,46,0,36,0,216,0,0,0,0,0,162,0,213,0,194,0,0,0,68,0,0,0,131,0,0,0,41,0,212,0,214,0,248,0,14,0,53,0,107,0,0,0,0,0,83,0,0,0,0,0,52,0,235,0,199,0,199,0,38,0,238,0,0,0,0,0,136,0,17,0,53,0,225,0,209,0,149,0,0,0,132,0,204,0,231,0,0,0,125,0,45,0,0,0,0,0,56,0,150,0,208,0,209,0,169,0,72,0,127,0,191,0,99,0,235,0,168,0,207,0,173,0,33,0,67,0,131,0,143,0,81,0,61,0,0,0,219,0,131,0,181,0,26,0,14,0,175,0,45,0,0,0,6,0,30,0,97,0,0,0,34,0,40,0,248,0,95,0,187,0,107,0,230,0,40,0,0,0,80,0,194,0,214,0,168,0,153,0,236,0,230,0,0,0,185,0,34,0,0,0,0,0,0,0,56,0,0,0,61,0,230,0,126,0,244,0,215,0,63,0,67,0,0,0,21,0,178,0,135,0,153,0,37,0,86,0,85,0,148,0,216,0,199,0,83,0,46,0,190,0,133,0,150,0,28,0,243,0,119,0,0,0,86,0,0,0,5,0,26,0,0,0,230,0,231,0,237,0,117,0,149,0,0,0,23,0,140,0,88,0,156,0,180,0,78,0,0,0,127,0,7,0,205,0,0,0,111,0,150,0,0,0,103,0,147,0,0,0,0,0,107,0,0,0,147,0,51,0,106,0,157,0,29,0,235,0,245,0,169,0,116,0,0,0,77,0,15,0,200,0,220,0,206,0,0,0,182,0,100,0,0,0,157,0,23,0,171,0,176,0,47,0,18,0,141,0,127,0,175,0,56,0,212,0,60,0,111,0,0,0,5,0,130,0,0,0,250,0,144,0,0,0,241,0,85,0,212,0,227,0,70,0,120,0,80,0,136,0,0,0,0,0,27,0,11,0,0,0,167,0,33,0,85,0,0,0,207,0,196,0,25,0,20,0,11,0,108,0,0,0,105,0,207,0,242,0,0,0,203,0,63,0,0,0,0,0,91,0,58,0,219,0,0,0,0,0,242,0,0,0,139,0,0,0,0,0,23,0,121,0,40,0,172,0,232,0,11,0,148,0,137,0,184,0,28,0,105,0,93,0,98,0,34,0,0,0,0,0,103,0,7,0,26,0,0,0,92,0,0,0,219,0,0,0,0,0,201,0,0,0,180,0,183,0,132,0,0,0,75,0,0,0,63,0,123,0,0,0,92,0,0,0,11,0,0,0,41,0,157,0,90,0,185,0,219,0,145,0,164,0,6,0,0,0,186,0,48,0,0,0,0,0,236,0,46,0,0,0,0,0,78,0,0,0,233,0,35,0,206,0,27,0,80,0,99,0,139,0,150,0,41,0,137,0,53,0,0,0,51,0,0,0,237,0,0,0,245,0,0,0,203,0,96,0,248,0,154,0,100,0,155,0,0,0,24,0,254,0,154,0,0,0,0,0,254,0,231,0,152,0,152,0,201,0,191,0,86,0,112,0,238,0,0,0,135,0,83,0,161,0,183,0,0,0,0,0,27,0,0,0,0,0,110,0,0,0,58,0,72,0,127,0,132,0,175,0,0,0,52,0,167,0,0,0,154,0,91,0,0,0,0,0,0,0,191,0,0,0,186,0,16,0,208,0,120,0,179,0,5,0,0,0,191,0,173,0,0,0,125,0,228,0,247,0,83,0,99,0,151,0,135,0,86,0,139,0,0,0,0,0,20,0,80,0,0,0,96,0,215,0,162,0,129,0,137,0,183,0,0,0,0,0,92,0,91,0,1,0,5,0,0,0,101,0,0,0,0,0,0,0,150,0,67,0,64,0,0,0,73,0,0,0,0,0,99,0,57,0,38,0,152,0,199,0,162,0,208,0,67,0,29,0,0,0,85,0,0,0,132,0,212,0,0,0,6,0,133,0,153,0,67,0,4,0,39,0,175,0,142,0,134,0,0,0,237,0,148,0,26,0,47,0,193,0,121,0,153,0,0,0,23,0,211,0,103,0,204,0,221,0,0,0,237,0,219,0,0,0,0,0,0,0,224,0,0,0,96,0,52,0,244,0,0,0,96,0,0,0,86,0,217,0,126,0,0,0,56,0,19,0,209,0,220,0,0,0,23,0,86,0,0,0,98,0,173,0,76,0,0,0,54,0,0,0,156,0,0,0,180,0,0,0,36,0,119,0,15,0,127,0,31,0,191,0,0,0,206,0,194,0,216,0,76,0,0,0,45,0,0,0,115,0,12,0,54,0,155,0,133,0,34,0,147,0,63,0,248,0,66,0,119,0,242,0,249,0,89,0,0,0,51,0,167,0,18,0,117,0,9,0,23,0,22,0,38,0,33,0,238,0,195,0,5,0,162,0,238,0,184,0,0,0,2,0,252,0,0,0,0,0,0,0,27,0,0,0,28,0,158,0,116,0,170,0,32,0,43,0,168,0,190,0,187,0,0,0,0,0,0,0,47,0,221,0,94,0,221,0,109,0,10,0,189,0,204,0,247,0,53,0,0,0,0,0,22,0,25,0,123,0,205,0,97,0,225,0,167,0,95,0,207,0,128,0,35,0,178,0,103,0,246,0,0,0,61,0,0,0,183,0,33,0,136,0,159,0,138,0,176,0,221,0,187,0,106,0,51,0,231,0,144,0,169,0,0,0,13,0,82,0,0,0,117,0,206,0,106,0,241,0,71,0,121,0,34,0,26,0,21,0,26,0,0,0,56,0,118,0,158,0,139,0,61,0,0,0,74,0,108,0,0,0,98,0,232,0,228,0);
signal scenario_full  : scenario_type := (0,0,56,31,52,31,52,30,249,31,249,30,44,31,166,31,166,30,239,31,173,31,34,31,252,31,252,30,136,31,136,30,168,31,37,31,34,31,128,31,33,31,48,31,8,31,190,31,110,31,48,31,56,31,188,31,46,31,36,31,216,31,216,30,216,29,162,31,213,31,194,31,194,30,68,31,68,30,131,31,131,30,41,31,212,31,214,31,248,31,14,31,53,31,107,31,107,30,107,29,83,31,83,30,83,29,52,31,235,31,199,31,199,31,38,31,238,31,238,30,238,29,136,31,17,31,53,31,225,31,209,31,149,31,149,30,132,31,204,31,231,31,231,30,125,31,45,31,45,30,45,29,56,31,150,31,208,31,209,31,169,31,72,31,127,31,191,31,99,31,235,31,168,31,207,31,173,31,33,31,67,31,131,31,143,31,81,31,61,31,61,30,219,31,131,31,181,31,26,31,14,31,175,31,45,31,45,30,6,31,30,31,97,31,97,30,34,31,40,31,248,31,95,31,187,31,107,31,230,31,40,31,40,30,80,31,194,31,214,31,168,31,153,31,236,31,230,31,230,30,185,31,34,31,34,30,34,29,34,28,56,31,56,30,61,31,230,31,126,31,244,31,215,31,63,31,67,31,67,30,21,31,178,31,135,31,153,31,37,31,86,31,85,31,148,31,216,31,199,31,83,31,46,31,190,31,133,31,150,31,28,31,243,31,119,31,119,30,86,31,86,30,5,31,26,31,26,30,230,31,231,31,237,31,117,31,149,31,149,30,23,31,140,31,88,31,156,31,180,31,78,31,78,30,127,31,7,31,205,31,205,30,111,31,150,31,150,30,103,31,147,31,147,30,147,29,107,31,107,30,147,31,51,31,106,31,157,31,29,31,235,31,245,31,169,31,116,31,116,30,77,31,15,31,200,31,220,31,206,31,206,30,182,31,100,31,100,30,157,31,23,31,171,31,176,31,47,31,18,31,141,31,127,31,175,31,56,31,212,31,60,31,111,31,111,30,5,31,130,31,130,30,250,31,144,31,144,30,241,31,85,31,212,31,227,31,70,31,120,31,80,31,136,31,136,30,136,29,27,31,11,31,11,30,167,31,33,31,85,31,85,30,207,31,196,31,25,31,20,31,11,31,108,31,108,30,105,31,207,31,242,31,242,30,203,31,63,31,63,30,63,29,91,31,58,31,219,31,219,30,219,29,242,31,242,30,139,31,139,30,139,29,23,31,121,31,40,31,172,31,232,31,11,31,148,31,137,31,184,31,28,31,105,31,93,31,98,31,34,31,34,30,34,29,103,31,7,31,26,31,26,30,92,31,92,30,219,31,219,30,219,29,201,31,201,30,180,31,183,31,132,31,132,30,75,31,75,30,63,31,123,31,123,30,92,31,92,30,11,31,11,30,41,31,157,31,90,31,185,31,219,31,145,31,164,31,6,31,6,30,186,31,48,31,48,30,48,29,236,31,46,31,46,30,46,29,78,31,78,30,233,31,35,31,206,31,27,31,80,31,99,31,139,31,150,31,41,31,137,31,53,31,53,30,51,31,51,30,237,31,237,30,245,31,245,30,203,31,96,31,248,31,154,31,100,31,155,31,155,30,24,31,254,31,154,31,154,30,154,29,254,31,231,31,152,31,152,31,201,31,191,31,86,31,112,31,238,31,238,30,135,31,83,31,161,31,183,31,183,30,183,29,27,31,27,30,27,29,110,31,110,30,58,31,72,31,127,31,132,31,175,31,175,30,52,31,167,31,167,30,154,31,91,31,91,30,91,29,91,28,191,31,191,30,186,31,16,31,208,31,120,31,179,31,5,31,5,30,191,31,173,31,173,30,125,31,228,31,247,31,83,31,99,31,151,31,135,31,86,31,139,31,139,30,139,29,20,31,80,31,80,30,96,31,215,31,162,31,129,31,137,31,183,31,183,30,183,29,92,31,91,31,1,31,5,31,5,30,101,31,101,30,101,29,101,28,150,31,67,31,64,31,64,30,73,31,73,30,73,29,99,31,57,31,38,31,152,31,199,31,162,31,208,31,67,31,29,31,29,30,85,31,85,30,132,31,212,31,212,30,6,31,133,31,153,31,67,31,4,31,39,31,175,31,142,31,134,31,134,30,237,31,148,31,26,31,47,31,193,31,121,31,153,31,153,30,23,31,211,31,103,31,204,31,221,31,221,30,237,31,219,31,219,30,219,29,219,28,224,31,224,30,96,31,52,31,244,31,244,30,96,31,96,30,86,31,217,31,126,31,126,30,56,31,19,31,209,31,220,31,220,30,23,31,86,31,86,30,98,31,173,31,76,31,76,30,54,31,54,30,156,31,156,30,180,31,180,30,36,31,119,31,15,31,127,31,31,31,191,31,191,30,206,31,194,31,216,31,76,31,76,30,45,31,45,30,115,31,12,31,54,31,155,31,133,31,34,31,147,31,63,31,248,31,66,31,119,31,242,31,249,31,89,31,89,30,51,31,167,31,18,31,117,31,9,31,23,31,22,31,38,31,33,31,238,31,195,31,5,31,162,31,238,31,184,31,184,30,2,31,252,31,252,30,252,29,252,28,27,31,27,30,28,31,158,31,116,31,170,31,32,31,43,31,168,31,190,31,187,31,187,30,187,29,187,28,47,31,221,31,94,31,221,31,109,31,10,31,189,31,204,31,247,31,53,31,53,30,53,29,22,31,25,31,123,31,205,31,97,31,225,31,167,31,95,31,207,31,128,31,35,31,178,31,103,31,246,31,246,30,61,31,61,30,183,31,33,31,136,31,159,31,138,31,176,31,221,31,187,31,106,31,51,31,231,31,144,31,169,31,169,30,13,31,82,31,82,30,117,31,206,31,106,31,241,31,71,31,121,31,34,31,26,31,21,31,26,31,26,30,56,31,118,31,158,31,139,31,61,31,61,30,74,31,108,31,108,30,98,31,232,31,228,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
