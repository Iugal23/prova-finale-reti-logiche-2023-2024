-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 312;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (157,0,28,0,0,0,248,0,0,0,152,0,127,0,151,0,41,0,74,0,117,0,100,0,130,0,132,0,189,0,249,0,244,0,212,0,175,0,198,0,62,0,221,0,216,0,252,0,142,0,18,0,122,0,0,0,147,0,162,0,91,0,156,0,11,0,168,0,62,0,124,0,67,0,69,0,120,0,157,0,19,0,219,0,161,0,191,0,8,0,109,0,129,0,108,0,96,0,148,0,208,0,130,0,179,0,0,0,20,0,245,0,24,0,118,0,95,0,140,0,0,0,24,0,124,0,43,0,112,0,25,0,131,0,114,0,134,0,125,0,112,0,93,0,124,0,243,0,92,0,67,0,0,0,84,0,213,0,101,0,119,0,0,0,81,0,161,0,0,0,0,0,164,0,35,0,150,0,112,0,68,0,82,0,242,0,191,0,27,0,51,0,0,0,175,0,225,0,16,0,0,0,129,0,108,0,0,0,99,0,235,0,0,0,0,0,22,0,0,0,237,0,134,0,0,0,95,0,0,0,105,0,10,0,195,0,25,0,251,0,196,0,21,0,240,0,0,0,106,0,0,0,0,0,178,0,239,0,0,0,62,0,89,0,13,0,0,0,192,0,161,0,210,0,210,0,243,0,13,0,0,0,24,0,0,0,94,0,235,0,0,0,138,0,142,0,189,0,0,0,48,0,226,0,117,0,105,0,69,0,30,0,86,0,130,0,42,0,0,0,206,0,207,0,33,0,46,0,19,0,143,0,162,0,0,0,0,0,0,0,214,0,195,0,0,0,17,0,214,0,251,0,178,0,0,0,250,0,46,0,0,0,1,0,20,0,147,0,68,0,235,0,153,0,22,0,0,0,17,0,234,0,91,0,119,0,77,0,217,0,0,0,184,0,219,0,162,0,29,0,49,0,156,0,29,0,115,0,202,0,55,0,124,0,0,0,195,0,57,0,56,0,62,0,96,0,136,0,247,0,0,0,0,0,209,0,0,0,137,0,37,0,105,0,0,0,107,0,231,0,0,0,56,0,214,0,0,0,246,0,47,0,55,0,146,0,82,0,181,0,232,0,154,0,0,0,180,0,113,0,193,0,195,0,11,0,72,0,166,0,160,0,98,0,104,0,195,0,136,0,239,0,217,0,123,0,0,0,141,0,94,0,168,0,255,0,202,0,161,0,67,0,255,0,0,0,47,0,0,0,7,0,252,0,0,0,106,0,5,0,146,0,215,0,129,0,242,0,0,0,146,0,114,0,0,0,0,0,0,0,93,0,246,0,0,0,0,0,232,0,57,0,198,0,206,0,205,0,88,0,0,0,89,0,0,0,50,0,140,0,179,0,123,0,119,0,147,0,115,0,88,0,28,0,213,0,204,0,163,0,146,0,0,0,0,0,234,0,48,0,164,0,145,0);
signal scenario_full  : scenario_type := (157,31,28,31,28,30,248,31,248,30,152,31,127,31,151,31,41,31,74,31,117,31,100,31,130,31,132,31,189,31,249,31,244,31,212,31,175,31,198,31,62,31,221,31,216,31,252,31,142,31,18,31,122,31,122,30,147,31,162,31,91,31,156,31,11,31,168,31,62,31,124,31,67,31,69,31,120,31,157,31,19,31,219,31,161,31,191,31,8,31,109,31,129,31,108,31,96,31,148,31,208,31,130,31,179,31,179,30,20,31,245,31,24,31,118,31,95,31,140,31,140,30,24,31,124,31,43,31,112,31,25,31,131,31,114,31,134,31,125,31,112,31,93,31,124,31,243,31,92,31,67,31,67,30,84,31,213,31,101,31,119,31,119,30,81,31,161,31,161,30,161,29,164,31,35,31,150,31,112,31,68,31,82,31,242,31,191,31,27,31,51,31,51,30,175,31,225,31,16,31,16,30,129,31,108,31,108,30,99,31,235,31,235,30,235,29,22,31,22,30,237,31,134,31,134,30,95,31,95,30,105,31,10,31,195,31,25,31,251,31,196,31,21,31,240,31,240,30,106,31,106,30,106,29,178,31,239,31,239,30,62,31,89,31,13,31,13,30,192,31,161,31,210,31,210,31,243,31,13,31,13,30,24,31,24,30,94,31,235,31,235,30,138,31,142,31,189,31,189,30,48,31,226,31,117,31,105,31,69,31,30,31,86,31,130,31,42,31,42,30,206,31,207,31,33,31,46,31,19,31,143,31,162,31,162,30,162,29,162,28,214,31,195,31,195,30,17,31,214,31,251,31,178,31,178,30,250,31,46,31,46,30,1,31,20,31,147,31,68,31,235,31,153,31,22,31,22,30,17,31,234,31,91,31,119,31,77,31,217,31,217,30,184,31,219,31,162,31,29,31,49,31,156,31,29,31,115,31,202,31,55,31,124,31,124,30,195,31,57,31,56,31,62,31,96,31,136,31,247,31,247,30,247,29,209,31,209,30,137,31,37,31,105,31,105,30,107,31,231,31,231,30,56,31,214,31,214,30,246,31,47,31,55,31,146,31,82,31,181,31,232,31,154,31,154,30,180,31,113,31,193,31,195,31,11,31,72,31,166,31,160,31,98,31,104,31,195,31,136,31,239,31,217,31,123,31,123,30,141,31,94,31,168,31,255,31,202,31,161,31,67,31,255,31,255,30,47,31,47,30,7,31,252,31,252,30,106,31,5,31,146,31,215,31,129,31,242,31,242,30,146,31,114,31,114,30,114,29,114,28,93,31,246,31,246,30,246,29,232,31,57,31,198,31,206,31,205,31,88,31,88,30,89,31,89,30,50,31,140,31,179,31,123,31,119,31,147,31,115,31,88,31,28,31,213,31,204,31,163,31,146,31,146,30,146,29,234,31,48,31,164,31,145,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
