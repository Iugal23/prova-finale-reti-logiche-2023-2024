-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 755;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,239,0,0,0,207,0,231,0,35,0,165,0,105,0,49,0,92,0,141,0,251,0,121,0,58,0,7,0,133,0,164,0,213,0,0,0,112,0,243,0,45,0,163,0,211,0,174,0,66,0,173,0,229,0,37,0,232,0,25,0,240,0,71,0,31,0,66,0,127,0,151,0,220,0,180,0,186,0,75,0,217,0,0,0,21,0,0,0,116,0,184,0,135,0,100,0,228,0,104,0,0,0,45,0,68,0,32,0,215,0,118,0,65,0,192,0,162,0,0,0,138,0,82,0,0,0,0,0,127,0,101,0,0,0,152,0,0,0,3,0,234,0,244,0,16,0,134,0,57,0,126,0,57,0,226,0,140,0,203,0,30,0,124,0,0,0,213,0,249,0,0,0,140,0,82,0,249,0,134,0,14,0,51,0,180,0,239,0,155,0,64,0,0,0,233,0,171,0,29,0,183,0,113,0,0,0,83,0,182,0,150,0,122,0,68,0,42,0,1,0,170,0,216,0,245,0,0,0,186,0,110,0,124,0,0,0,99,0,1,0,219,0,234,0,0,0,160,0,225,0,0,0,0,0,0,0,4,0,63,0,150,0,85,0,44,0,127,0,228,0,135,0,102,0,90,0,57,0,117,0,26,0,110,0,0,0,187,0,167,0,0,0,244,0,54,0,243,0,0,0,172,0,199,0,191,0,96,0,91,0,53,0,23,0,42,0,136,0,0,0,0,0,92,0,83,0,248,0,73,0,185,0,1,0,76,0,218,0,241,0,154,0,0,0,147,0,167,0,31,0,0,0,95,0,83,0,30,0,154,0,128,0,0,0,183,0,242,0,32,0,114,0,3,0,63,0,236,0,224,0,0,0,247,0,0,0,41,0,196,0,58,0,167,0,158,0,0,0,169,0,23,0,206,0,194,0,54,0,128,0,7,0,0,0,47,0,50,0,125,0,73,0,0,0,0,0,0,0,188,0,0,0,0,0,170,0,216,0,148,0,69,0,0,0,234,0,91,0,232,0,124,0,0,0,54,0,4,0,0,0,125,0,148,0,222,0,51,0,247,0,74,0,245,0,198,0,82,0,168,0,135,0,179,0,0,0,201,0,83,0,70,0,0,0,0,0,39,0,152,0,0,0,86,0,0,0,87,0,215,0,18,0,4,0,1,0,219,0,246,0,164,0,106,0,137,0,165,0,254,0,0,0,243,0,253,0,22,0,0,0,0,0,0,0,233,0,140,0,0,0,0,0,15,0,41,0,62,0,0,0,200,0,91,0,27,0,0,0,143,0,38,0,188,0,128,0,131,0,48,0,234,0,0,0,228,0,16,0,173,0,58,0,0,0,71,0,186,0,162,0,128,0,179,0,255,0,78,0,161,0,30,0,32,0,97,0,130,0,185,0,191,0,189,0,6,0,229,0,157,0,202,0,41,0,148,0,118,0,103,0,73,0,126,0,0,0,213,0,0,0,194,0,223,0,0,0,238,0,0,0,210,0,66,0,208,0,103,0,137,0,169,0,67,0,0,0,72,0,0,0,240,0,167,0,0,0,137,0,0,0,0,0,8,0,35,0,124,0,74,0,0,0,54,0,73,0,10,0,25,0,254,0,44,0,253,0,160,0,0,0,161,0,164,0,116,0,88,0,125,0,0,0,172,0,247,0,81,0,4,0,0,0,57,0,0,0,220,0,102,0,123,0,56,0,145,0,100,0,0,0,103,0,160,0,169,0,0,0,90,0,147,0,143,0,0,0,89,0,57,0,137,0,109,0,211,0,0,0,251,0,129,0,79,0,118,0,97,0,192,0,0,0,171,0,92,0,94,0,125,0,0,0,91,0,22,0,222,0,86,0,37,0,0,0,167,0,176,0,45,0,0,0,128,0,0,0,245,0,124,0,3,0,246,0,0,0,88,0,40,0,0,0,189,0,63,0,0,0,220,0,44,0,90,0,49,0,0,0,0,0,180,0,103,0,118,0,0,0,107,0,68,0,27,0,190,0,0,0,0,0,205,0,96,0,0,0,53,0,244,0,24,0,129,0,0,0,59,0,0,0,111,0,226,0,33,0,0,0,217,0,77,0,152,0,92,0,210,0,223,0,0,0,234,0,35,0,26,0,0,0,149,0,131,0,61,0,78,0,0,0,24,0,0,0,16,0,196,0,0,0,40,0,0,0,0,0,206,0,0,0,76,0,187,0,172,0,165,0,251,0,182,0,0,0,25,0,181,0,119,0,235,0,52,0,255,0,18,0,95,0,180,0,128,0,115,0,126,0,243,0,67,0,0,0,84,0,183,0,0,0,124,0,212,0,86,0,46,0,0,0,243,0,0,0,0,0,67,0,168,0,0,0,16,0,0,0,231,0,254,0,62,0,0,0,43,0,64,0,221,0,0,0,0,0,52,0,68,0,10,0,116,0,131,0,126,0,141,0,21,0,83,0,74,0,233,0,47,0,154,0,0,0,0,0,0,0,154,0,217,0,65,0,183,0,104,0,10,0,0,0,156,0,0,0,197,0,157,0,0,0,49,0,0,0,180,0,0,0,1,0,0,0,0,0,9,0,34,0,26,0,118,0,64,0,40,0,39,0,168,0,0,0,91,0,244,0,241,0,45,0,172,0,168,0,76,0,0,0,212,0,167,0,82,0,191,0,0,0,182,0,87,0,205,0,235,0,147,0,128,0,0,0,250,0,106,0,120,0,158,0,79,0,0,0,0,0,159,0,183,0,0,0,102,0,230,0,22,0,118,0,0,0,30,0,0,0,0,0,237,0,90,0,23,0,95,0,0,0,0,0,0,0,0,0,140,0,48,0,217,0,0,0,0,0,112,0,95,0,117,0,195,0,0,0,0,0,15,0,133,0,158,0,247,0,91,0,10,0,0,0,77,0,106,0,222,0,0,0,225,0,0,0,128,0,132,0,31,0,0,0,219,0,160,0,0,0,162,0,255,0,151,0,90,0,227,0,77,0,81,0,0,0,237,0,185,0,7,0,151,0,101,0,6,0,107,0,117,0,186,0,25,0,0,0,121,0,152,0,61,0,179,0,236,0,0,0,113,0,223,0,209,0,214,0,25,0,54,0,176,0,20,0,0,0,218,0,169,0,0,0,187,0,96,0,205,0,0,0,219,0,52,0,27,0,243,0,186,0,0,0,73,0,124,0,6,0,225,0,0,0,8,0,151,0,223,0,11,0,0,0,0,0,0,0,0,0,224,0,214,0,32,0,100,0,0,0,213,0,0,0,178,0,204,0,235,0,235,0,33,0,171,0,243,0,59,0,168,0,26,0,224,0,0,0,239,0,112,0,77,0,230,0,66,0,88,0,105,0,0,0,131,0,116,0,231,0,0,0,219,0,213,0,227,0,128,0,1,0,208,0,91,0,125,0,153,0,164,0);
signal scenario_full  : scenario_type := (0,0,239,31,239,30,207,31,231,31,35,31,165,31,105,31,49,31,92,31,141,31,251,31,121,31,58,31,7,31,133,31,164,31,213,31,213,30,112,31,243,31,45,31,163,31,211,31,174,31,66,31,173,31,229,31,37,31,232,31,25,31,240,31,71,31,31,31,66,31,127,31,151,31,220,31,180,31,186,31,75,31,217,31,217,30,21,31,21,30,116,31,184,31,135,31,100,31,228,31,104,31,104,30,45,31,68,31,32,31,215,31,118,31,65,31,192,31,162,31,162,30,138,31,82,31,82,30,82,29,127,31,101,31,101,30,152,31,152,30,3,31,234,31,244,31,16,31,134,31,57,31,126,31,57,31,226,31,140,31,203,31,30,31,124,31,124,30,213,31,249,31,249,30,140,31,82,31,249,31,134,31,14,31,51,31,180,31,239,31,155,31,64,31,64,30,233,31,171,31,29,31,183,31,113,31,113,30,83,31,182,31,150,31,122,31,68,31,42,31,1,31,170,31,216,31,245,31,245,30,186,31,110,31,124,31,124,30,99,31,1,31,219,31,234,31,234,30,160,31,225,31,225,30,225,29,225,28,4,31,63,31,150,31,85,31,44,31,127,31,228,31,135,31,102,31,90,31,57,31,117,31,26,31,110,31,110,30,187,31,167,31,167,30,244,31,54,31,243,31,243,30,172,31,199,31,191,31,96,31,91,31,53,31,23,31,42,31,136,31,136,30,136,29,92,31,83,31,248,31,73,31,185,31,1,31,76,31,218,31,241,31,154,31,154,30,147,31,167,31,31,31,31,30,95,31,83,31,30,31,154,31,128,31,128,30,183,31,242,31,32,31,114,31,3,31,63,31,236,31,224,31,224,30,247,31,247,30,41,31,196,31,58,31,167,31,158,31,158,30,169,31,23,31,206,31,194,31,54,31,128,31,7,31,7,30,47,31,50,31,125,31,73,31,73,30,73,29,73,28,188,31,188,30,188,29,170,31,216,31,148,31,69,31,69,30,234,31,91,31,232,31,124,31,124,30,54,31,4,31,4,30,125,31,148,31,222,31,51,31,247,31,74,31,245,31,198,31,82,31,168,31,135,31,179,31,179,30,201,31,83,31,70,31,70,30,70,29,39,31,152,31,152,30,86,31,86,30,87,31,215,31,18,31,4,31,1,31,219,31,246,31,164,31,106,31,137,31,165,31,254,31,254,30,243,31,253,31,22,31,22,30,22,29,22,28,233,31,140,31,140,30,140,29,15,31,41,31,62,31,62,30,200,31,91,31,27,31,27,30,143,31,38,31,188,31,128,31,131,31,48,31,234,31,234,30,228,31,16,31,173,31,58,31,58,30,71,31,186,31,162,31,128,31,179,31,255,31,78,31,161,31,30,31,32,31,97,31,130,31,185,31,191,31,189,31,6,31,229,31,157,31,202,31,41,31,148,31,118,31,103,31,73,31,126,31,126,30,213,31,213,30,194,31,223,31,223,30,238,31,238,30,210,31,66,31,208,31,103,31,137,31,169,31,67,31,67,30,72,31,72,30,240,31,167,31,167,30,137,31,137,30,137,29,8,31,35,31,124,31,74,31,74,30,54,31,73,31,10,31,25,31,254,31,44,31,253,31,160,31,160,30,161,31,164,31,116,31,88,31,125,31,125,30,172,31,247,31,81,31,4,31,4,30,57,31,57,30,220,31,102,31,123,31,56,31,145,31,100,31,100,30,103,31,160,31,169,31,169,30,90,31,147,31,143,31,143,30,89,31,57,31,137,31,109,31,211,31,211,30,251,31,129,31,79,31,118,31,97,31,192,31,192,30,171,31,92,31,94,31,125,31,125,30,91,31,22,31,222,31,86,31,37,31,37,30,167,31,176,31,45,31,45,30,128,31,128,30,245,31,124,31,3,31,246,31,246,30,88,31,40,31,40,30,189,31,63,31,63,30,220,31,44,31,90,31,49,31,49,30,49,29,180,31,103,31,118,31,118,30,107,31,68,31,27,31,190,31,190,30,190,29,205,31,96,31,96,30,53,31,244,31,24,31,129,31,129,30,59,31,59,30,111,31,226,31,33,31,33,30,217,31,77,31,152,31,92,31,210,31,223,31,223,30,234,31,35,31,26,31,26,30,149,31,131,31,61,31,78,31,78,30,24,31,24,30,16,31,196,31,196,30,40,31,40,30,40,29,206,31,206,30,76,31,187,31,172,31,165,31,251,31,182,31,182,30,25,31,181,31,119,31,235,31,52,31,255,31,18,31,95,31,180,31,128,31,115,31,126,31,243,31,67,31,67,30,84,31,183,31,183,30,124,31,212,31,86,31,46,31,46,30,243,31,243,30,243,29,67,31,168,31,168,30,16,31,16,30,231,31,254,31,62,31,62,30,43,31,64,31,221,31,221,30,221,29,52,31,68,31,10,31,116,31,131,31,126,31,141,31,21,31,83,31,74,31,233,31,47,31,154,31,154,30,154,29,154,28,154,31,217,31,65,31,183,31,104,31,10,31,10,30,156,31,156,30,197,31,157,31,157,30,49,31,49,30,180,31,180,30,1,31,1,30,1,29,9,31,34,31,26,31,118,31,64,31,40,31,39,31,168,31,168,30,91,31,244,31,241,31,45,31,172,31,168,31,76,31,76,30,212,31,167,31,82,31,191,31,191,30,182,31,87,31,205,31,235,31,147,31,128,31,128,30,250,31,106,31,120,31,158,31,79,31,79,30,79,29,159,31,183,31,183,30,102,31,230,31,22,31,118,31,118,30,30,31,30,30,30,29,237,31,90,31,23,31,95,31,95,30,95,29,95,28,95,27,140,31,48,31,217,31,217,30,217,29,112,31,95,31,117,31,195,31,195,30,195,29,15,31,133,31,158,31,247,31,91,31,10,31,10,30,77,31,106,31,222,31,222,30,225,31,225,30,128,31,132,31,31,31,31,30,219,31,160,31,160,30,162,31,255,31,151,31,90,31,227,31,77,31,81,31,81,30,237,31,185,31,7,31,151,31,101,31,6,31,107,31,117,31,186,31,25,31,25,30,121,31,152,31,61,31,179,31,236,31,236,30,113,31,223,31,209,31,214,31,25,31,54,31,176,31,20,31,20,30,218,31,169,31,169,30,187,31,96,31,205,31,205,30,219,31,52,31,27,31,243,31,186,31,186,30,73,31,124,31,6,31,225,31,225,30,8,31,151,31,223,31,11,31,11,30,11,29,11,28,11,27,224,31,214,31,32,31,100,31,100,30,213,31,213,30,178,31,204,31,235,31,235,31,33,31,171,31,243,31,59,31,168,31,26,31,224,31,224,30,239,31,112,31,77,31,230,31,66,31,88,31,105,31,105,30,131,31,116,31,231,31,231,30,219,31,213,31,227,31,128,31,1,31,208,31,91,31,125,31,153,31,164,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
