-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 487;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (245,0,187,0,63,0,117,0,251,0,232,0,69,0,183,0,0,0,236,0,199,0,0,0,239,0,85,0,222,0,111,0,0,0,0,0,0,0,99,0,131,0,222,0,220,0,0,0,119,0,44,0,212,0,0,0,0,0,0,0,60,0,168,0,104,0,0,0,171,0,44,0,116,0,2,0,5,0,102,0,128,0,219,0,252,0,0,0,3,0,52,0,0,0,0,0,0,0,138,0,12,0,0,0,193,0,0,0,4,0,46,0,221,0,0,0,0,0,188,0,240,0,42,0,28,0,137,0,239,0,244,0,178,0,13,0,89,0,248,0,114,0,0,0,253,0,118,0,163,0,69,0,251,0,0,0,205,0,172,0,0,0,49,0,0,0,172,0,0,0,82,0,19,0,146,0,80,0,15,0,150,0,33,0,52,0,231,0,75,0,0,0,0,0,0,0,133,0,28,0,104,0,167,0,61,0,0,0,0,0,189,0,182,0,0,0,0,0,0,0,0,0,1,0,120,0,215,0,5,0,186,0,94,0,0,0,97,0,0,0,41,0,90,0,48,0,0,0,182,0,0,0,193,0,223,0,236,0,0,0,217,0,11,0,210,0,7,0,182,0,243,0,0,0,5,0,69,0,193,0,227,0,211,0,150,0,91,0,206,0,7,0,0,0,79,0,8,0,111,0,0,0,18,0,55,0,181,0,229,0,202,0,112,0,109,0,0,0,164,0,43,0,151,0,109,0,125,0,167,0,0,0,6,0,220,0,202,0,0,0,14,0,124,0,244,0,155,0,248,0,168,0,208,0,78,0,76,0,78,0,0,0,171,0,0,0,0,0,231,0,0,0,78,0,0,0,110,0,2,0,52,0,0,0,30,0,201,0,128,0,0,0,25,0,72,0,104,0,0,0,131,0,0,0,0,0,209,0,156,0,161,0,0,0,54,0,0,0,39,0,200,0,173,0,0,0,0,0,145,0,11,0,0,0,0,0,71,0,42,0,97,0,54,0,141,0,0,0,10,0,195,0,38,0,13,0,137,0,242,0,75,0,75,0,54,0,0,0,0,0,132,0,0,0,232,0,244,0,126,0,223,0,0,0,64,0,34,0,0,0,179,0,39,0,35,0,249,0,60,0,184,0,97,0,248,0,195,0,230,0,143,0,229,0,214,0,212,0,0,0,152,0,251,0,254,0,51,0,180,0,125,0,223,0,0,0,159,0,14,0,250,0,163,0,181,0,15,0,92,0,244,0,144,0,203,0,105,0,167,0,14,0,93,0,0,0,135,0,141,0,0,0,168,0,193,0,126,0,181,0,117,0,114,0,211,0,168,0,66,0,199,0,40,0,5,0,119,0,205,0,82,0,223,0,102,0,191,0,229,0,243,0,50,0,19,0,0,0,0,0,216,0,120,0,145,0,135,0,167,0,0,0,0,0,248,0,180,0,204,0,23,0,22,0,181,0,146,0,146,0,9,0,68,0,98,0,92,0,39,0,146,0,0,0,22,0,92,0,173,0,0,0,26,0,233,0,136,0,105,0,184,0,224,0,0,0,165,0,65,0,0,0,57,0,249,0,182,0,119,0,239,0,202,0,135,0,0,0,196,0,138,0,190,0,243,0,185,0,0,0,67,0,37,0,4,0,0,0,212,0,0,0,58,0,53,0,160,0,14,0,0,0,0,0,76,0,194,0,201,0,142,0,184,0,141,0,18,0,146,0,82,0,70,0,80,0,246,0,246,0,182,0,205,0,206,0,203,0,0,0,180,0,253,0,141,0,0,0,6,0,173,0,244,0,37,0,228,0,107,0,0,0,0,0,0,0,0,0,236,0,0,0,104,0,40,0,27,0,0,0,150,0,0,0,0,0,238,0,155,0,102,0,254,0,249,0,221,0,0,0,250,0,48,0,0,0,97,0,212,0,0,0,225,0,150,0,0,0,186,0,1,0,147,0,242,0,205,0,0,0,0,0,58,0,136,0,0,0,49,0,245,0,206,0,88,0,242,0,136,0,16,0,53,0,228,0,47,0,197,0,0,0,221,0,163,0,240,0,0,0,21,0,79,0,221,0,0,0,102,0,196,0,130,0,235,0,0,0,224,0,0,0,101,0,248,0,0,0,123,0,106,0,116,0,43,0,87,0,196,0,0,0,213,0,0,0,0,0,63,0,140,0,0,0,225,0,144,0,148,0,70,0,19,0);
signal scenario_full  : scenario_type := (245,31,187,31,63,31,117,31,251,31,232,31,69,31,183,31,183,30,236,31,199,31,199,30,239,31,85,31,222,31,111,31,111,30,111,29,111,28,99,31,131,31,222,31,220,31,220,30,119,31,44,31,212,31,212,30,212,29,212,28,60,31,168,31,104,31,104,30,171,31,44,31,116,31,2,31,5,31,102,31,128,31,219,31,252,31,252,30,3,31,52,31,52,30,52,29,52,28,138,31,12,31,12,30,193,31,193,30,4,31,46,31,221,31,221,30,221,29,188,31,240,31,42,31,28,31,137,31,239,31,244,31,178,31,13,31,89,31,248,31,114,31,114,30,253,31,118,31,163,31,69,31,251,31,251,30,205,31,172,31,172,30,49,31,49,30,172,31,172,30,82,31,19,31,146,31,80,31,15,31,150,31,33,31,52,31,231,31,75,31,75,30,75,29,75,28,133,31,28,31,104,31,167,31,61,31,61,30,61,29,189,31,182,31,182,30,182,29,182,28,182,27,1,31,120,31,215,31,5,31,186,31,94,31,94,30,97,31,97,30,41,31,90,31,48,31,48,30,182,31,182,30,193,31,223,31,236,31,236,30,217,31,11,31,210,31,7,31,182,31,243,31,243,30,5,31,69,31,193,31,227,31,211,31,150,31,91,31,206,31,7,31,7,30,79,31,8,31,111,31,111,30,18,31,55,31,181,31,229,31,202,31,112,31,109,31,109,30,164,31,43,31,151,31,109,31,125,31,167,31,167,30,6,31,220,31,202,31,202,30,14,31,124,31,244,31,155,31,248,31,168,31,208,31,78,31,76,31,78,31,78,30,171,31,171,30,171,29,231,31,231,30,78,31,78,30,110,31,2,31,52,31,52,30,30,31,201,31,128,31,128,30,25,31,72,31,104,31,104,30,131,31,131,30,131,29,209,31,156,31,161,31,161,30,54,31,54,30,39,31,200,31,173,31,173,30,173,29,145,31,11,31,11,30,11,29,71,31,42,31,97,31,54,31,141,31,141,30,10,31,195,31,38,31,13,31,137,31,242,31,75,31,75,31,54,31,54,30,54,29,132,31,132,30,232,31,244,31,126,31,223,31,223,30,64,31,34,31,34,30,179,31,39,31,35,31,249,31,60,31,184,31,97,31,248,31,195,31,230,31,143,31,229,31,214,31,212,31,212,30,152,31,251,31,254,31,51,31,180,31,125,31,223,31,223,30,159,31,14,31,250,31,163,31,181,31,15,31,92,31,244,31,144,31,203,31,105,31,167,31,14,31,93,31,93,30,135,31,141,31,141,30,168,31,193,31,126,31,181,31,117,31,114,31,211,31,168,31,66,31,199,31,40,31,5,31,119,31,205,31,82,31,223,31,102,31,191,31,229,31,243,31,50,31,19,31,19,30,19,29,216,31,120,31,145,31,135,31,167,31,167,30,167,29,248,31,180,31,204,31,23,31,22,31,181,31,146,31,146,31,9,31,68,31,98,31,92,31,39,31,146,31,146,30,22,31,92,31,173,31,173,30,26,31,233,31,136,31,105,31,184,31,224,31,224,30,165,31,65,31,65,30,57,31,249,31,182,31,119,31,239,31,202,31,135,31,135,30,196,31,138,31,190,31,243,31,185,31,185,30,67,31,37,31,4,31,4,30,212,31,212,30,58,31,53,31,160,31,14,31,14,30,14,29,76,31,194,31,201,31,142,31,184,31,141,31,18,31,146,31,82,31,70,31,80,31,246,31,246,31,182,31,205,31,206,31,203,31,203,30,180,31,253,31,141,31,141,30,6,31,173,31,244,31,37,31,228,31,107,31,107,30,107,29,107,28,107,27,236,31,236,30,104,31,40,31,27,31,27,30,150,31,150,30,150,29,238,31,155,31,102,31,254,31,249,31,221,31,221,30,250,31,48,31,48,30,97,31,212,31,212,30,225,31,150,31,150,30,186,31,1,31,147,31,242,31,205,31,205,30,205,29,58,31,136,31,136,30,49,31,245,31,206,31,88,31,242,31,136,31,16,31,53,31,228,31,47,31,197,31,197,30,221,31,163,31,240,31,240,30,21,31,79,31,221,31,221,30,102,31,196,31,130,31,235,31,235,30,224,31,224,30,101,31,248,31,248,30,123,31,106,31,116,31,43,31,87,31,196,31,196,30,213,31,213,30,213,29,63,31,140,31,140,30,225,31,144,31,148,31,70,31,19,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
