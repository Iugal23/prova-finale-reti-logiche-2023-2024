-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_683 is
end project_tb_683;

architecture project_tb_arch_683 of project_tb_683 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 252;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,108,0,96,0,0,0,0,0,127,0,175,0,165,0,213,0,34,0,0,0,87,0,0,0,0,0,213,0,203,0,122,0,0,0,0,0,181,0,14,0,39,0,225,0,220,0,186,0,190,0,189,0,199,0,75,0,28,0,99,0,110,0,212,0,142,0,173,0,3,0,149,0,124,0,30,0,220,0,0,0,190,0,0,0,241,0,100,0,77,0,0,0,173,0,186,0,0,0,224,0,72,0,27,0,3,0,179,0,198,0,23,0,75,0,77,0,75,0,0,0,103,0,189,0,241,0,21,0,56,0,249,0,216,0,147,0,51,0,157,0,241,0,250,0,45,0,133,0,2,0,106,0,41,0,164,0,2,0,12,0,77,0,246,0,36,0,0,0,8,0,167,0,132,0,91,0,245,0,127,0,199,0,0,0,81,0,213,0,0,0,6,0,186,0,128,0,145,0,75,0,201,0,29,0,95,0,123,0,87,0,105,0,152,0,0,0,0,0,213,0,192,0,192,0,0,0,237,0,182,0,174,0,186,0,0,0,73,0,253,0,0,0,66,0,173,0,0,0,143,0,0,0,251,0,168,0,87,0,190,0,129,0,160,0,207,0,0,0,215,0,159,0,0,0,0,0,59,0,32,0,0,0,0,0,221,0,0,0,0,0,125,0,106,0,0,0,180,0,38,0,0,0,113,0,53,0,132,0,231,0,173,0,92,0,161,0,117,0,0,0,0,0,109,0,0,0,109,0,54,0,172,0,147,0,0,0,100,0,243,0,154,0,153,0,155,0,204,0,143,0,39,0,0,0,0,0,165,0,112,0,170,0,48,0,75,0,108,0,94,0,0,0,196,0,119,0,187,0,79,0,179,0,163,0,127,0,0,0,2,0,134,0,166,0,171,0,188,0,0,0,93,0,101,0,161,0,0,0,158,0,51,0,185,0,127,0,0,0,203,0,247,0,215,0,101,0,172,0,18,0,170,0,36,0,21,0,135,0,239,0,229,0,52,0,125,0,0,0,0,0,246,0,41,0,184,0,58,0,0,0,188,0,135,0,234,0,45,0,18,0,36,0,150,0,0,0,52,0,183,0,0,0,0,0,33,0,0,0,250,0,0,0,161,0,23,0,242,0,158,0,56,0);
signal scenario_full  : scenario_type := (0,0,108,31,96,31,96,30,96,29,127,31,175,31,165,31,213,31,34,31,34,30,87,31,87,30,87,29,213,31,203,31,122,31,122,30,122,29,181,31,14,31,39,31,225,31,220,31,186,31,190,31,189,31,199,31,75,31,28,31,99,31,110,31,212,31,142,31,173,31,3,31,149,31,124,31,30,31,220,31,220,30,190,31,190,30,241,31,100,31,77,31,77,30,173,31,186,31,186,30,224,31,72,31,27,31,3,31,179,31,198,31,23,31,75,31,77,31,75,31,75,30,103,31,189,31,241,31,21,31,56,31,249,31,216,31,147,31,51,31,157,31,241,31,250,31,45,31,133,31,2,31,106,31,41,31,164,31,2,31,12,31,77,31,246,31,36,31,36,30,8,31,167,31,132,31,91,31,245,31,127,31,199,31,199,30,81,31,213,31,213,30,6,31,186,31,128,31,145,31,75,31,201,31,29,31,95,31,123,31,87,31,105,31,152,31,152,30,152,29,213,31,192,31,192,31,192,30,237,31,182,31,174,31,186,31,186,30,73,31,253,31,253,30,66,31,173,31,173,30,143,31,143,30,251,31,168,31,87,31,190,31,129,31,160,31,207,31,207,30,215,31,159,31,159,30,159,29,59,31,32,31,32,30,32,29,221,31,221,30,221,29,125,31,106,31,106,30,180,31,38,31,38,30,113,31,53,31,132,31,231,31,173,31,92,31,161,31,117,31,117,30,117,29,109,31,109,30,109,31,54,31,172,31,147,31,147,30,100,31,243,31,154,31,153,31,155,31,204,31,143,31,39,31,39,30,39,29,165,31,112,31,170,31,48,31,75,31,108,31,94,31,94,30,196,31,119,31,187,31,79,31,179,31,163,31,127,31,127,30,2,31,134,31,166,31,171,31,188,31,188,30,93,31,101,31,161,31,161,30,158,31,51,31,185,31,127,31,127,30,203,31,247,31,215,31,101,31,172,31,18,31,170,31,36,31,21,31,135,31,239,31,229,31,52,31,125,31,125,30,125,29,246,31,41,31,184,31,58,31,58,30,188,31,135,31,234,31,45,31,18,31,36,31,150,31,150,30,52,31,183,31,183,30,183,29,33,31,33,30,250,31,250,30,161,31,23,31,242,31,158,31,56,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
