-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_420 is
end project_tb_420;

architecture project_tb_arch_420 of project_tb_420 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 276;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (55,0,0,0,60,0,0,0,148,0,81,0,0,0,200,0,191,0,127,0,0,0,201,0,134,0,25,0,243,0,168,0,213,0,180,0,54,0,122,0,0,0,188,0,115,0,0,0,180,0,61,0,119,0,245,0,67,0,0,0,221,0,38,0,0,0,224,0,162,0,242,0,175,0,26,0,188,0,0,0,178,0,74,0,121,0,120,0,108,0,67,0,166,0,223,0,28,0,94,0,90,0,73,0,213,0,234,0,134,0,57,0,31,0,233,0,161,0,47,0,0,0,157,0,214,0,0,0,236,0,0,0,214,0,176,0,249,0,231,0,187,0,78,0,190,0,141,0,43,0,74,0,158,0,236,0,0,0,41,0,51,0,0,0,82,0,143,0,211,0,157,0,250,0,147,0,75,0,34,0,169,0,31,0,165,0,222,0,165,0,22,0,0,0,97,0,0,0,175,0,53,0,80,0,236,0,0,0,200,0,26,0,247,0,0,0,27,0,106,0,117,0,249,0,9,0,213,0,130,0,255,0,215,0,205,0,2,0,26,0,0,0,0,0,122,0,44,0,60,0,115,0,192,0,253,0,0,0,66,0,179,0,188,0,79,0,57,0,0,0,168,0,71,0,0,0,0,0,136,0,114,0,75,0,0,0,134,0,185,0,229,0,24,0,139,0,10,0,170,0,0,0,0,0,53,0,52,0,42,0,211,0,82,0,19,0,29,0,111,0,2,0,3,0,139,0,0,0,240,0,0,0,162,0,98,0,173,0,6,0,202,0,206,0,15,0,232,0,0,0,238,0,0,0,170,0,240,0,0,0,7,0,176,0,227,0,150,0,175,0,188,0,152,0,171,0,20,0,109,0,16,0,33,0,15,0,0,0,160,0,81,0,215,0,12,0,17,0,0,0,0,0,0,0,160,0,77,0,216,0,115,0,250,0,48,0,211,0,206,0,90,0,95,0,50,0,0,0,65,0,89,0,0,0,139,0,124,0,0,0,233,0,252,0,188,0,0,0,0,0,111,0,1,0,26,0,240,0,25,0,185,0,39,0,0,0,18,0,0,0,95,0,194,0,176,0,191,0,0,0,82,0,242,0,0,0,219,0,7,0,0,0,1,0,209,0,126,0,241,0,238,0,136,0,0,0,129,0,93,0,138,0,90,0,251,0,159,0,0,0,20,0,0,0,186,0,190,0,0,0,244,0,0,0,91,0,28,0,237,0,0,0,96,0,190,0,215,0,69,0,14,0);
signal scenario_full  : scenario_type := (55,31,55,30,60,31,60,30,148,31,81,31,81,30,200,31,191,31,127,31,127,30,201,31,134,31,25,31,243,31,168,31,213,31,180,31,54,31,122,31,122,30,188,31,115,31,115,30,180,31,61,31,119,31,245,31,67,31,67,30,221,31,38,31,38,30,224,31,162,31,242,31,175,31,26,31,188,31,188,30,178,31,74,31,121,31,120,31,108,31,67,31,166,31,223,31,28,31,94,31,90,31,73,31,213,31,234,31,134,31,57,31,31,31,233,31,161,31,47,31,47,30,157,31,214,31,214,30,236,31,236,30,214,31,176,31,249,31,231,31,187,31,78,31,190,31,141,31,43,31,74,31,158,31,236,31,236,30,41,31,51,31,51,30,82,31,143,31,211,31,157,31,250,31,147,31,75,31,34,31,169,31,31,31,165,31,222,31,165,31,22,31,22,30,97,31,97,30,175,31,53,31,80,31,236,31,236,30,200,31,26,31,247,31,247,30,27,31,106,31,117,31,249,31,9,31,213,31,130,31,255,31,215,31,205,31,2,31,26,31,26,30,26,29,122,31,44,31,60,31,115,31,192,31,253,31,253,30,66,31,179,31,188,31,79,31,57,31,57,30,168,31,71,31,71,30,71,29,136,31,114,31,75,31,75,30,134,31,185,31,229,31,24,31,139,31,10,31,170,31,170,30,170,29,53,31,52,31,42,31,211,31,82,31,19,31,29,31,111,31,2,31,3,31,139,31,139,30,240,31,240,30,162,31,98,31,173,31,6,31,202,31,206,31,15,31,232,31,232,30,238,31,238,30,170,31,240,31,240,30,7,31,176,31,227,31,150,31,175,31,188,31,152,31,171,31,20,31,109,31,16,31,33,31,15,31,15,30,160,31,81,31,215,31,12,31,17,31,17,30,17,29,17,28,160,31,77,31,216,31,115,31,250,31,48,31,211,31,206,31,90,31,95,31,50,31,50,30,65,31,89,31,89,30,139,31,124,31,124,30,233,31,252,31,188,31,188,30,188,29,111,31,1,31,26,31,240,31,25,31,185,31,39,31,39,30,18,31,18,30,95,31,194,31,176,31,191,31,191,30,82,31,242,31,242,30,219,31,7,31,7,30,1,31,209,31,126,31,241,31,238,31,136,31,136,30,129,31,93,31,138,31,90,31,251,31,159,31,159,30,20,31,20,30,186,31,190,31,190,30,244,31,244,30,91,31,28,31,237,31,237,30,96,31,190,31,215,31,69,31,14,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
