-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_473 is
end project_tb_473;

architecture project_tb_arch_473 of project_tb_473 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 673;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (6,0,102,0,153,0,0,0,185,0,177,0,100,0,174,0,201,0,115,0,145,0,168,0,0,0,65,0,160,0,0,0,0,0,57,0,85,0,8,0,0,0,242,0,55,0,159,0,67,0,230,0,160,0,20,0,87,0,94,0,14,0,53,0,59,0,65,0,241,0,99,0,205,0,198,0,0,0,142,0,22,0,235,0,92,0,254,0,26,0,223,0,95,0,167,0,132,0,145,0,98,0,121,0,195,0,240,0,213,0,0,0,46,0,124,0,144,0,12,0,0,0,246,0,64,0,172,0,176,0,135,0,222,0,146,0,35,0,140,0,150,0,209,0,189,0,162,0,127,0,96,0,121,0,163,0,85,0,0,0,172,0,140,0,169,0,0,0,0,0,50,0,101,0,134,0,0,0,141,0,182,0,215,0,242,0,35,0,240,0,0,0,152,0,83,0,0,0,25,0,78,0,144,0,170,0,0,0,148,0,12,0,176,0,57,0,66,0,0,0,203,0,16,0,191,0,53,0,0,0,127,0,188,0,0,0,18,0,89,0,109,0,0,0,0,0,20,0,199,0,40,0,98,0,10,0,205,0,0,0,250,0,156,0,105,0,0,0,154,0,232,0,0,0,241,0,3,0,97,0,84,0,175,0,139,0,123,0,24,0,91,0,198,0,133,0,94,0,199,0,66,0,115,0,0,0,0,0,0,0,0,0,84,0,20,0,222,0,0,0,7,0,0,0,58,0,40,0,122,0,164,0,177,0,239,0,96,0,0,0,57,0,38,0,248,0,94,0,100,0,228,0,44,0,0,0,0,0,69,0,19,0,113,0,55,0,0,0,132,0,146,0,163,0,41,0,61,0,49,0,28,0,147,0,80,0,104,0,80,0,18,0,29,0,154,0,85,0,171,0,24,0,215,0,232,0,185,0,0,0,55,0,193,0,35,0,60,0,232,0,86,0,10,0,225,0,155,0,211,0,0,0,114,0,102,0,0,0,0,0,183,0,0,0,0,0,228,0,0,0,0,0,15,0,105,0,155,0,183,0,0,0,128,0,56,0,0,0,149,0,0,0,200,0,242,0,0,0,149,0,2,0,160,0,96,0,223,0,82,0,0,0,169,0,0,0,179,0,238,0,40,0,58,0,0,0,119,0,147,0,0,0,254,0,98,0,183,0,0,0,253,0,0,0,151,0,93,0,207,0,79,0,79,0,110,0,92,0,8,0,238,0,240,0,106,0,109,0,25,0,0,0,122,0,232,0,0,0,0,0,0,0,247,0,95,0,62,0,49,0,227,0,222,0,15,0,158,0,0,0,85,0,131,0,223,0,0,0,108,0,34,0,0,0,0,0,47,0,50,0,131,0,216,0,224,0,0,0,15,0,101,0,0,0,0,0,79,0,130,0,0,0,0,0,149,0,0,0,71,0,22,0,219,0,0,0,0,0,157,0,0,0,200,0,237,0,0,0,81,0,0,0,0,0,0,0,123,0,114,0,31,0,72,0,233,0,131,0,0,0,205,0,0,0,0,0,94,0,157,0,0,0,189,0,206,0,234,0,66,0,0,0,80,0,36,0,222,0,192,0,16,0,0,0,58,0,58,0,123,0,178,0,32,0,0,0,49,0,0,0,189,0,224,0,16,0,200,0,0,0,245,0,125,0,149,0,0,0,237,0,0,0,81,0,128,0,160,0,0,0,0,0,55,0,146,0,0,0,11,0,209,0,76,0,90,0,96,0,136,0,248,0,0,0,136,0,159,0,176,0,194,0,112,0,179,0,114,0,200,0,0,0,255,0,154,0,232,0,9,0,5,0,0,0,117,0,0,0,0,0,181,0,2,0,117,0,0,0,0,0,30,0,142,0,148,0,21,0,46,0,254,0,101,0,0,0,84,0,222,0,98,0,47,0,136,0,2,0,0,0,165,0,0,0,0,0,196,0,0,0,62,0,191,0,22,0,162,0,108,0,223,0,80,0,89,0,0,0,89,0,147,0,35,0,157,0,19,0,0,0,191,0,113,0,0,0,0,0,165,0,0,0,193,0,64,0,110,0,246,0,105,0,188,0,255,0,53,0,181,0,92,0,10,0,251,0,221,0,251,0,0,0,216,0,0,0,201,0,123,0,235,0,91,0,191,0,217,0,61,0,135,0,0,0,72,0,222,0,161,0,0,0,22,0,42,0,149,0,136,0,210,0,69,0,221,0,62,0,253,0,67,0,42,0,106,0,251,0,79,0,5,0,110,0,72,0,0,0,0,0,130,0,0,0,48,0,246,0,46,0,107,0,252,0,152,0,77,0,177,0,165,0,233,0,115,0,178,0,252,0,188,0,152,0,243,0,34,0,188,0,191,0,65,0,81,0,120,0,63,0,64,0,6,0,151,0,189,0,0,0,71,0,0,0,241,0,243,0,6,0,172,0,0,0,0,0,118,0,131,0,182,0,118,0,124,0,183,0,69,0,0,0,76,0,85,0,66,0,215,0,206,0,164,0,0,0,205,0,0,0,94,0,174,0,126,0,3,0,91,0,214,0,0,0,164,0,2,0,33,0,87,0,210,0,0,0,80,0,215,0,0,0,152,0,24,0,0,0,74,0,132,0,0,0,55,0,115,0,22,0,134,0,74,0,0,0,211,0,138,0,227,0,122,0,69,0,102,0,225,0,219,0,9,0,189,0,236,0,15,0,105,0,65,0,183,0,80,0,112,0,127,0,16,0,0,0,15,0,41,0,220,0,0,0,65,0,211,0,137,0,210,0,120,0,0,0,168,0,208,0,129,0,19,0,151,0,0,0,25,0,218,0,3,0,201,0,0,0,106,0,179,0,105,0,34,0,47,0,0,0,0,0,0,0,33,0,4,0,17,0,161,0,0,0,212,0,148,0,118,0,239,0,0,0,64,0,0,0,0,0,218,0,132,0,214,0,211,0,35,0,198,0,86,0,105,0,41,0,83,0,12,0,146,0,0,0,225,0,166,0,211,0,0,0,249,0,237,0,151,0,164,0,230,0,65,0,200,0,161,0,0,0,179,0,148,0);
signal scenario_full  : scenario_type := (6,31,102,31,153,31,153,30,185,31,177,31,100,31,174,31,201,31,115,31,145,31,168,31,168,30,65,31,160,31,160,30,160,29,57,31,85,31,8,31,8,30,242,31,55,31,159,31,67,31,230,31,160,31,20,31,87,31,94,31,14,31,53,31,59,31,65,31,241,31,99,31,205,31,198,31,198,30,142,31,22,31,235,31,92,31,254,31,26,31,223,31,95,31,167,31,132,31,145,31,98,31,121,31,195,31,240,31,213,31,213,30,46,31,124,31,144,31,12,31,12,30,246,31,64,31,172,31,176,31,135,31,222,31,146,31,35,31,140,31,150,31,209,31,189,31,162,31,127,31,96,31,121,31,163,31,85,31,85,30,172,31,140,31,169,31,169,30,169,29,50,31,101,31,134,31,134,30,141,31,182,31,215,31,242,31,35,31,240,31,240,30,152,31,83,31,83,30,25,31,78,31,144,31,170,31,170,30,148,31,12,31,176,31,57,31,66,31,66,30,203,31,16,31,191,31,53,31,53,30,127,31,188,31,188,30,18,31,89,31,109,31,109,30,109,29,20,31,199,31,40,31,98,31,10,31,205,31,205,30,250,31,156,31,105,31,105,30,154,31,232,31,232,30,241,31,3,31,97,31,84,31,175,31,139,31,123,31,24,31,91,31,198,31,133,31,94,31,199,31,66,31,115,31,115,30,115,29,115,28,115,27,84,31,20,31,222,31,222,30,7,31,7,30,58,31,40,31,122,31,164,31,177,31,239,31,96,31,96,30,57,31,38,31,248,31,94,31,100,31,228,31,44,31,44,30,44,29,69,31,19,31,113,31,55,31,55,30,132,31,146,31,163,31,41,31,61,31,49,31,28,31,147,31,80,31,104,31,80,31,18,31,29,31,154,31,85,31,171,31,24,31,215,31,232,31,185,31,185,30,55,31,193,31,35,31,60,31,232,31,86,31,10,31,225,31,155,31,211,31,211,30,114,31,102,31,102,30,102,29,183,31,183,30,183,29,228,31,228,30,228,29,15,31,105,31,155,31,183,31,183,30,128,31,56,31,56,30,149,31,149,30,200,31,242,31,242,30,149,31,2,31,160,31,96,31,223,31,82,31,82,30,169,31,169,30,179,31,238,31,40,31,58,31,58,30,119,31,147,31,147,30,254,31,98,31,183,31,183,30,253,31,253,30,151,31,93,31,207,31,79,31,79,31,110,31,92,31,8,31,238,31,240,31,106,31,109,31,25,31,25,30,122,31,232,31,232,30,232,29,232,28,247,31,95,31,62,31,49,31,227,31,222,31,15,31,158,31,158,30,85,31,131,31,223,31,223,30,108,31,34,31,34,30,34,29,47,31,50,31,131,31,216,31,224,31,224,30,15,31,101,31,101,30,101,29,79,31,130,31,130,30,130,29,149,31,149,30,71,31,22,31,219,31,219,30,219,29,157,31,157,30,200,31,237,31,237,30,81,31,81,30,81,29,81,28,123,31,114,31,31,31,72,31,233,31,131,31,131,30,205,31,205,30,205,29,94,31,157,31,157,30,189,31,206,31,234,31,66,31,66,30,80,31,36,31,222,31,192,31,16,31,16,30,58,31,58,31,123,31,178,31,32,31,32,30,49,31,49,30,189,31,224,31,16,31,200,31,200,30,245,31,125,31,149,31,149,30,237,31,237,30,81,31,128,31,160,31,160,30,160,29,55,31,146,31,146,30,11,31,209,31,76,31,90,31,96,31,136,31,248,31,248,30,136,31,159,31,176,31,194,31,112,31,179,31,114,31,200,31,200,30,255,31,154,31,232,31,9,31,5,31,5,30,117,31,117,30,117,29,181,31,2,31,117,31,117,30,117,29,30,31,142,31,148,31,21,31,46,31,254,31,101,31,101,30,84,31,222,31,98,31,47,31,136,31,2,31,2,30,165,31,165,30,165,29,196,31,196,30,62,31,191,31,22,31,162,31,108,31,223,31,80,31,89,31,89,30,89,31,147,31,35,31,157,31,19,31,19,30,191,31,113,31,113,30,113,29,165,31,165,30,193,31,64,31,110,31,246,31,105,31,188,31,255,31,53,31,181,31,92,31,10,31,251,31,221,31,251,31,251,30,216,31,216,30,201,31,123,31,235,31,91,31,191,31,217,31,61,31,135,31,135,30,72,31,222,31,161,31,161,30,22,31,42,31,149,31,136,31,210,31,69,31,221,31,62,31,253,31,67,31,42,31,106,31,251,31,79,31,5,31,110,31,72,31,72,30,72,29,130,31,130,30,48,31,246,31,46,31,107,31,252,31,152,31,77,31,177,31,165,31,233,31,115,31,178,31,252,31,188,31,152,31,243,31,34,31,188,31,191,31,65,31,81,31,120,31,63,31,64,31,6,31,151,31,189,31,189,30,71,31,71,30,241,31,243,31,6,31,172,31,172,30,172,29,118,31,131,31,182,31,118,31,124,31,183,31,69,31,69,30,76,31,85,31,66,31,215,31,206,31,164,31,164,30,205,31,205,30,94,31,174,31,126,31,3,31,91,31,214,31,214,30,164,31,2,31,33,31,87,31,210,31,210,30,80,31,215,31,215,30,152,31,24,31,24,30,74,31,132,31,132,30,55,31,115,31,22,31,134,31,74,31,74,30,211,31,138,31,227,31,122,31,69,31,102,31,225,31,219,31,9,31,189,31,236,31,15,31,105,31,65,31,183,31,80,31,112,31,127,31,16,31,16,30,15,31,41,31,220,31,220,30,65,31,211,31,137,31,210,31,120,31,120,30,168,31,208,31,129,31,19,31,151,31,151,30,25,31,218,31,3,31,201,31,201,30,106,31,179,31,105,31,34,31,47,31,47,30,47,29,47,28,33,31,4,31,17,31,161,31,161,30,212,31,148,31,118,31,239,31,239,30,64,31,64,30,64,29,218,31,132,31,214,31,211,31,35,31,198,31,86,31,105,31,41,31,83,31,12,31,146,31,146,30,225,31,166,31,211,31,211,30,249,31,237,31,151,31,164,31,230,31,65,31,200,31,161,31,161,30,179,31,148,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
