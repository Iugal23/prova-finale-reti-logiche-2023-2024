-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_928 is
end project_tb_928;

architecture project_tb_arch_928 of project_tb_928 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 569;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (126,0,131,0,0,0,185,0,232,0,36,0,0,0,207,0,250,0,178,0,234,0,0,0,86,0,141,0,255,0,189,0,218,0,137,0,226,0,36,0,231,0,195,0,111,0,60,0,85,0,0,0,0,0,210,0,87,0,238,0,77,0,6,0,88,0,0,0,167,0,135,0,0,0,204,0,10,0,145,0,211,0,219,0,0,0,204,0,38,0,0,0,0,0,170,0,251,0,137,0,0,0,0,0,223,0,0,0,0,0,0,0,85,0,85,0,43,0,27,0,177,0,25,0,0,0,38,0,10,0,0,0,0,0,222,0,0,0,32,0,105,0,159,0,0,0,0,0,40,0,241,0,97,0,35,0,50,0,217,0,0,0,128,0,0,0,95,0,235,0,237,0,143,0,37,0,68,0,255,0,2,0,10,0,134,0,33,0,0,0,128,0,163,0,109,0,52,0,0,0,126,0,130,0,157,0,101,0,103,0,76,0,235,0,89,0,0,0,210,0,209,0,241,0,21,0,82,0,205,0,180,0,104,0,163,0,14,0,65,0,205,0,116,0,212,0,28,0,224,0,118,0,80,0,194,0,249,0,0,0,11,0,99,0,7,0,157,0,250,0,80,0,9,0,0,0,0,0,0,0,212,0,0,0,0,0,215,0,75,0,22,0,0,0,207,0,144,0,176,0,119,0,240,0,0,0,141,0,0,0,220,0,181,0,55,0,222,0,246,0,14,0,143,0,12,0,156,0,179,0,0,0,1,0,0,0,216,0,46,0,252,0,0,0,122,0,14,0,225,0,98,0,246,0,249,0,134,0,171,0,0,0,119,0,0,0,0,0,0,0,38,0,0,0,171,0,139,0,0,0,0,0,119,0,62,0,97,0,0,0,234,0,19,0,138,0,0,0,113,0,235,0,38,0,173,0,233,0,0,0,11,0,6,0,133,0,82,0,4,0,98,0,113,0,21,0,114,0,200,0,88,0,122,0,112,0,0,0,247,0,0,0,163,0,0,0,142,0,0,0,0,0,46,0,211,0,226,0,186,0,96,0,0,0,227,0,26,0,215,0,99,0,213,0,171,0,126,0,56,0,11,0,0,0,61,0,249,0,71,0,183,0,0,0,0,0,96,0,25,0,98,0,0,0,151,0,178,0,105,0,186,0,174,0,0,0,193,0,0,0,159,0,77,0,66,0,177,0,245,0,138,0,221,0,106,0,114,0,0,0,16,0,1,0,200,0,0,0,0,0,197,0,211,0,161,0,28,0,0,0,205,0,226,0,201,0,109,0,0,0,214,0,68,0,16,0,29,0,24,0,237,0,82,0,148,0,233,0,174,0,0,0,251,0,227,0,0,0,48,0,77,0,121,0,142,0,146,0,34,0,41,0,246,0,173,0,197,0,189,0,243,0,170,0,74,0,53,0,0,0,66,0,189,0,10,0,82,0,99,0,46,0,115,0,86,0,61,0,193,0,164,0,137,0,0,0,199,0,54,0,93,0,18,0,0,0,160,0,159,0,212,0,247,0,17,0,5,0,188,0,132,0,0,0,71,0,6,0,37,0,78,0,34,0,40,0,30,0,223,0,203,0,50,0,84,0,134,0,84,0,243,0,0,0,83,0,136,0,0,0,175,0,0,0,254,0,210,0,185,0,172,0,76,0,248,0,0,0,206,0,69,0,128,0,33,0,0,0,243,0,41,0,198,0,165,0,0,0,99,0,0,0,38,0,184,0,0,0,242,0,164,0,99,0,0,0,0,0,234,0,72,0,117,0,82,0,98,0,83,0,20,0,2,0,3,0,0,0,238,0,0,0,0,0,50,0,130,0,48,0,43,0,53,0,118,0,14,0,137,0,0,0,210,0,57,0,0,0,142,0,160,0,194,0,0,0,0,0,0,0,80,0,184,0,214,0,0,0,135,0,217,0,174,0,68,0,72,0,97,0,98,0,49,0,221,0,0,0,110,0,145,0,0,0,175,0,0,0,216,0,167,0,35,0,85,0,207,0,107,0,245,0,107,0,0,0,91,0,99,0,227,0,142,0,0,0,108,0,182,0,210,0,205,0,59,0,167,0,0,0,249,0,243,0,251,0,118,0,133,0,109,0,43,0,0,0,169,0,65,0,232,0,21,0,107,0,117,0,242,0,165,0,162,0,216,0,5,0,62,0,197,0,0,0,87,0,175,0,0,0,195,0,138,0,127,0,77,0,219,0,0,0,13,0,0,0,0,0,22,0,1,0,99,0,0,0,91,0,162,0,27,0,157,0,75,0,144,0,0,0,0,0,2,0,240,0,247,0,249,0,243,0,81,0,235,0,65,0,97,0,18,0,163,0,0,0,236,0,194,0,136,0,43,0,161,0,11,0,0,0,86,0,212,0,97,0,0,0,254,0,0,0,240,0,0,0,104,0,79,0,58,0,40,0,88,0,0,0,177,0,160,0,220,0,188,0,227,0,0,0,0,0,155,0,12,0,202,0,161,0,65,0,0,0,135,0,0,0,186,0,0,0,24,0,74,0,42,0,232,0,141,0,109,0,115,0,0,0,223,0,241,0,164,0,205,0,233,0);
signal scenario_full  : scenario_type := (126,31,131,31,131,30,185,31,232,31,36,31,36,30,207,31,250,31,178,31,234,31,234,30,86,31,141,31,255,31,189,31,218,31,137,31,226,31,36,31,231,31,195,31,111,31,60,31,85,31,85,30,85,29,210,31,87,31,238,31,77,31,6,31,88,31,88,30,167,31,135,31,135,30,204,31,10,31,145,31,211,31,219,31,219,30,204,31,38,31,38,30,38,29,170,31,251,31,137,31,137,30,137,29,223,31,223,30,223,29,223,28,85,31,85,31,43,31,27,31,177,31,25,31,25,30,38,31,10,31,10,30,10,29,222,31,222,30,32,31,105,31,159,31,159,30,159,29,40,31,241,31,97,31,35,31,50,31,217,31,217,30,128,31,128,30,95,31,235,31,237,31,143,31,37,31,68,31,255,31,2,31,10,31,134,31,33,31,33,30,128,31,163,31,109,31,52,31,52,30,126,31,130,31,157,31,101,31,103,31,76,31,235,31,89,31,89,30,210,31,209,31,241,31,21,31,82,31,205,31,180,31,104,31,163,31,14,31,65,31,205,31,116,31,212,31,28,31,224,31,118,31,80,31,194,31,249,31,249,30,11,31,99,31,7,31,157,31,250,31,80,31,9,31,9,30,9,29,9,28,212,31,212,30,212,29,215,31,75,31,22,31,22,30,207,31,144,31,176,31,119,31,240,31,240,30,141,31,141,30,220,31,181,31,55,31,222,31,246,31,14,31,143,31,12,31,156,31,179,31,179,30,1,31,1,30,216,31,46,31,252,31,252,30,122,31,14,31,225,31,98,31,246,31,249,31,134,31,171,31,171,30,119,31,119,30,119,29,119,28,38,31,38,30,171,31,139,31,139,30,139,29,119,31,62,31,97,31,97,30,234,31,19,31,138,31,138,30,113,31,235,31,38,31,173,31,233,31,233,30,11,31,6,31,133,31,82,31,4,31,98,31,113,31,21,31,114,31,200,31,88,31,122,31,112,31,112,30,247,31,247,30,163,31,163,30,142,31,142,30,142,29,46,31,211,31,226,31,186,31,96,31,96,30,227,31,26,31,215,31,99,31,213,31,171,31,126,31,56,31,11,31,11,30,61,31,249,31,71,31,183,31,183,30,183,29,96,31,25,31,98,31,98,30,151,31,178,31,105,31,186,31,174,31,174,30,193,31,193,30,159,31,77,31,66,31,177,31,245,31,138,31,221,31,106,31,114,31,114,30,16,31,1,31,200,31,200,30,200,29,197,31,211,31,161,31,28,31,28,30,205,31,226,31,201,31,109,31,109,30,214,31,68,31,16,31,29,31,24,31,237,31,82,31,148,31,233,31,174,31,174,30,251,31,227,31,227,30,48,31,77,31,121,31,142,31,146,31,34,31,41,31,246,31,173,31,197,31,189,31,243,31,170,31,74,31,53,31,53,30,66,31,189,31,10,31,82,31,99,31,46,31,115,31,86,31,61,31,193,31,164,31,137,31,137,30,199,31,54,31,93,31,18,31,18,30,160,31,159,31,212,31,247,31,17,31,5,31,188,31,132,31,132,30,71,31,6,31,37,31,78,31,34,31,40,31,30,31,223,31,203,31,50,31,84,31,134,31,84,31,243,31,243,30,83,31,136,31,136,30,175,31,175,30,254,31,210,31,185,31,172,31,76,31,248,31,248,30,206,31,69,31,128,31,33,31,33,30,243,31,41,31,198,31,165,31,165,30,99,31,99,30,38,31,184,31,184,30,242,31,164,31,99,31,99,30,99,29,234,31,72,31,117,31,82,31,98,31,83,31,20,31,2,31,3,31,3,30,238,31,238,30,238,29,50,31,130,31,48,31,43,31,53,31,118,31,14,31,137,31,137,30,210,31,57,31,57,30,142,31,160,31,194,31,194,30,194,29,194,28,80,31,184,31,214,31,214,30,135,31,217,31,174,31,68,31,72,31,97,31,98,31,49,31,221,31,221,30,110,31,145,31,145,30,175,31,175,30,216,31,167,31,35,31,85,31,207,31,107,31,245,31,107,31,107,30,91,31,99,31,227,31,142,31,142,30,108,31,182,31,210,31,205,31,59,31,167,31,167,30,249,31,243,31,251,31,118,31,133,31,109,31,43,31,43,30,169,31,65,31,232,31,21,31,107,31,117,31,242,31,165,31,162,31,216,31,5,31,62,31,197,31,197,30,87,31,175,31,175,30,195,31,138,31,127,31,77,31,219,31,219,30,13,31,13,30,13,29,22,31,1,31,99,31,99,30,91,31,162,31,27,31,157,31,75,31,144,31,144,30,144,29,2,31,240,31,247,31,249,31,243,31,81,31,235,31,65,31,97,31,18,31,163,31,163,30,236,31,194,31,136,31,43,31,161,31,11,31,11,30,86,31,212,31,97,31,97,30,254,31,254,30,240,31,240,30,104,31,79,31,58,31,40,31,88,31,88,30,177,31,160,31,220,31,188,31,227,31,227,30,227,29,155,31,12,31,202,31,161,31,65,31,65,30,135,31,135,30,186,31,186,30,24,31,74,31,42,31,232,31,141,31,109,31,115,31,115,30,223,31,241,31,164,31,205,31,233,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
