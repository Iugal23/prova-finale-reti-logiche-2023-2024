-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 790;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (95,0,47,0,179,0,28,0,100,0,40,0,249,0,137,0,108,0,119,0,90,0,0,0,34,0,2,0,28,0,120,0,1,0,0,0,16,0,218,0,106,0,214,0,102,0,160,0,91,0,163,0,206,0,61,0,159,0,214,0,75,0,207,0,245,0,152,0,246,0,141,0,182,0,174,0,143,0,209,0,59,0,0,0,55,0,0,0,102,0,0,0,213,0,23,0,207,0,63,0,58,0,182,0,27,0,252,0,137,0,50,0,21,0,109,0,0,0,211,0,0,0,204,0,238,0,15,0,234,0,0,0,57,0,13,0,23,0,37,0,5,0,0,0,0,0,242,0,103,0,143,0,201,0,82,0,156,0,0,0,98,0,89,0,45,0,200,0,21,0,113,0,145,0,215,0,171,0,89,0,184,0,0,0,140,0,222,0,0,0,86,0,184,0,150,0,52,0,9,0,216,0,116,0,221,0,147,0,145,0,59,0,217,0,187,0,137,0,195,0,0,0,89,0,107,0,0,0,196,0,212,0,76,0,0,0,0,0,168,0,78,0,140,0,141,0,221,0,0,0,244,0,80,0,185,0,138,0,85,0,0,0,15,0,16,0,0,0,209,0,0,0,0,0,161,0,0,0,32,0,193,0,145,0,0,0,17,0,6,0,0,0,126,0,0,0,80,0,0,0,173,0,0,0,48,0,0,0,66,0,254,0,215,0,139,0,113,0,243,0,150,0,0,0,213,0,35,0,24,0,0,0,205,0,0,0,90,0,60,0,162,0,221,0,113,0,55,0,0,0,128,0,98,0,208,0,177,0,133,0,129,0,238,0,54,0,145,0,102,0,12,0,133,0,222,0,94,0,204,0,136,0,234,0,9,0,202,0,16,0,105,0,254,0,0,0,116,0,74,0,100,0,57,0,48,0,24,0,204,0,247,0,47,0,86,0,217,0,2,0,183,0,241,0,0,0,157,0,165,0,86,0,0,0,128,0,241,0,228,0,0,0,33,0,28,0,1,0,81,0,125,0,68,0,0,0,117,0,137,0,0,0,3,0,157,0,84,0,182,0,75,0,0,0,0,0,124,0,0,0,104,0,43,0,0,0,245,0,32,0,119,0,0,0,173,0,231,0,104,0,160,0,166,0,129,0,127,0,35,0,183,0,89,0,27,0,66,0,50,0,136,0,4,0,29,0,131,0,124,0,192,0,168,0,87,0,97,0,49,0,253,0,0,0,0,0,0,0,105,0,110,0,80,0,170,0,6,0,115,0,0,0,132,0,133,0,241,0,218,0,121,0,135,0,174,0,0,0,0,0,132,0,41,0,98,0,250,0,144,0,252,0,124,0,0,0,234,0,34,0,197,0,0,0,180,0,178,0,127,0,0,0,36,0,0,0,118,0,193,0,65,0,228,0,122,0,0,0,255,0,0,0,92,0,103,0,195,0,250,0,89,0,221,0,235,0,0,0,0,0,97,0,214,0,205,0,244,0,61,0,0,0,0,0,127,0,0,0,142,0,107,0,0,0,0,0,69,0,114,0,215,0,88,0,78,0,23,0,178,0,62,0,70,0,199,0,245,0,82,0,40,0,117,0,0,0,127,0,36,0,147,0,38,0,106,0,0,0,171,0,173,0,28,0,188,0,15,0,56,0,150,0,129,0,0,0,0,0,212,0,221,0,0,0,92,0,66,0,31,0,0,0,162,0,186,0,168,0,0,0,177,0,249,0,46,0,215,0,0,0,115,0,236,0,12,0,197,0,12,0,240,0,139,0,106,0,248,0,79,0,47,0,15,0,51,0,0,0,227,0,237,0,136,0,249,0,203,0,64,0,235,0,222,0,0,0,227,0,88,0,0,0,0,0,14,0,116,0,0,0,232,0,0,0,3,0,208,0,85,0,166,0,0,0,102,0,241,0,124,0,103,0,22,0,1,0,58,0,154,0,9,0,0,0,246,0,39,0,187,0,94,0,0,0,115,0,121,0,158,0,0,0,0,0,139,0,65,0,168,0,0,0,146,0,0,0,155,0,23,0,63,0,15,0,46,0,16,0,148,0,129,0,161,0,81,0,188,0,0,0,14,0,201,0,84,0,79,0,179,0,61,0,135,0,0,0,233,0,51,0,74,0,251,0,228,0,137,0,0,0,0,0,222,0,236,0,17,0,0,0,241,0,0,0,237,0,141,0,233,0,82,0,202,0,76,0,62,0,29,0,182,0,245,0,154,0,77,0,37,0,30,0,2,0,0,0,0,0,63,0,190,0,74,0,134,0,97,0,22,0,19,0,206,0,37,0,172,0,136,0,12,0,0,0,0,0,80,0,0,0,193,0,212,0,127,0,239,0,98,0,144,0,0,0,0,0,79,0,211,0,0,0,141,0,0,0,230,0,31,0,171,0,113,0,247,0,86,0,0,0,7,0,190,0,0,0,95,0,248,0,173,0,120,0,73,0,0,0,242,0,149,0,213,0,0,0,140,0,21,0,197,0,195,0,0,0,31,0,185,0,49,0,12,0,87,0,166,0,225,0,209,0,193,0,210,0,0,0,95,0,191,0,0,0,0,0,184,0,216,0,5,0,168,0,208,0,206,0,45,0,76,0,164,0,89,0,0,0,44,0,0,0,0,0,77,0,50,0,0,0,83,0,22,0,83,0,1,0,68,0,220,0,75,0,100,0,180,0,245,0,0,0,0,0,0,0,133,0,219,0,230,0,219,0,184,0,240,0,245,0,0,0,0,0,194,0,46,0,117,0,35,0,160,0,225,0,1,0,49,0,243,0,172,0,31,0,186,0,0,0,24,0,135,0,11,0,198,0,0,0,40,0,103,0,102,0,25,0,128,0,12,0,0,0,103,0,67,0,177,0,231,0,238,0,94,0,222,0,71,0,169,0,173,0,245,0,0,0,185,0,243,0,39,0,32,0,88,0,153,0,151,0,0,0,84,0,244,0,43,0,0,0,212,0,218,0,30,0,132,0,0,0,233,0,115,0,121,0,106,0,228,0,43,0,0,0,220,0,94,0,211,0,0,0,13,0,221,0,243,0,34,0,0,0,227,0,130,0,82,0,35,0,15,0,236,0,151,0,69,0,166,0,172,0,28,0,0,0,173,0,151,0,113,0,205,0,9,0,243,0,222,0,29,0,97,0,20,0,173,0,49,0,236,0,0,0,9,0,232,0,130,0,14,0,180,0,0,0,131,0,0,0,8,0,180,0,211,0,6,0,78,0,8,0,251,0,60,0,201,0,0,0,64,0,4,0,0,0,82,0,0,0,0,0,190,0,24,0,189,0,0,0,178,0,122,0,105,0,112,0,0,0,111,0,247,0,0,0,0,0,46,0,93,0,0,0,198,0,172,0,228,0,115,0,153,0,156,0,191,0,220,0,85,0,194,0,77,0,80,0,110,0,20,0,96,0,158,0,199,0,170,0,25,0,231,0,77,0,3,0,89,0,250,0,130,0,189,0,56,0,211,0,107,0,0,0,14,0,106,0,61,0,63,0,88,0,77,0,247,0,1,0,208,0,0,0,183,0,214,0,199,0,191,0,0,0,170,0,223,0);
signal scenario_full  : scenario_type := (95,31,47,31,179,31,28,31,100,31,40,31,249,31,137,31,108,31,119,31,90,31,90,30,34,31,2,31,28,31,120,31,1,31,1,30,16,31,218,31,106,31,214,31,102,31,160,31,91,31,163,31,206,31,61,31,159,31,214,31,75,31,207,31,245,31,152,31,246,31,141,31,182,31,174,31,143,31,209,31,59,31,59,30,55,31,55,30,102,31,102,30,213,31,23,31,207,31,63,31,58,31,182,31,27,31,252,31,137,31,50,31,21,31,109,31,109,30,211,31,211,30,204,31,238,31,15,31,234,31,234,30,57,31,13,31,23,31,37,31,5,31,5,30,5,29,242,31,103,31,143,31,201,31,82,31,156,31,156,30,98,31,89,31,45,31,200,31,21,31,113,31,145,31,215,31,171,31,89,31,184,31,184,30,140,31,222,31,222,30,86,31,184,31,150,31,52,31,9,31,216,31,116,31,221,31,147,31,145,31,59,31,217,31,187,31,137,31,195,31,195,30,89,31,107,31,107,30,196,31,212,31,76,31,76,30,76,29,168,31,78,31,140,31,141,31,221,31,221,30,244,31,80,31,185,31,138,31,85,31,85,30,15,31,16,31,16,30,209,31,209,30,209,29,161,31,161,30,32,31,193,31,145,31,145,30,17,31,6,31,6,30,126,31,126,30,80,31,80,30,173,31,173,30,48,31,48,30,66,31,254,31,215,31,139,31,113,31,243,31,150,31,150,30,213,31,35,31,24,31,24,30,205,31,205,30,90,31,60,31,162,31,221,31,113,31,55,31,55,30,128,31,98,31,208,31,177,31,133,31,129,31,238,31,54,31,145,31,102,31,12,31,133,31,222,31,94,31,204,31,136,31,234,31,9,31,202,31,16,31,105,31,254,31,254,30,116,31,74,31,100,31,57,31,48,31,24,31,204,31,247,31,47,31,86,31,217,31,2,31,183,31,241,31,241,30,157,31,165,31,86,31,86,30,128,31,241,31,228,31,228,30,33,31,28,31,1,31,81,31,125,31,68,31,68,30,117,31,137,31,137,30,3,31,157,31,84,31,182,31,75,31,75,30,75,29,124,31,124,30,104,31,43,31,43,30,245,31,32,31,119,31,119,30,173,31,231,31,104,31,160,31,166,31,129,31,127,31,35,31,183,31,89,31,27,31,66,31,50,31,136,31,4,31,29,31,131,31,124,31,192,31,168,31,87,31,97,31,49,31,253,31,253,30,253,29,253,28,105,31,110,31,80,31,170,31,6,31,115,31,115,30,132,31,133,31,241,31,218,31,121,31,135,31,174,31,174,30,174,29,132,31,41,31,98,31,250,31,144,31,252,31,124,31,124,30,234,31,34,31,197,31,197,30,180,31,178,31,127,31,127,30,36,31,36,30,118,31,193,31,65,31,228,31,122,31,122,30,255,31,255,30,92,31,103,31,195,31,250,31,89,31,221,31,235,31,235,30,235,29,97,31,214,31,205,31,244,31,61,31,61,30,61,29,127,31,127,30,142,31,107,31,107,30,107,29,69,31,114,31,215,31,88,31,78,31,23,31,178,31,62,31,70,31,199,31,245,31,82,31,40,31,117,31,117,30,127,31,36,31,147,31,38,31,106,31,106,30,171,31,173,31,28,31,188,31,15,31,56,31,150,31,129,31,129,30,129,29,212,31,221,31,221,30,92,31,66,31,31,31,31,30,162,31,186,31,168,31,168,30,177,31,249,31,46,31,215,31,215,30,115,31,236,31,12,31,197,31,12,31,240,31,139,31,106,31,248,31,79,31,47,31,15,31,51,31,51,30,227,31,237,31,136,31,249,31,203,31,64,31,235,31,222,31,222,30,227,31,88,31,88,30,88,29,14,31,116,31,116,30,232,31,232,30,3,31,208,31,85,31,166,31,166,30,102,31,241,31,124,31,103,31,22,31,1,31,58,31,154,31,9,31,9,30,246,31,39,31,187,31,94,31,94,30,115,31,121,31,158,31,158,30,158,29,139,31,65,31,168,31,168,30,146,31,146,30,155,31,23,31,63,31,15,31,46,31,16,31,148,31,129,31,161,31,81,31,188,31,188,30,14,31,201,31,84,31,79,31,179,31,61,31,135,31,135,30,233,31,51,31,74,31,251,31,228,31,137,31,137,30,137,29,222,31,236,31,17,31,17,30,241,31,241,30,237,31,141,31,233,31,82,31,202,31,76,31,62,31,29,31,182,31,245,31,154,31,77,31,37,31,30,31,2,31,2,30,2,29,63,31,190,31,74,31,134,31,97,31,22,31,19,31,206,31,37,31,172,31,136,31,12,31,12,30,12,29,80,31,80,30,193,31,212,31,127,31,239,31,98,31,144,31,144,30,144,29,79,31,211,31,211,30,141,31,141,30,230,31,31,31,171,31,113,31,247,31,86,31,86,30,7,31,190,31,190,30,95,31,248,31,173,31,120,31,73,31,73,30,242,31,149,31,213,31,213,30,140,31,21,31,197,31,195,31,195,30,31,31,185,31,49,31,12,31,87,31,166,31,225,31,209,31,193,31,210,31,210,30,95,31,191,31,191,30,191,29,184,31,216,31,5,31,168,31,208,31,206,31,45,31,76,31,164,31,89,31,89,30,44,31,44,30,44,29,77,31,50,31,50,30,83,31,22,31,83,31,1,31,68,31,220,31,75,31,100,31,180,31,245,31,245,30,245,29,245,28,133,31,219,31,230,31,219,31,184,31,240,31,245,31,245,30,245,29,194,31,46,31,117,31,35,31,160,31,225,31,1,31,49,31,243,31,172,31,31,31,186,31,186,30,24,31,135,31,11,31,198,31,198,30,40,31,103,31,102,31,25,31,128,31,12,31,12,30,103,31,67,31,177,31,231,31,238,31,94,31,222,31,71,31,169,31,173,31,245,31,245,30,185,31,243,31,39,31,32,31,88,31,153,31,151,31,151,30,84,31,244,31,43,31,43,30,212,31,218,31,30,31,132,31,132,30,233,31,115,31,121,31,106,31,228,31,43,31,43,30,220,31,94,31,211,31,211,30,13,31,221,31,243,31,34,31,34,30,227,31,130,31,82,31,35,31,15,31,236,31,151,31,69,31,166,31,172,31,28,31,28,30,173,31,151,31,113,31,205,31,9,31,243,31,222,31,29,31,97,31,20,31,173,31,49,31,236,31,236,30,9,31,232,31,130,31,14,31,180,31,180,30,131,31,131,30,8,31,180,31,211,31,6,31,78,31,8,31,251,31,60,31,201,31,201,30,64,31,4,31,4,30,82,31,82,30,82,29,190,31,24,31,189,31,189,30,178,31,122,31,105,31,112,31,112,30,111,31,247,31,247,30,247,29,46,31,93,31,93,30,198,31,172,31,228,31,115,31,153,31,156,31,191,31,220,31,85,31,194,31,77,31,80,31,110,31,20,31,96,31,158,31,199,31,170,31,25,31,231,31,77,31,3,31,89,31,250,31,130,31,189,31,56,31,211,31,107,31,107,30,14,31,106,31,61,31,63,31,88,31,77,31,247,31,1,31,208,31,208,30,183,31,214,31,199,31,191,31,191,30,170,31,223,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
