-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 814;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,58,0,18,0,0,0,39,0,197,0,0,0,143,0,0,0,214,0,0,0,238,0,95,0,204,0,173,0,179,0,184,0,94,0,68,0,0,0,76,0,0,0,18,0,235,0,176,0,0,0,61,0,220,0,157,0,56,0,0,0,174,0,108,0,196,0,43,0,35,0,194,0,202,0,78,0,156,0,187,0,0,0,245,0,77,0,0,0,51,0,0,0,137,0,193,0,203,0,93,0,120,0,27,0,0,0,250,0,252,0,234,0,0,0,244,0,225,0,29,0,211,0,108,0,236,0,85,0,244,0,62,0,0,0,240,0,14,0,190,0,0,0,0,0,249,0,213,0,217,0,183,0,210,0,152,0,150,0,216,0,193,0,231,0,144,0,59,0,97,0,32,0,0,0,0,0,247,0,160,0,210,0,64,0,196,0,157,0,102,0,163,0,74,0,227,0,137,0,0,0,85,0,199,0,100,0,207,0,244,0,132,0,180,0,0,0,27,0,0,0,161,0,152,0,147,0,110,0,162,0,25,0,0,0,77,0,0,0,113,0,182,0,164,0,69,0,0,0,230,0,3,0,36,0,134,0,137,0,0,0,102,0,166,0,99,0,0,0,114,0,6,0,96,0,0,0,136,0,105,0,0,0,61,0,139,0,37,0,179,0,153,0,147,0,127,0,245,0,203,0,74,0,254,0,99,0,142,0,163,0,208,0,28,0,15,0,0,0,247,0,120,0,201,0,144,0,9,0,137,0,164,0,0,0,97,0,103,0,0,0,27,0,132,0,242,0,90,0,246,0,111,0,0,0,157,0,17,0,194,0,240,0,255,0,202,0,46,0,0,0,241,0,30,0,52,0,0,0,74,0,130,0,0,0,34,0,221,0,113,0,247,0,233,0,0,0,81,0,26,0,16,0,38,0,39,0,72,0,0,0,0,0,143,0,195,0,138,0,0,0,105,0,33,0,22,0,192,0,156,0,232,0,5,0,0,0,212,0,99,0,39,0,129,0,77,0,36,0,202,0,52,0,237,0,0,0,191,0,0,0,136,0,0,0,150,0,80,0,21,0,242,0,0,0,0,0,158,0,0,0,0,0,144,0,209,0,210,0,84,0,156,0,0,0,20,0,0,0,160,0,209,0,189,0,137,0,144,0,0,0,171,0,202,0,156,0,178,0,115,0,0,0,0,0,211,0,61,0,112,0,244,0,196,0,7,0,221,0,90,0,153,0,124,0,0,0,65,0,96,0,214,0,73,0,171,0,0,0,80,0,26,0,157,0,227,0,254,0,144,0,67,0,252,0,181,0,251,0,235,0,9,0,0,0,111,0,0,0,0,0,146,0,161,0,0,0,83,0,246,0,142,0,0,0,207,0,221,0,0,0,59,0,40,0,58,0,232,0,195,0,163,0,187,0,173,0,135,0,183,0,93,0,0,0,97,0,131,0,0,0,237,0,223,0,88,0,187,0,156,0,23,0,222,0,32,0,143,0,22,0,206,0,0,0,0,0,0,0,98,0,71,0,167,0,135,0,19,0,109,0,101,0,146,0,229,0,242,0,63,0,171,0,0,0,39,0,15,0,0,0,121,0,64,0,2,0,190,0,100,0,220,0,2,0,68,0,0,0,0,0,0,0,0,0,26,0,152,0,0,0,82,0,0,0,252,0,174,0,58,0,135,0,195,0,0,0,114,0,0,0,0,0,0,0,237,0,59,0,227,0,201,0,223,0,0,0,32,0,149,0,97,0,0,0,0,0,0,0,103,0,94,0,167,0,239,0,165,0,228,0,219,0,107,0,167,0,196,0,0,0,42,0,47,0,146,0,89,0,29,0,0,0,79,0,53,0,157,0,145,0,180,0,226,0,205,0,0,0,0,0,35,0,124,0,0,0,58,0,100,0,99,0,0,0,142,0,3,0,245,0,243,0,225,0,0,0,12,0,255,0,221,0,94,0,0,0,213,0,48,0,3,0,177,0,201,0,0,0,116,0,213,0,0,0,167,0,0,0,0,0,239,0,240,0,109,0,192,0,0,0,9,0,229,0,0,0,0,0,175,0,250,0,164,0,149,0,164,0,76,0,0,0,199,0,191,0,0,0,247,0,0,0,1,0,0,0,120,0,135,0,135,0,96,0,119,0,101,0,122,0,0,0,169,0,54,0,39,0,231,0,32,0,165,0,85,0,65,0,219,0,101,0,168,0,15,0,137,0,0,0,187,0,135,0,33,0,77,0,217,0,0,0,208,0,153,0,149,0,62,0,165,0,151,0,189,0,13,0,0,0,0,0,251,0,19,0,0,0,38,0,0,0,214,0,68,0,30,0,114,0,191,0,95,0,117,0,154,0,232,0,146,0,74,0,173,0,0,0,106,0,236,0,237,0,131,0,0,0,184,0,33,0,224,0,209,0,211,0,0,0,155,0,151,0,60,0,238,0,182,0,0,0,197,0,28,0,29,0,240,0,183,0,0,0,27,0,221,0,167,0,59,0,75,0,160,0,217,0,229,0,44,0,0,0,94,0,195,0,231,0,70,0,0,0,17,0,165,0,164,0,247,0,84,0,0,0,21,0,33,0,0,0,229,0,0,0,72,0,0,0,144,0,0,0,106,0,149,0,158,0,0,0,81,0,154,0,66,0,212,0,38,0,85,0,232,0,0,0,15,0,0,0,214,0,8,0,129,0,135,0,4,0,241,0,159,0,225,0,12,0,115,0,47,0,8,0,193,0,243,0,1,0,161,0,44,0,69,0,198,0,192,0,0,0,15,0,40,0,245,0,243,0,227,0,0,0,166,0,58,0,94,0,0,0,240,0,88,0,138,0,0,0,166,0,69,0,0,0,0,0,0,0,40,0,134,0,0,0,63,0,116,0,225,0,83,0,48,0,123,0,161,0,230,0,156,0,30,0,228,0,136,0,56,0,183,0,0,0,166,0,0,0,231,0,0,0,9,0,99,0,157,0,195,0,170,0,94,0,16,0,38,0,164,0,54,0,196,0,0,0,196,0,0,0,194,0,248,0,55,0,239,0,75,0,67,0,12,0,208,0,59,0,43,0,4,0,0,0,166,0,0,0,78,0,52,0,0,0,144,0,108,0,0,0,78,0,0,0,0,0,109,0,192,0,223,0,69,0,0,0,137,0,46,0,55,0,45,0,84,0,145,0,86,0,71,0,0,0,197,0,237,0,0,0,143,0,135,0,0,0,0,0,53,0,2,0,0,0,89,0,167,0,39,0,179,0,0,0,139,0,109,0,1,0,193,0,8,0,37,0,0,0,82,0,62,0,83,0,0,0,98,0,40,0,65,0,0,0,0,0,226,0,74,0,0,0,166,0,244,0,102,0,0,0,0,0,90,0,112,0,0,0,156,0,136,0,56,0,0,0,5,0,38,0,182,0,215,0,25,0,30,0,1,0,14,0,186,0,0,0,185,0,194,0,90,0,42,0,186,0,4,0,0,0,85,0,119,0,7,0,121,0,203,0,169,0,0,0,209,0,228,0,112,0,0,0,0,0,154,0,93,0,125,0,55,0,247,0,36,0,25,0,104,0,201,0,0,0,219,0,43,0,180,0,24,0,112,0,75,0,187,0,177,0,104,0,62,0,204,0,145,0,168,0,0,0,226,0,172,0,0,0,76,0,0,0,206,0,111,0,147,0,163,0,0,0);
signal scenario_full  : scenario_type := (0,0,58,31,18,31,18,30,39,31,197,31,197,30,143,31,143,30,214,31,214,30,238,31,95,31,204,31,173,31,179,31,184,31,94,31,68,31,68,30,76,31,76,30,18,31,235,31,176,31,176,30,61,31,220,31,157,31,56,31,56,30,174,31,108,31,196,31,43,31,35,31,194,31,202,31,78,31,156,31,187,31,187,30,245,31,77,31,77,30,51,31,51,30,137,31,193,31,203,31,93,31,120,31,27,31,27,30,250,31,252,31,234,31,234,30,244,31,225,31,29,31,211,31,108,31,236,31,85,31,244,31,62,31,62,30,240,31,14,31,190,31,190,30,190,29,249,31,213,31,217,31,183,31,210,31,152,31,150,31,216,31,193,31,231,31,144,31,59,31,97,31,32,31,32,30,32,29,247,31,160,31,210,31,64,31,196,31,157,31,102,31,163,31,74,31,227,31,137,31,137,30,85,31,199,31,100,31,207,31,244,31,132,31,180,31,180,30,27,31,27,30,161,31,152,31,147,31,110,31,162,31,25,31,25,30,77,31,77,30,113,31,182,31,164,31,69,31,69,30,230,31,3,31,36,31,134,31,137,31,137,30,102,31,166,31,99,31,99,30,114,31,6,31,96,31,96,30,136,31,105,31,105,30,61,31,139,31,37,31,179,31,153,31,147,31,127,31,245,31,203,31,74,31,254,31,99,31,142,31,163,31,208,31,28,31,15,31,15,30,247,31,120,31,201,31,144,31,9,31,137,31,164,31,164,30,97,31,103,31,103,30,27,31,132,31,242,31,90,31,246,31,111,31,111,30,157,31,17,31,194,31,240,31,255,31,202,31,46,31,46,30,241,31,30,31,52,31,52,30,74,31,130,31,130,30,34,31,221,31,113,31,247,31,233,31,233,30,81,31,26,31,16,31,38,31,39,31,72,31,72,30,72,29,143,31,195,31,138,31,138,30,105,31,33,31,22,31,192,31,156,31,232,31,5,31,5,30,212,31,99,31,39,31,129,31,77,31,36,31,202,31,52,31,237,31,237,30,191,31,191,30,136,31,136,30,150,31,80,31,21,31,242,31,242,30,242,29,158,31,158,30,158,29,144,31,209,31,210,31,84,31,156,31,156,30,20,31,20,30,160,31,209,31,189,31,137,31,144,31,144,30,171,31,202,31,156,31,178,31,115,31,115,30,115,29,211,31,61,31,112,31,244,31,196,31,7,31,221,31,90,31,153,31,124,31,124,30,65,31,96,31,214,31,73,31,171,31,171,30,80,31,26,31,157,31,227,31,254,31,144,31,67,31,252,31,181,31,251,31,235,31,9,31,9,30,111,31,111,30,111,29,146,31,161,31,161,30,83,31,246,31,142,31,142,30,207,31,221,31,221,30,59,31,40,31,58,31,232,31,195,31,163,31,187,31,173,31,135,31,183,31,93,31,93,30,97,31,131,31,131,30,237,31,223,31,88,31,187,31,156,31,23,31,222,31,32,31,143,31,22,31,206,31,206,30,206,29,206,28,98,31,71,31,167,31,135,31,19,31,109,31,101,31,146,31,229,31,242,31,63,31,171,31,171,30,39,31,15,31,15,30,121,31,64,31,2,31,190,31,100,31,220,31,2,31,68,31,68,30,68,29,68,28,68,27,26,31,152,31,152,30,82,31,82,30,252,31,174,31,58,31,135,31,195,31,195,30,114,31,114,30,114,29,114,28,237,31,59,31,227,31,201,31,223,31,223,30,32,31,149,31,97,31,97,30,97,29,97,28,103,31,94,31,167,31,239,31,165,31,228,31,219,31,107,31,167,31,196,31,196,30,42,31,47,31,146,31,89,31,29,31,29,30,79,31,53,31,157,31,145,31,180,31,226,31,205,31,205,30,205,29,35,31,124,31,124,30,58,31,100,31,99,31,99,30,142,31,3,31,245,31,243,31,225,31,225,30,12,31,255,31,221,31,94,31,94,30,213,31,48,31,3,31,177,31,201,31,201,30,116,31,213,31,213,30,167,31,167,30,167,29,239,31,240,31,109,31,192,31,192,30,9,31,229,31,229,30,229,29,175,31,250,31,164,31,149,31,164,31,76,31,76,30,199,31,191,31,191,30,247,31,247,30,1,31,1,30,120,31,135,31,135,31,96,31,119,31,101,31,122,31,122,30,169,31,54,31,39,31,231,31,32,31,165,31,85,31,65,31,219,31,101,31,168,31,15,31,137,31,137,30,187,31,135,31,33,31,77,31,217,31,217,30,208,31,153,31,149,31,62,31,165,31,151,31,189,31,13,31,13,30,13,29,251,31,19,31,19,30,38,31,38,30,214,31,68,31,30,31,114,31,191,31,95,31,117,31,154,31,232,31,146,31,74,31,173,31,173,30,106,31,236,31,237,31,131,31,131,30,184,31,33,31,224,31,209,31,211,31,211,30,155,31,151,31,60,31,238,31,182,31,182,30,197,31,28,31,29,31,240,31,183,31,183,30,27,31,221,31,167,31,59,31,75,31,160,31,217,31,229,31,44,31,44,30,94,31,195,31,231,31,70,31,70,30,17,31,165,31,164,31,247,31,84,31,84,30,21,31,33,31,33,30,229,31,229,30,72,31,72,30,144,31,144,30,106,31,149,31,158,31,158,30,81,31,154,31,66,31,212,31,38,31,85,31,232,31,232,30,15,31,15,30,214,31,8,31,129,31,135,31,4,31,241,31,159,31,225,31,12,31,115,31,47,31,8,31,193,31,243,31,1,31,161,31,44,31,69,31,198,31,192,31,192,30,15,31,40,31,245,31,243,31,227,31,227,30,166,31,58,31,94,31,94,30,240,31,88,31,138,31,138,30,166,31,69,31,69,30,69,29,69,28,40,31,134,31,134,30,63,31,116,31,225,31,83,31,48,31,123,31,161,31,230,31,156,31,30,31,228,31,136,31,56,31,183,31,183,30,166,31,166,30,231,31,231,30,9,31,99,31,157,31,195,31,170,31,94,31,16,31,38,31,164,31,54,31,196,31,196,30,196,31,196,30,194,31,248,31,55,31,239,31,75,31,67,31,12,31,208,31,59,31,43,31,4,31,4,30,166,31,166,30,78,31,52,31,52,30,144,31,108,31,108,30,78,31,78,30,78,29,109,31,192,31,223,31,69,31,69,30,137,31,46,31,55,31,45,31,84,31,145,31,86,31,71,31,71,30,197,31,237,31,237,30,143,31,135,31,135,30,135,29,53,31,2,31,2,30,89,31,167,31,39,31,179,31,179,30,139,31,109,31,1,31,193,31,8,31,37,31,37,30,82,31,62,31,83,31,83,30,98,31,40,31,65,31,65,30,65,29,226,31,74,31,74,30,166,31,244,31,102,31,102,30,102,29,90,31,112,31,112,30,156,31,136,31,56,31,56,30,5,31,38,31,182,31,215,31,25,31,30,31,1,31,14,31,186,31,186,30,185,31,194,31,90,31,42,31,186,31,4,31,4,30,85,31,119,31,7,31,121,31,203,31,169,31,169,30,209,31,228,31,112,31,112,30,112,29,154,31,93,31,125,31,55,31,247,31,36,31,25,31,104,31,201,31,201,30,219,31,43,31,180,31,24,31,112,31,75,31,187,31,177,31,104,31,62,31,204,31,145,31,168,31,168,30,226,31,172,31,172,30,76,31,76,30,206,31,111,31,147,31,163,31,163,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
