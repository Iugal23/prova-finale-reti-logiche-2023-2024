-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 310;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (47,0,168,0,189,0,10,0,218,0,18,0,0,0,156,0,148,0,174,0,0,0,0,0,0,0,63,0,0,0,14,0,59,0,0,0,154,0,0,0,98,0,0,0,112,0,101,0,124,0,39,0,0,0,41,0,104,0,119,0,248,0,169,0,0,0,0,0,0,0,10,0,31,0,109,0,207,0,101,0,108,0,142,0,73,0,45,0,213,0,54,0,31,0,63,0,202,0,106,0,234,0,217,0,109,0,0,0,198,0,219,0,192,0,122,0,0,0,0,0,84,0,125,0,79,0,159,0,254,0,61,0,164,0,227,0,0,0,83,0,144,0,14,0,92,0,100,0,190,0,14,0,0,0,98,0,0,0,0,0,68,0,148,0,108,0,0,0,16,0,140,0,72,0,0,0,235,0,194,0,81,0,177,0,29,0,95,0,0,0,0,0,198,0,96,0,247,0,158,0,99,0,112,0,170,0,117,0,173,0,181,0,234,0,111,0,36,0,5,0,27,0,0,0,188,0,12,0,29,0,107,0,0,0,198,0,203,0,66,0,122,0,243,0,94,0,103,0,226,0,60,0,84,0,77,0,23,0,0,0,150,0,0,0,69,0,129,0,25,0,215,0,164,0,85,0,141,0,250,0,73,0,0,0,178,0,22,0,184,0,134,0,53,0,215,0,98,0,156,0,254,0,244,0,0,0,0,0,163,0,0,0,0,0,220,0,202,0,64,0,2,0,33,0,90,0,187,0,66,0,66,0,29,0,0,0,0,0,12,0,108,0,0,0,223,0,0,0,39,0,244,0,131,0,11,0,85,0,0,0,0,0,105,0,18,0,228,0,245,0,0,0,122,0,188,0,145,0,8,0,111,0,17,0,0,0,211,0,0,0,0,0,104,0,9,0,113,0,92,0,162,0,151,0,227,0,0,0,248,0,212,0,133,0,83,0,0,0,0,0,127,0,220,0,0,0,120,0,0,0,25,0,139,0,40,0,147,0,46,0,139,0,225,0,148,0,0,0,86,0,61,0,9,0,0,0,78,0,75,0,112,0,0,0,177,0,0,0,97,0,0,0,230,0,208,0,62,0,60,0,236,0,211,0,114,0,184,0,11,0,118,0,196,0,154,0,238,0,0,0,224,0,138,0,74,0,0,0,45,0,0,0,194,0,96,0,0,0,233,0,195,0,146,0,68,0,186,0,144,0,137,0,0,0,254,0,230,0,197,0,140,0,212,0,218,0,72,0,0,0,31,0,171,0,157,0,121,0,26,0,201,0,86,0,0,0,100,0,0,0,160,0,70,0,61,0,0,0,112,0,52,0,216,0,0,0,97,0,0,0,0,0,123,0,21,0,81,0,0,0,189,0,0,0,0,0,0,0,0,0,134,0,103,0,204,0,0,0,0,0);
signal scenario_full  : scenario_type := (47,31,168,31,189,31,10,31,218,31,18,31,18,30,156,31,148,31,174,31,174,30,174,29,174,28,63,31,63,30,14,31,59,31,59,30,154,31,154,30,98,31,98,30,112,31,101,31,124,31,39,31,39,30,41,31,104,31,119,31,248,31,169,31,169,30,169,29,169,28,10,31,31,31,109,31,207,31,101,31,108,31,142,31,73,31,45,31,213,31,54,31,31,31,63,31,202,31,106,31,234,31,217,31,109,31,109,30,198,31,219,31,192,31,122,31,122,30,122,29,84,31,125,31,79,31,159,31,254,31,61,31,164,31,227,31,227,30,83,31,144,31,14,31,92,31,100,31,190,31,14,31,14,30,98,31,98,30,98,29,68,31,148,31,108,31,108,30,16,31,140,31,72,31,72,30,235,31,194,31,81,31,177,31,29,31,95,31,95,30,95,29,198,31,96,31,247,31,158,31,99,31,112,31,170,31,117,31,173,31,181,31,234,31,111,31,36,31,5,31,27,31,27,30,188,31,12,31,29,31,107,31,107,30,198,31,203,31,66,31,122,31,243,31,94,31,103,31,226,31,60,31,84,31,77,31,23,31,23,30,150,31,150,30,69,31,129,31,25,31,215,31,164,31,85,31,141,31,250,31,73,31,73,30,178,31,22,31,184,31,134,31,53,31,215,31,98,31,156,31,254,31,244,31,244,30,244,29,163,31,163,30,163,29,220,31,202,31,64,31,2,31,33,31,90,31,187,31,66,31,66,31,29,31,29,30,29,29,12,31,108,31,108,30,223,31,223,30,39,31,244,31,131,31,11,31,85,31,85,30,85,29,105,31,18,31,228,31,245,31,245,30,122,31,188,31,145,31,8,31,111,31,17,31,17,30,211,31,211,30,211,29,104,31,9,31,113,31,92,31,162,31,151,31,227,31,227,30,248,31,212,31,133,31,83,31,83,30,83,29,127,31,220,31,220,30,120,31,120,30,25,31,139,31,40,31,147,31,46,31,139,31,225,31,148,31,148,30,86,31,61,31,9,31,9,30,78,31,75,31,112,31,112,30,177,31,177,30,97,31,97,30,230,31,208,31,62,31,60,31,236,31,211,31,114,31,184,31,11,31,118,31,196,31,154,31,238,31,238,30,224,31,138,31,74,31,74,30,45,31,45,30,194,31,96,31,96,30,233,31,195,31,146,31,68,31,186,31,144,31,137,31,137,30,254,31,230,31,197,31,140,31,212,31,218,31,72,31,72,30,31,31,171,31,157,31,121,31,26,31,201,31,86,31,86,30,100,31,100,30,160,31,70,31,61,31,61,30,112,31,52,31,216,31,216,30,97,31,97,30,97,29,123,31,21,31,81,31,81,30,189,31,189,30,189,29,189,28,189,27,134,31,103,31,204,31,204,30,204,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
