-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_156 is
end project_tb_156;

architecture project_tb_arch_156 of project_tb_156 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 268;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (181,0,0,0,0,0,49,0,49,0,32,0,108,0,160,0,0,0,123,0,111,0,0,0,0,0,0,0,0,0,0,0,234,0,193,0,214,0,0,0,252,0,0,0,0,0,249,0,10,0,14,0,0,0,53,0,162,0,235,0,20,0,35,0,90,0,92,0,208,0,0,0,84,0,146,0,0,0,158,0,174,0,228,0,0,0,172,0,156,0,215,0,190,0,0,0,92,0,158,0,65,0,158,0,0,0,32,0,0,0,211,0,192,0,0,0,237,0,176,0,30,0,213,0,18,0,0,0,125,0,236,0,181,0,0,0,117,0,186,0,28,0,0,0,156,0,89,0,116,0,149,0,107,0,205,0,158,0,231,0,214,0,131,0,2,0,0,0,0,0,161,0,128,0,169,0,0,0,117,0,167,0,237,0,196,0,0,0,74,0,0,0,189,0,0,0,174,0,173,0,107,0,0,0,113,0,104,0,93,0,153,0,0,0,206,0,45,0,198,0,124,0,0,0,130,0,24,0,207,0,43,0,17,0,0,0,181,0,15,0,0,0,237,0,0,0,158,0,111,0,2,0,211,0,0,0,188,0,0,0,0,0,173,0,0,0,0,0,0,0,196,0,95,0,166,0,56,0,251,0,77,0,54,0,45,0,0,0,0,0,11,0,99,0,232,0,213,0,67,0,94,0,192,0,120,0,74,0,174,0,0,0,115,0,220,0,153,0,0,0,129,0,87,0,0,0,126,0,107,0,45,0,123,0,133,0,126,0,33,0,70,0,96,0,217,0,103,0,45,0,0,0,161,0,34,0,0,0,0,0,84,0,64,0,102,0,162,0,0,0,88,0,12,0,0,0,229,0,99,0,24,0,12,0,0,0,132,0,19,0,136,0,45,0,158,0,0,0,84,0,58,0,213,0,53,0,201,0,64,0,229,0,110,0,202,0,237,0,238,0,227,0,145,0,114,0,15,0,92,0,0,0,252,0,195,0,231,0,0,0,171,0,0,0,117,0,89,0,194,0,0,0,0,0,171,0,49,0,230,0,230,0,69,0,61,0,142,0,58,0,214,0,220,0,160,0,48,0,159,0,41,0,90,0,105,0,177,0,153,0,0,0,254,0,0,0,236,0,0,0,254,0,134,0,52,0,145,0,122,0,101,0,119,0,158,0,0,0,192,0,96,0,0,0,152,0,73,0,10,0,124,0,245,0,110,0);
signal scenario_full  : scenario_type := (181,31,181,30,181,29,49,31,49,31,32,31,108,31,160,31,160,30,123,31,111,31,111,30,111,29,111,28,111,27,111,26,234,31,193,31,214,31,214,30,252,31,252,30,252,29,249,31,10,31,14,31,14,30,53,31,162,31,235,31,20,31,35,31,90,31,92,31,208,31,208,30,84,31,146,31,146,30,158,31,174,31,228,31,228,30,172,31,156,31,215,31,190,31,190,30,92,31,158,31,65,31,158,31,158,30,32,31,32,30,211,31,192,31,192,30,237,31,176,31,30,31,213,31,18,31,18,30,125,31,236,31,181,31,181,30,117,31,186,31,28,31,28,30,156,31,89,31,116,31,149,31,107,31,205,31,158,31,231,31,214,31,131,31,2,31,2,30,2,29,161,31,128,31,169,31,169,30,117,31,167,31,237,31,196,31,196,30,74,31,74,30,189,31,189,30,174,31,173,31,107,31,107,30,113,31,104,31,93,31,153,31,153,30,206,31,45,31,198,31,124,31,124,30,130,31,24,31,207,31,43,31,17,31,17,30,181,31,15,31,15,30,237,31,237,30,158,31,111,31,2,31,211,31,211,30,188,31,188,30,188,29,173,31,173,30,173,29,173,28,196,31,95,31,166,31,56,31,251,31,77,31,54,31,45,31,45,30,45,29,11,31,99,31,232,31,213,31,67,31,94,31,192,31,120,31,74,31,174,31,174,30,115,31,220,31,153,31,153,30,129,31,87,31,87,30,126,31,107,31,45,31,123,31,133,31,126,31,33,31,70,31,96,31,217,31,103,31,45,31,45,30,161,31,34,31,34,30,34,29,84,31,64,31,102,31,162,31,162,30,88,31,12,31,12,30,229,31,99,31,24,31,12,31,12,30,132,31,19,31,136,31,45,31,158,31,158,30,84,31,58,31,213,31,53,31,201,31,64,31,229,31,110,31,202,31,237,31,238,31,227,31,145,31,114,31,15,31,92,31,92,30,252,31,195,31,231,31,231,30,171,31,171,30,117,31,89,31,194,31,194,30,194,29,171,31,49,31,230,31,230,31,69,31,61,31,142,31,58,31,214,31,220,31,160,31,48,31,159,31,41,31,90,31,105,31,177,31,153,31,153,30,254,31,254,30,236,31,236,30,254,31,134,31,52,31,145,31,122,31,101,31,119,31,158,31,158,30,192,31,96,31,96,30,152,31,73,31,10,31,124,31,245,31,110,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
