-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 188;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (145,0,93,0,0,0,4,0,73,0,98,0,176,0,0,0,0,0,58,0,0,0,60,0,97,0,159,0,0,0,36,0,0,0,232,0,206,0,115,0,62,0,32,0,246,0,95,0,113,0,12,0,0,0,76,0,98,0,0,0,4,0,110,0,0,0,102,0,0,0,173,0,137,0,125,0,179,0,191,0,91,0,197,0,51,0,9,0,169,0,132,0,114,0,0,0,222,0,229,0,68,0,169,0,224,0,0,0,228,0,45,0,210,0,0,0,30,0,76,0,0,0,252,0,246,0,97,0,0,0,8,0,28,0,112,0,138,0,0,0,90,0,0,0,29,0,71,0,0,0,0,0,237,0,154,0,224,0,98,0,227,0,0,0,158,0,107,0,68,0,0,0,0,0,229,0,216,0,238,0,0,0,72,0,198,0,0,0,0,0,177,0,203,0,0,0,154,0,156,0,11,0,99,0,28,0,17,0,53,0,255,0,179,0,138,0,203,0,39,0,0,0,53,0,51,0,0,0,179,0,17,0,106,0,124,0,129,0,183,0,105,0,31,0,77,0,144,0,0,0,20,0,151,0,61,0,82,0,6,0,159,0,24,0,212,0,102,0,16,0,176,0,11,0,156,0,0,0,193,0,255,0,0,0,232,0,0,0,211,0,99,0,125,0,137,0,0,0,60,0,206,0,236,0,132,0,85,0,59,0,124,0,0,0,131,0,24,0,235,0,0,0,42,0,130,0,126,0,253,0,28,0,226,0,210,0,213,0,152,0,12,0,184,0,208,0,212,0,0,0,0,0,174,0,99,0,65,0,0,0,92,0,72,0,255,0,199,0,30,0,0,0,0,0,156,0);
signal scenario_full  : scenario_type := (145,31,93,31,93,30,4,31,73,31,98,31,176,31,176,30,176,29,58,31,58,30,60,31,97,31,159,31,159,30,36,31,36,30,232,31,206,31,115,31,62,31,32,31,246,31,95,31,113,31,12,31,12,30,76,31,98,31,98,30,4,31,110,31,110,30,102,31,102,30,173,31,137,31,125,31,179,31,191,31,91,31,197,31,51,31,9,31,169,31,132,31,114,31,114,30,222,31,229,31,68,31,169,31,224,31,224,30,228,31,45,31,210,31,210,30,30,31,76,31,76,30,252,31,246,31,97,31,97,30,8,31,28,31,112,31,138,31,138,30,90,31,90,30,29,31,71,31,71,30,71,29,237,31,154,31,224,31,98,31,227,31,227,30,158,31,107,31,68,31,68,30,68,29,229,31,216,31,238,31,238,30,72,31,198,31,198,30,198,29,177,31,203,31,203,30,154,31,156,31,11,31,99,31,28,31,17,31,53,31,255,31,179,31,138,31,203,31,39,31,39,30,53,31,51,31,51,30,179,31,17,31,106,31,124,31,129,31,183,31,105,31,31,31,77,31,144,31,144,30,20,31,151,31,61,31,82,31,6,31,159,31,24,31,212,31,102,31,16,31,176,31,11,31,156,31,156,30,193,31,255,31,255,30,232,31,232,30,211,31,99,31,125,31,137,31,137,30,60,31,206,31,236,31,132,31,85,31,59,31,124,31,124,30,131,31,24,31,235,31,235,30,42,31,130,31,126,31,253,31,28,31,226,31,210,31,213,31,152,31,12,31,184,31,208,31,212,31,212,30,212,29,174,31,99,31,65,31,65,30,92,31,72,31,255,31,199,31,30,31,30,30,30,29,156,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
