-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 394;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (75,0,226,0,73,0,227,0,100,0,46,0,0,0,226,0,175,0,150,0,198,0,7,0,0,0,1,0,0,0,49,0,14,0,200,0,242,0,0,0,252,0,0,0,33,0,250,0,212,0,0,0,94,0,155,0,0,0,63,0,246,0,209,0,65,0,133,0,0,0,148,0,0,0,38,0,0,0,226,0,62,0,195,0,237,0,0,0,48,0,39,0,0,0,34,0,127,0,153,0,0,0,105,0,53,0,101,0,0,0,182,0,130,0,119,0,0,0,123,0,17,0,242,0,0,0,40,0,20,0,0,0,137,0,65,0,115,0,210,0,80,0,0,0,255,0,232,0,6,0,29,0,0,0,180,0,55,0,251,0,0,0,225,0,0,0,0,0,149,0,0,0,19,0,96,0,0,0,192,0,21,0,115,0,0,0,86,0,7,0,0,0,25,0,36,0,239,0,164,0,191,0,180,0,216,0,0,0,83,0,159,0,9,0,0,0,82,0,206,0,0,0,67,0,60,0,203,0,88,0,51,0,229,0,220,0,63,0,0,0,0,0,152,0,43,0,198,0,41,0,59,0,76,0,0,0,32,0,244,0,94,0,203,0,83,0,17,0,0,0,23,0,81,0,227,0,0,0,242,0,58,0,124,0,251,0,87,0,0,0,215,0,250,0,240,0,0,0,0,0,95,0,16,0,0,0,195,0,162,0,75,0,136,0,0,0,0,0,77,0,0,0,186,0,204,0,0,0,69,0,0,0,130,0,112,0,18,0,24,0,0,0,0,0,45,0,104,0,127,0,192,0,0,0,55,0,58,0,136,0,179,0,0,0,225,0,0,0,99,0,48,0,160,0,41,0,121,0,0,0,183,0,27,0,0,0,151,0,89,0,86,0,136,0,178,0,139,0,204,0,240,0,37,0,216,0,0,0,70,0,0,0,169,0,0,0,145,0,126,0,115,0,164,0,64,0,0,0,58,0,198,0,237,0,47,0,138,0,155,0,30,0,220,0,153,0,196,0,95,0,124,0,125,0,54,0,158,0,89,0,236,0,217,0,225,0,0,0,0,0,87,0,237,0,0,0,177,0,0,0,157,0,156,0,207,0,0,0,177,0,213,0,123,0,0,0,216,0,183,0,0,0,41,0,8,0,0,0,103,0,88,0,61,0,27,0,222,0,64,0,250,0,3,0,28,0,43,0,238,0,137,0,208,0,26,0,189,0,243,0,51,0,0,0,0,0,8,0,0,0,0,0,24,0,29,0,0,0,8,0,240,0,134,0,147,0,230,0,28,0,0,0,103,0,214,0,8,0,158,0,0,0,192,0,186,0,13,0,122,0,55,0,214,0,51,0,239,0,177,0,0,0,0,0,112,0,63,0,162,0,126,0,32,0,144,0,237,0,0,0,200,0,224,0,71,0,132,0,242,0,117,0,82,0,0,0,226,0,190,0,113,0,202,0,96,0,32,0,145,0,0,0,0,0,17,0,0,0,173,0,45,0,213,0,161,0,144,0,55,0,0,0,202,0,50,0,117,0,22,0,126,0,0,0,169,0,92,0,0,0,0,0,47,0,8,0,0,0,217,0,181,0,0,0,29,0,198,0,211,0,0,0,218,0,0,0,144,0,220,0,255,0,0,0,19,0,199,0,117,0,14,0,72,0,16,0,40,0,223,0,122,0,154,0,172,0,109,0,159,0,0,0,114,0,18,0,0,0,122,0,177,0,95,0,179,0,0,0,65,0,224,0,118,0,67,0,10,0,116,0,75,0,252,0,98,0,24,0);
signal scenario_full  : scenario_type := (75,31,226,31,73,31,227,31,100,31,46,31,46,30,226,31,175,31,150,31,198,31,7,31,7,30,1,31,1,30,49,31,14,31,200,31,242,31,242,30,252,31,252,30,33,31,250,31,212,31,212,30,94,31,155,31,155,30,63,31,246,31,209,31,65,31,133,31,133,30,148,31,148,30,38,31,38,30,226,31,62,31,195,31,237,31,237,30,48,31,39,31,39,30,34,31,127,31,153,31,153,30,105,31,53,31,101,31,101,30,182,31,130,31,119,31,119,30,123,31,17,31,242,31,242,30,40,31,20,31,20,30,137,31,65,31,115,31,210,31,80,31,80,30,255,31,232,31,6,31,29,31,29,30,180,31,55,31,251,31,251,30,225,31,225,30,225,29,149,31,149,30,19,31,96,31,96,30,192,31,21,31,115,31,115,30,86,31,7,31,7,30,25,31,36,31,239,31,164,31,191,31,180,31,216,31,216,30,83,31,159,31,9,31,9,30,82,31,206,31,206,30,67,31,60,31,203,31,88,31,51,31,229,31,220,31,63,31,63,30,63,29,152,31,43,31,198,31,41,31,59,31,76,31,76,30,32,31,244,31,94,31,203,31,83,31,17,31,17,30,23,31,81,31,227,31,227,30,242,31,58,31,124,31,251,31,87,31,87,30,215,31,250,31,240,31,240,30,240,29,95,31,16,31,16,30,195,31,162,31,75,31,136,31,136,30,136,29,77,31,77,30,186,31,204,31,204,30,69,31,69,30,130,31,112,31,18,31,24,31,24,30,24,29,45,31,104,31,127,31,192,31,192,30,55,31,58,31,136,31,179,31,179,30,225,31,225,30,99,31,48,31,160,31,41,31,121,31,121,30,183,31,27,31,27,30,151,31,89,31,86,31,136,31,178,31,139,31,204,31,240,31,37,31,216,31,216,30,70,31,70,30,169,31,169,30,145,31,126,31,115,31,164,31,64,31,64,30,58,31,198,31,237,31,47,31,138,31,155,31,30,31,220,31,153,31,196,31,95,31,124,31,125,31,54,31,158,31,89,31,236,31,217,31,225,31,225,30,225,29,87,31,237,31,237,30,177,31,177,30,157,31,156,31,207,31,207,30,177,31,213,31,123,31,123,30,216,31,183,31,183,30,41,31,8,31,8,30,103,31,88,31,61,31,27,31,222,31,64,31,250,31,3,31,28,31,43,31,238,31,137,31,208,31,26,31,189,31,243,31,51,31,51,30,51,29,8,31,8,30,8,29,24,31,29,31,29,30,8,31,240,31,134,31,147,31,230,31,28,31,28,30,103,31,214,31,8,31,158,31,158,30,192,31,186,31,13,31,122,31,55,31,214,31,51,31,239,31,177,31,177,30,177,29,112,31,63,31,162,31,126,31,32,31,144,31,237,31,237,30,200,31,224,31,71,31,132,31,242,31,117,31,82,31,82,30,226,31,190,31,113,31,202,31,96,31,32,31,145,31,145,30,145,29,17,31,17,30,173,31,45,31,213,31,161,31,144,31,55,31,55,30,202,31,50,31,117,31,22,31,126,31,126,30,169,31,92,31,92,30,92,29,47,31,8,31,8,30,217,31,181,31,181,30,29,31,198,31,211,31,211,30,218,31,218,30,144,31,220,31,255,31,255,30,19,31,199,31,117,31,14,31,72,31,16,31,40,31,223,31,122,31,154,31,172,31,109,31,159,31,159,30,114,31,18,31,18,30,122,31,177,31,95,31,179,31,179,30,65,31,224,31,118,31,67,31,10,31,116,31,75,31,252,31,98,31,24,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
