-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_942 is
end project_tb_942;

architecture project_tb_arch_942 of project_tb_942 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 291;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (9,0,154,0,104,0,147,0,16,0,20,0,92,0,134,0,77,0,146,0,15,0,202,0,75,0,0,0,129,0,58,0,29,0,149,0,237,0,224,0,133,0,78,0,151,0,192,0,0,0,0,0,54,0,0,0,82,0,0,0,99,0,0,0,38,0,0,0,0,0,156,0,233,0,0,0,0,0,19,0,22,0,41,0,65,0,46,0,129,0,25,0,229,0,139,0,0,0,54,0,0,0,5,0,245,0,241,0,46,0,0,0,110,0,195,0,0,0,113,0,3,0,229,0,164,0,3,0,116,0,0,0,0,0,228,0,51,0,104,0,123,0,64,0,254,0,0,0,245,0,112,0,98,0,52,0,150,0,0,0,69,0,184,0,0,0,135,0,0,0,77,0,38,0,120,0,207,0,55,0,51,0,0,0,221,0,254,0,94,0,28,0,0,0,34,0,82,0,0,0,55,0,168,0,67,0,80,0,156,0,32,0,131,0,97,0,0,0,80,0,243,0,6,0,182,0,82,0,0,0,130,0,237,0,56,0,226,0,0,0,87,0,208,0,14,0,0,0,76,0,163,0,163,0,238,0,190,0,166,0,56,0,209,0,0,0,75,0,65,0,69,0,102,0,8,0,55,0,127,0,0,0,0,0,0,0,181,0,215,0,147,0,0,0,0,0,130,0,200,0,235,0,125,0,216,0,160,0,0,0,0,0,242,0,3,0,136,0,246,0,243,0,0,0,89,0,238,0,130,0,43,0,40,0,0,0,0,0,141,0,0,0,200,0,252,0,0,0,201,0,202,0,155,0,178,0,253,0,15,0,210,0,20,0,27,0,213,0,2,0,192,0,154,0,75,0,97,0,20,0,12,0,0,0,0,0,165,0,20,0,254,0,179,0,56,0,79,0,92,0,232,0,98,0,62,0,143,0,5,0,39,0,131,0,233,0,213,0,238,0,0,0,237,0,0,0,17,0,90,0,0,0,139,0,167,0,48,0,12,0,45,0,220,0,127,0,0,0,178,0,239,0,3,0,179,0,0,0,13,0,23,0,169,0,160,0,217,0,245,0,24,0,13,0,51,0,98,0,130,0,168,0,71,0,217,0,161,0,4,0,109,0,0,0,196,0,199,0,117,0,0,0,97,0,213,0,117,0,0,0,104,0,41,0,183,0,0,0,174,0,196,0,185,0,38,0,247,0,142,0,68,0,171,0,4,0,225,0,72,0,200,0,188,0,0,0,73,0,8,0,0,0,196,0,0,0,91,0,166,0,152,0,100,0,180,0,224,0,191,0,218,0,56,0,169,0,3,0,175,0,253,0);
signal scenario_full  : scenario_type := (9,31,154,31,104,31,147,31,16,31,20,31,92,31,134,31,77,31,146,31,15,31,202,31,75,31,75,30,129,31,58,31,29,31,149,31,237,31,224,31,133,31,78,31,151,31,192,31,192,30,192,29,54,31,54,30,82,31,82,30,99,31,99,30,38,31,38,30,38,29,156,31,233,31,233,30,233,29,19,31,22,31,41,31,65,31,46,31,129,31,25,31,229,31,139,31,139,30,54,31,54,30,5,31,245,31,241,31,46,31,46,30,110,31,195,31,195,30,113,31,3,31,229,31,164,31,3,31,116,31,116,30,116,29,228,31,51,31,104,31,123,31,64,31,254,31,254,30,245,31,112,31,98,31,52,31,150,31,150,30,69,31,184,31,184,30,135,31,135,30,77,31,38,31,120,31,207,31,55,31,51,31,51,30,221,31,254,31,94,31,28,31,28,30,34,31,82,31,82,30,55,31,168,31,67,31,80,31,156,31,32,31,131,31,97,31,97,30,80,31,243,31,6,31,182,31,82,31,82,30,130,31,237,31,56,31,226,31,226,30,87,31,208,31,14,31,14,30,76,31,163,31,163,31,238,31,190,31,166,31,56,31,209,31,209,30,75,31,65,31,69,31,102,31,8,31,55,31,127,31,127,30,127,29,127,28,181,31,215,31,147,31,147,30,147,29,130,31,200,31,235,31,125,31,216,31,160,31,160,30,160,29,242,31,3,31,136,31,246,31,243,31,243,30,89,31,238,31,130,31,43,31,40,31,40,30,40,29,141,31,141,30,200,31,252,31,252,30,201,31,202,31,155,31,178,31,253,31,15,31,210,31,20,31,27,31,213,31,2,31,192,31,154,31,75,31,97,31,20,31,12,31,12,30,12,29,165,31,20,31,254,31,179,31,56,31,79,31,92,31,232,31,98,31,62,31,143,31,5,31,39,31,131,31,233,31,213,31,238,31,238,30,237,31,237,30,17,31,90,31,90,30,139,31,167,31,48,31,12,31,45,31,220,31,127,31,127,30,178,31,239,31,3,31,179,31,179,30,13,31,23,31,169,31,160,31,217,31,245,31,24,31,13,31,51,31,98,31,130,31,168,31,71,31,217,31,161,31,4,31,109,31,109,30,196,31,199,31,117,31,117,30,97,31,213,31,117,31,117,30,104,31,41,31,183,31,183,30,174,31,196,31,185,31,38,31,247,31,142,31,68,31,171,31,4,31,225,31,72,31,200,31,188,31,188,30,73,31,8,31,8,30,196,31,196,30,91,31,166,31,152,31,100,31,180,31,224,31,191,31,218,31,56,31,169,31,3,31,175,31,253,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
