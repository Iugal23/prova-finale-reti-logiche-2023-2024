-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_241 is
end project_tb_241;

architecture project_tb_arch_241 of project_tb_241 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 693;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (180,0,255,0,195,0,20,0,56,0,205,0,168,0,245,0,0,0,68,0,8,0,47,0,120,0,212,0,0,0,112,0,119,0,175,0,208,0,62,0,0,0,206,0,45,0,255,0,32,0,146,0,175,0,0,0,73,0,189,0,0,0,184,0,14,0,210,0,21,0,1,0,69,0,204,0,0,0,56,0,0,0,219,0,49,0,156,0,0,0,65,0,97,0,0,0,0,0,66,0,104,0,105,0,0,0,0,0,75,0,0,0,18,0,48,0,212,0,98,0,92,0,84,0,219,0,14,0,182,0,98,0,15,0,40,0,246,0,53,0,0,0,60,0,0,0,39,0,65,0,84,0,248,0,252,0,207,0,128,0,53,0,99,0,28,0,26,0,101,0,47,0,118,0,29,0,254,0,230,0,168,0,0,0,0,0,48,0,92,0,151,0,189,0,213,0,35,0,88,0,69,0,144,0,68,0,213,0,40,0,0,0,182,0,217,0,70,0,141,0,210,0,0,0,125,0,64,0,252,0,196,0,16,0,131,0,0,0,82,0,21,0,141,0,202,0,147,0,252,0,45,0,151,0,0,0,236,0,200,0,30,0,49,0,92,0,58,0,136,0,105,0,29,0,38,0,81,0,0,0,118,0,231,0,188,0,72,0,88,0,104,0,199,0,202,0,65,0,118,0,180,0,0,0,154,0,17,0,0,0,191,0,71,0,225,0,24,0,37,0,99,0,0,0,203,0,95,0,114,0,0,0,240,0,191,0,122,0,108,0,238,0,0,0,0,0,176,0,71,0,241,0,1,0,139,0,246,0,154,0,56,0,255,0,0,0,161,0,163,0,6,0,113,0,215,0,177,0,120,0,0,0,140,0,131,0,0,0,162,0,46,0,0,0,108,0,154,0,155,0,24,0,135,0,152,0,136,0,29,0,7,0,6,0,101,0,201,0,111,0,180,0,0,0,159,0,0,0,61,0,179,0,146,0,11,0,133,0,32,0,153,0,41,0,219,0,243,0,177,0,252,0,93,0,58,0,0,0,107,0,55,0,7,0,172,0,7,0,242,0,93,0,165,0,187,0,30,0,246,0,39,0,163,0,131,0,198,0,20,0,57,0,0,0,199,0,19,0,234,0,168,0,220,0,204,0,6,0,17,0,42,0,0,0,182,0,149,0,181,0,127,0,108,0,186,0,249,0,66,0,0,0,110,0,0,0,215,0,0,0,0,0,9,0,9,0,25,0,0,0,0,0,73,0,80,0,235,0,149,0,0,0,0,0,40,0,16,0,228,0,203,0,119,0,0,0,192,0,184,0,140,0,47,0,0,0,195,0,103,0,0,0,0,0,109,0,96,0,169,0,0,0,232,0,140,0,103,0,157,0,162,0,178,0,0,0,143,0,214,0,0,0,204,0,0,0,230,0,53,0,0,0,183,0,0,0,0,0,0,0,34,0,141,0,15,0,0,0,121,0,45,0,33,0,205,0,222,0,194,0,0,0,201,0,109,0,0,0,89,0,90,0,143,0,4,0,137,0,122,0,2,0,142,0,78,0,113,0,191,0,255,0,0,0,251,0,0,0,73,0,50,0,172,0,246,0,0,0,0,0,42,0,152,0,178,0,73,0,0,0,172,0,176,0,8,0,0,0,20,0,203,0,65,0,9,0,142,0,59,0,0,0,127,0,234,0,0,0,226,0,190,0,222,0,103,0,186,0,43,0,111,0,153,0,111,0,139,0,0,0,233,0,198,0,146,0,220,0,49,0,202,0,0,0,195,0,150,0,229,0,25,0,0,0,161,0,93,0,148,0,0,0,152,0,230,0,191,0,21,0,0,0,107,0,15,0,166,0,22,0,0,0,82,0,58,0,63,0,92,0,163,0,2,0,126,0,199,0,38,0,144,0,189,0,192,0,253,0,0,0,0,0,133,0,198,0,82,0,61,0,106,0,156,0,225,0,251,0,238,0,0,0,6,0,101,0,187,0,0,0,44,0,107,0,80,0,184,0,15,0,124,0,173,0,193,0,53,0,124,0,143,0,217,0,204,0,65,0,49,0,7,0,0,0,72,0,228,0,199,0,156,0,0,0,63,0,237,0,0,0,87,0,108,0,217,0,0,0,0,0,151,0,119,0,0,0,111,0,154,0,61,0,194,0,126,0,0,0,165,0,182,0,110,0,0,0,220,0,249,0,34,0,51,0,0,0,210,0,0,0,148,0,165,0,129,0,201,0,127,0,66,0,197,0,224,0,186,0,94,0,77,0,37,0,24,0,77,0,0,0,81,0,0,0,170,0,233,0,0,0,81,0,23,0,63,0,148,0,46,0,39,0,124,0,203,0,57,0,0,0,201,0,235,0,182,0,198,0,151,0,101,0,172,0,255,0,193,0,213,0,98,0,2,0,174,0,0,0,93,0,63,0,0,0,191,0,72,0,172,0,20,0,69,0,26,0,194,0,0,0,245,0,122,0,0,0,156,0,219,0,0,0,8,0,35,0,28,0,174,0,5,0,6,0,111,0,137,0,94,0,163,0,227,0,0,0,137,0,33,0,126,0,70,0,225,0,180,0,252,0,232,0,0,0,199,0,212,0,164,0,25,0,0,0,34,0,74,0,147,0,83,0,148,0,0,0,159,0,184,0,250,0,4,0,161,0,155,0,0,0,195,0,0,0,0,0,89,0,179,0,68,0,72,0,135,0,203,0,163,0,37,0,143,0,9,0,81,0,163,0,220,0,237,0,0,0,0,0,146,0,0,0,225,0,124,0,14,0,0,0,193,0,7,0,0,0,104,0,101,0,130,0,161,0,41,0,128,0,226,0,20,0,209,0,0,0,61,0,0,0,179,0,45,0,44,0,141,0,242,0,189,0,61,0,192,0,145,0,0,0,118,0,120,0,192,0,101,0,64,0,0,0,34,0,238,0,250,0,203,0,123,0,76,0,56,0,103,0,227,0,238,0,37,0,0,0,0,0,0,0,78,0,199,0,48,0,58,0,52,0,0,0,252,0,60,0,220,0,204,0,71,0,111,0,148,0,124,0,0,0,104,0,108,0,176,0,241,0,0,0,33,0,157,0,253,0,3,0,69,0,84,0,244,0,251,0,7,0,124,0,138,0,0,0,177,0);
signal scenario_full  : scenario_type := (180,31,255,31,195,31,20,31,56,31,205,31,168,31,245,31,245,30,68,31,8,31,47,31,120,31,212,31,212,30,112,31,119,31,175,31,208,31,62,31,62,30,206,31,45,31,255,31,32,31,146,31,175,31,175,30,73,31,189,31,189,30,184,31,14,31,210,31,21,31,1,31,69,31,204,31,204,30,56,31,56,30,219,31,49,31,156,31,156,30,65,31,97,31,97,30,97,29,66,31,104,31,105,31,105,30,105,29,75,31,75,30,18,31,48,31,212,31,98,31,92,31,84,31,219,31,14,31,182,31,98,31,15,31,40,31,246,31,53,31,53,30,60,31,60,30,39,31,65,31,84,31,248,31,252,31,207,31,128,31,53,31,99,31,28,31,26,31,101,31,47,31,118,31,29,31,254,31,230,31,168,31,168,30,168,29,48,31,92,31,151,31,189,31,213,31,35,31,88,31,69,31,144,31,68,31,213,31,40,31,40,30,182,31,217,31,70,31,141,31,210,31,210,30,125,31,64,31,252,31,196,31,16,31,131,31,131,30,82,31,21,31,141,31,202,31,147,31,252,31,45,31,151,31,151,30,236,31,200,31,30,31,49,31,92,31,58,31,136,31,105,31,29,31,38,31,81,31,81,30,118,31,231,31,188,31,72,31,88,31,104,31,199,31,202,31,65,31,118,31,180,31,180,30,154,31,17,31,17,30,191,31,71,31,225,31,24,31,37,31,99,31,99,30,203,31,95,31,114,31,114,30,240,31,191,31,122,31,108,31,238,31,238,30,238,29,176,31,71,31,241,31,1,31,139,31,246,31,154,31,56,31,255,31,255,30,161,31,163,31,6,31,113,31,215,31,177,31,120,31,120,30,140,31,131,31,131,30,162,31,46,31,46,30,108,31,154,31,155,31,24,31,135,31,152,31,136,31,29,31,7,31,6,31,101,31,201,31,111,31,180,31,180,30,159,31,159,30,61,31,179,31,146,31,11,31,133,31,32,31,153,31,41,31,219,31,243,31,177,31,252,31,93,31,58,31,58,30,107,31,55,31,7,31,172,31,7,31,242,31,93,31,165,31,187,31,30,31,246,31,39,31,163,31,131,31,198,31,20,31,57,31,57,30,199,31,19,31,234,31,168,31,220,31,204,31,6,31,17,31,42,31,42,30,182,31,149,31,181,31,127,31,108,31,186,31,249,31,66,31,66,30,110,31,110,30,215,31,215,30,215,29,9,31,9,31,25,31,25,30,25,29,73,31,80,31,235,31,149,31,149,30,149,29,40,31,16,31,228,31,203,31,119,31,119,30,192,31,184,31,140,31,47,31,47,30,195,31,103,31,103,30,103,29,109,31,96,31,169,31,169,30,232,31,140,31,103,31,157,31,162,31,178,31,178,30,143,31,214,31,214,30,204,31,204,30,230,31,53,31,53,30,183,31,183,30,183,29,183,28,34,31,141,31,15,31,15,30,121,31,45,31,33,31,205,31,222,31,194,31,194,30,201,31,109,31,109,30,89,31,90,31,143,31,4,31,137,31,122,31,2,31,142,31,78,31,113,31,191,31,255,31,255,30,251,31,251,30,73,31,50,31,172,31,246,31,246,30,246,29,42,31,152,31,178,31,73,31,73,30,172,31,176,31,8,31,8,30,20,31,203,31,65,31,9,31,142,31,59,31,59,30,127,31,234,31,234,30,226,31,190,31,222,31,103,31,186,31,43,31,111,31,153,31,111,31,139,31,139,30,233,31,198,31,146,31,220,31,49,31,202,31,202,30,195,31,150,31,229,31,25,31,25,30,161,31,93,31,148,31,148,30,152,31,230,31,191,31,21,31,21,30,107,31,15,31,166,31,22,31,22,30,82,31,58,31,63,31,92,31,163,31,2,31,126,31,199,31,38,31,144,31,189,31,192,31,253,31,253,30,253,29,133,31,198,31,82,31,61,31,106,31,156,31,225,31,251,31,238,31,238,30,6,31,101,31,187,31,187,30,44,31,107,31,80,31,184,31,15,31,124,31,173,31,193,31,53,31,124,31,143,31,217,31,204,31,65,31,49,31,7,31,7,30,72,31,228,31,199,31,156,31,156,30,63,31,237,31,237,30,87,31,108,31,217,31,217,30,217,29,151,31,119,31,119,30,111,31,154,31,61,31,194,31,126,31,126,30,165,31,182,31,110,31,110,30,220,31,249,31,34,31,51,31,51,30,210,31,210,30,148,31,165,31,129,31,201,31,127,31,66,31,197,31,224,31,186,31,94,31,77,31,37,31,24,31,77,31,77,30,81,31,81,30,170,31,233,31,233,30,81,31,23,31,63,31,148,31,46,31,39,31,124,31,203,31,57,31,57,30,201,31,235,31,182,31,198,31,151,31,101,31,172,31,255,31,193,31,213,31,98,31,2,31,174,31,174,30,93,31,63,31,63,30,191,31,72,31,172,31,20,31,69,31,26,31,194,31,194,30,245,31,122,31,122,30,156,31,219,31,219,30,8,31,35,31,28,31,174,31,5,31,6,31,111,31,137,31,94,31,163,31,227,31,227,30,137,31,33,31,126,31,70,31,225,31,180,31,252,31,232,31,232,30,199,31,212,31,164,31,25,31,25,30,34,31,74,31,147,31,83,31,148,31,148,30,159,31,184,31,250,31,4,31,161,31,155,31,155,30,195,31,195,30,195,29,89,31,179,31,68,31,72,31,135,31,203,31,163,31,37,31,143,31,9,31,81,31,163,31,220,31,237,31,237,30,237,29,146,31,146,30,225,31,124,31,14,31,14,30,193,31,7,31,7,30,104,31,101,31,130,31,161,31,41,31,128,31,226,31,20,31,209,31,209,30,61,31,61,30,179,31,45,31,44,31,141,31,242,31,189,31,61,31,192,31,145,31,145,30,118,31,120,31,192,31,101,31,64,31,64,30,34,31,238,31,250,31,203,31,123,31,76,31,56,31,103,31,227,31,238,31,37,31,37,30,37,29,37,28,78,31,199,31,48,31,58,31,52,31,52,30,252,31,60,31,220,31,204,31,71,31,111,31,148,31,124,31,124,30,104,31,108,31,176,31,241,31,241,30,33,31,157,31,253,31,3,31,69,31,84,31,244,31,251,31,7,31,124,31,138,31,138,30,177,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
