-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 346;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,103,0,222,0,0,0,214,0,9,0,52,0,183,0,24,0,215,0,140,0,89,0,214,0,102,0,255,0,26,0,86,0,148,0,69,0,34,0,84,0,236,0,147,0,84,0,38,0,71,0,0,0,177,0,72,0,155,0,0,0,167,0,215,0,0,0,45,0,255,0,119,0,165,0,207,0,91,0,41,0,227,0,51,0,165,0,79,0,37,0,77,0,243,0,23,0,216,0,204,0,0,0,105,0,73,0,55,0,65,0,0,0,142,0,118,0,0,0,63,0,157,0,62,0,41,0,96,0,69,0,245,0,152,0,0,0,37,0,32,0,102,0,54,0,38,0,0,0,192,0,127,0,0,0,0,0,60,0,126,0,167,0,55,0,0,0,185,0,184,0,66,0,151,0,153,0,146,0,181,0,0,0,197,0,220,0,164,0,5,0,35,0,70,0,223,0,0,0,0,0,25,0,0,0,94,0,236,0,113,0,0,0,250,0,204,0,18,0,173,0,45,0,135,0,250,0,139,0,228,0,173,0,0,0,0,0,48,0,101,0,143,0,142,0,110,0,152,0,0,0,107,0,146,0,139,0,106,0,125,0,0,0,168,0,163,0,116,0,91,0,187,0,65,0,84,0,67,0,205,0,233,0,253,0,0,0,111,0,67,0,0,0,186,0,87,0,249,0,85,0,131,0,133,0,133,0,13,0,161,0,43,0,45,0,0,0,85,0,163,0,146,0,217,0,213,0,0,0,26,0,214,0,82,0,74,0,0,0,16,0,104,0,0,0,114,0,212,0,0,0,147,0,34,0,115,0,228,0,215,0,42,0,0,0,81,0,202,0,181,0,18,0,147,0,29,0,40,0,45,0,191,0,0,0,120,0,26,0,66,0,0,0,93,0,26,0,113,0,109,0,193,0,107,0,0,0,0,0,158,0,0,0,231,0,79,0,245,0,226,0,0,0,70,0,229,0,0,0,135,0,167,0,165,0,0,0,86,0,90,0,0,0,238,0,0,0,0,0,147,0,157,0,0,0,146,0,21,0,106,0,204,0,0,0,225,0,215,0,81,0,217,0,128,0,130,0,219,0,10,0,80,0,187,0,0,0,87,0,183,0,232,0,6,0,0,0,87,0,0,0,0,0,152,0,162,0,133,0,132,0,0,0,196,0,150,0,207,0,114,0,0,0,133,0,0,0,0,0,223,0,134,0,0,0,217,0,0,0,22,0,138,0,137,0,0,0,32,0,103,0,150,0,251,0,6,0,25,0,183,0,97,0,197,0,0,0,216,0,8,0,92,0,237,0,64,0,245,0,0,0,0,0,0,0,67,0,238,0,186,0,206,0,217,0,49,0,120,0,61,0,144,0,202,0,166,0,114,0,188,0,122,0,0,0,79,0,232,0,148,0,91,0,174,0,194,0,82,0,182,0,15,0,204,0,235,0,129,0,219,0,0,0,65,0,112,0,139,0,82,0,240,0,144,0,82,0,171,0,219,0,120,0,164,0,123,0,246,0,0,0,70,0,0,0,35,0,229,0,12,0,27,0,0,0,161,0,58,0);
signal scenario_full  : scenario_type := (0,0,0,0,103,31,222,31,222,30,214,31,9,31,52,31,183,31,24,31,215,31,140,31,89,31,214,31,102,31,255,31,26,31,86,31,148,31,69,31,34,31,84,31,236,31,147,31,84,31,38,31,71,31,71,30,177,31,72,31,155,31,155,30,167,31,215,31,215,30,45,31,255,31,119,31,165,31,207,31,91,31,41,31,227,31,51,31,165,31,79,31,37,31,77,31,243,31,23,31,216,31,204,31,204,30,105,31,73,31,55,31,65,31,65,30,142,31,118,31,118,30,63,31,157,31,62,31,41,31,96,31,69,31,245,31,152,31,152,30,37,31,32,31,102,31,54,31,38,31,38,30,192,31,127,31,127,30,127,29,60,31,126,31,167,31,55,31,55,30,185,31,184,31,66,31,151,31,153,31,146,31,181,31,181,30,197,31,220,31,164,31,5,31,35,31,70,31,223,31,223,30,223,29,25,31,25,30,94,31,236,31,113,31,113,30,250,31,204,31,18,31,173,31,45,31,135,31,250,31,139,31,228,31,173,31,173,30,173,29,48,31,101,31,143,31,142,31,110,31,152,31,152,30,107,31,146,31,139,31,106,31,125,31,125,30,168,31,163,31,116,31,91,31,187,31,65,31,84,31,67,31,205,31,233,31,253,31,253,30,111,31,67,31,67,30,186,31,87,31,249,31,85,31,131,31,133,31,133,31,13,31,161,31,43,31,45,31,45,30,85,31,163,31,146,31,217,31,213,31,213,30,26,31,214,31,82,31,74,31,74,30,16,31,104,31,104,30,114,31,212,31,212,30,147,31,34,31,115,31,228,31,215,31,42,31,42,30,81,31,202,31,181,31,18,31,147,31,29,31,40,31,45,31,191,31,191,30,120,31,26,31,66,31,66,30,93,31,26,31,113,31,109,31,193,31,107,31,107,30,107,29,158,31,158,30,231,31,79,31,245,31,226,31,226,30,70,31,229,31,229,30,135,31,167,31,165,31,165,30,86,31,90,31,90,30,238,31,238,30,238,29,147,31,157,31,157,30,146,31,21,31,106,31,204,31,204,30,225,31,215,31,81,31,217,31,128,31,130,31,219,31,10,31,80,31,187,31,187,30,87,31,183,31,232,31,6,31,6,30,87,31,87,30,87,29,152,31,162,31,133,31,132,31,132,30,196,31,150,31,207,31,114,31,114,30,133,31,133,30,133,29,223,31,134,31,134,30,217,31,217,30,22,31,138,31,137,31,137,30,32,31,103,31,150,31,251,31,6,31,25,31,183,31,97,31,197,31,197,30,216,31,8,31,92,31,237,31,64,31,245,31,245,30,245,29,245,28,67,31,238,31,186,31,206,31,217,31,49,31,120,31,61,31,144,31,202,31,166,31,114,31,188,31,122,31,122,30,79,31,232,31,148,31,91,31,174,31,194,31,82,31,182,31,15,31,204,31,235,31,129,31,219,31,219,30,65,31,112,31,139,31,82,31,240,31,144,31,82,31,171,31,219,31,120,31,164,31,123,31,246,31,246,30,70,31,70,30,35,31,229,31,12,31,27,31,27,30,161,31,58,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
