-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 890;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (190,0,28,0,0,0,99,0,194,0,156,0,0,0,253,0,131,0,0,0,0,0,225,0,162,0,169,0,37,0,101,0,82,0,37,0,0,0,0,0,13,0,172,0,61,0,0,0,229,0,226,0,0,0,151,0,42,0,94,0,0,0,164,0,88,0,10,0,0,0,105,0,0,0,0,0,0,0,156,0,0,0,110,0,9,0,222,0,157,0,0,0,9,0,0,0,131,0,197,0,106,0,0,0,229,0,58,0,0,0,203,0,220,0,198,0,146,0,0,0,0,0,83,0,9,0,149,0,6,0,12,0,0,0,77,0,0,0,155,0,94,0,192,0,0,0,187,0,232,0,238,0,0,0,46,0,209,0,54,0,30,0,0,0,98,0,118,0,0,0,151,0,253,0,135,0,180,0,0,0,115,0,113,0,15,0,0,0,0,0,144,0,64,0,50,0,222,0,84,0,190,0,67,0,136,0,44,0,81,0,75,0,0,0,0,0,0,0,42,0,0,0,0,0,202,0,229,0,85,0,79,0,42,0,79,0,98,0,0,0,27,0,34,0,126,0,108,0,114,0,207,0,216,0,119,0,167,0,0,0,117,0,47,0,242,0,0,0,79,0,131,0,63,0,151,0,78,0,0,0,248,0,112,0,159,0,8,0,248,0,114,0,0,0,0,0,213,0,215,0,67,0,88,0,110,0,25,0,0,0,0,0,0,0,228,0,43,0,77,0,0,0,134,0,35,0,163,0,40,0,164,0,85,0,0,0,0,0,85,0,220,0,116,0,128,0,142,0,225,0,0,0,176,0,101,0,143,0,24,0,196,0,0,0,186,0,202,0,0,0,169,0,102,0,12,0,0,0,127,0,147,0,207,0,0,0,80,0,73,0,0,0,55,0,185,0,127,0,93,0,241,0,197,0,42,0,192,0,232,0,110,0,195,0,192,0,39,0,113,0,66,0,208,0,251,0,0,0,71,0,0,0,110,0,24,0,0,0,28,0,184,0,145,0,128,0,79,0,6,0,0,0,200,0,230,0,254,0,239,0,222,0,116,0,227,0,213,0,36,0,216,0,60,0,117,0,215,0,179,0,157,0,241,0,36,0,0,0,228,0,25,0,229,0,202,0,79,0,83,0,170,0,236,0,212,0,79,0,194,0,110,0,49,0,227,0,189,0,69,0,0,0,37,0,184,0,206,0,62,0,177,0,0,0,245,0,140,0,0,0,0,0,0,0,197,0,0,0,0,0,196,0,38,0,29,0,147,0,0,0,131,0,115,0,114,0,0,0,0,0,211,0,45,0,12,0,172,0,3,0,223,0,91,0,160,0,246,0,0,0,3,0,17,0,0,0,158,0,94,0,0,0,207,0,7,0,171,0,0,0,194,0,222,0,71,0,0,0,164,0,133,0,0,0,0,0,40,0,196,0,96,0,82,0,227,0,83,0,177,0,34,0,84,0,56,0,98,0,161,0,183,0,0,0,104,0,66,0,0,0,121,0,188,0,180,0,251,0,190,0,0,0,254,0,83,0,204,0,171,0,0,0,156,0,51,0,135,0,207,0,234,0,117,0,90,0,3,0,253,0,0,0,111,0,112,0,112,0,0,0,224,0,0,0,0,0,172,0,37,0,242,0,0,0,19,0,0,0,85,0,74,0,0,0,160,0,255,0,0,0,110,0,175,0,0,0,36,0,138,0,0,0,114,0,5,0,198,0,201,0,57,0,236,0,63,0,33,0,138,0,0,0,14,0,142,0,96,0,179,0,0,0,112,0,73,0,8,0,0,0,64,0,24,0,179,0,128,0,45,0,0,0,126,0,0,0,191,0,17,0,202,0,0,0,0,0,119,0,26,0,145,0,0,0,129,0,220,0,193,0,56,0,0,0,193,0,119,0,255,0,113,0,83,0,64,0,175,0,247,0,167,0,176,0,187,0,0,0,127,0,210,0,109,0,71,0,131,0,54,0,235,0,0,0,7,0,194,0,53,0,79,0,240,0,246,0,57,0,156,0,144,0,43,0,8,0,214,0,0,0,85,0,193,0,239,0,70,0,109,0,190,0,14,0,121,0,26,0,168,0,129,0,214,0,23,0,0,0,220,0,0,0,3,0,105,0,213,0,119,0,36,0,151,0,201,0,0,0,205,0,197,0,0,0,199,0,36,0,21,0,0,0,0,0,142,0,244,0,196,0,162,0,183,0,10,0,155,0,0,0,34,0,214,0,241,0,247,0,139,0,0,0,47,0,0,0,49,0,234,0,200,0,61,0,0,0,0,0,153,0,225,0,32,0,171,0,246,0,90,0,109,0,0,0,150,0,26,0,191,0,232,0,0,0,253,0,59,0,154,0,72,0,185,0,204,0,112,0,48,0,203,0,219,0,85,0,36,0,20,0,166,0,56,0,184,0,140,0,13,0,0,0,188,0,177,0,254,0,43,0,42,0,138,0,246,0,93,0,0,0,87,0,150,0,150,0,32,0,207,0,142,0,0,0,67,0,164,0,59,0,40,0,55,0,43,0,91,0,40,0,0,0,254,0,144,0,143,0,193,0,0,0,203,0,47,0,26,0,55,0,135,0,127,0,165,0,201,0,131,0,183,0,0,0,155,0,222,0,0,0,29,0,124,0,30,0,173,0,0,0,0,0,176,0,25,0,0,0,0,0,238,0,54,0,8,0,108,0,136,0,170,0,0,0,57,0,0,0,158,0,27,0,143,0,0,0,0,0,43,0,0,0,146,0,229,0,187,0,221,0,0,0,0,0,0,0,243,0,0,0,53,0,124,0,89,0,46,0,0,0,0,0,252,0,161,0,39,0,0,0,218,0,233,0,0,0,6,0,34,0,137,0,109,0,60,0,98,0,172,0,229,0,157,0,192,0,46,0,60,0,201,0,7,0,163,0,238,0,221,0,128,0,15,0,186,0,184,0,198,0,125,0,149,0,0,0,0,0,0,0,0,0,248,0,179,0,180,0,94,0,66,0,234,0,207,0,129,0,232,0,0,0,221,0,89,0,243,0,0,0,29,0,250,0,129,0,151,0,190,0,44,0,211,0,221,0,235,0,15,0,36,0,90,0,0,0,170,0,198,0,59,0,0,0,233,0,208,0,0,0,32,0,173,0,98,0,39,0,182,0,0,0,161,0,156,0,39,0,223,0,4,0,243,0,106,0,0,0,19,0,51,0,15,0,107,0,84,0,209,0,152,0,38,0,0,0,190,0,228,0,132,0,0,0,0,0,232,0,0,0,203,0,243,0,244,0,20,0,0,0,0,0,9,0,101,0,115,0,0,0,178,0,162,0,0,0,55,0,0,0,55,0,0,0,187,0,23,0,0,0,163,0,151,0,170,0,73,0,82,0,26,0,0,0,49,0,192,0,0,0,253,0,163,0,16,0,31,0,181,0,117,0,21,0,56,0,251,0,112,0,6,0,0,0,133,0,0,0,7,0,154,0,17,0,0,0,239,0,151,0,18,0,96,0,64,0,80,0,228,0,0,0,73,0,0,0,113,0,228,0,237,0,159,0,60,0,167,0,0,0,0,0,105,0,183,0,0,0,49,0,209,0,132,0,70,0,114,0,191,0,174,0,214,0,0,0,243,0,231,0,0,0,235,0,0,0,0,0,0,0,123,0,4,0,70,0,180,0,212,0,231,0,214,0,90,0,247,0,0,0,48,0,172,0,138,0,163,0,0,0,46,0,0,0,0,0,107,0,29,0,0,0,161,0,0,0,53,0,194,0,0,0,145,0,0,0,244,0,40,0,84,0,78,0,192,0,62,0,0,0,83,0,152,0,0,0,0,0,232,0,0,0,150,0,171,0,48,0,165,0,176,0,0,0,255,0,0,0,139,0,29,0,241,0,159,0,150,0,0,0,94,0,61,0,30,0,207,0,148,0,30,0,140,0,246,0,0,0,71,0,144,0,0,0,144,0,158,0,144,0,147,0,172,0,213,0,2,0,180,0,0,0,152,0,28,0,79,0,26,0,0,0,98,0,0,0,167,0,0,0);
signal scenario_full  : scenario_type := (190,31,28,31,28,30,99,31,194,31,156,31,156,30,253,31,131,31,131,30,131,29,225,31,162,31,169,31,37,31,101,31,82,31,37,31,37,30,37,29,13,31,172,31,61,31,61,30,229,31,226,31,226,30,151,31,42,31,94,31,94,30,164,31,88,31,10,31,10,30,105,31,105,30,105,29,105,28,156,31,156,30,110,31,9,31,222,31,157,31,157,30,9,31,9,30,131,31,197,31,106,31,106,30,229,31,58,31,58,30,203,31,220,31,198,31,146,31,146,30,146,29,83,31,9,31,149,31,6,31,12,31,12,30,77,31,77,30,155,31,94,31,192,31,192,30,187,31,232,31,238,31,238,30,46,31,209,31,54,31,30,31,30,30,98,31,118,31,118,30,151,31,253,31,135,31,180,31,180,30,115,31,113,31,15,31,15,30,15,29,144,31,64,31,50,31,222,31,84,31,190,31,67,31,136,31,44,31,81,31,75,31,75,30,75,29,75,28,42,31,42,30,42,29,202,31,229,31,85,31,79,31,42,31,79,31,98,31,98,30,27,31,34,31,126,31,108,31,114,31,207,31,216,31,119,31,167,31,167,30,117,31,47,31,242,31,242,30,79,31,131,31,63,31,151,31,78,31,78,30,248,31,112,31,159,31,8,31,248,31,114,31,114,30,114,29,213,31,215,31,67,31,88,31,110,31,25,31,25,30,25,29,25,28,228,31,43,31,77,31,77,30,134,31,35,31,163,31,40,31,164,31,85,31,85,30,85,29,85,31,220,31,116,31,128,31,142,31,225,31,225,30,176,31,101,31,143,31,24,31,196,31,196,30,186,31,202,31,202,30,169,31,102,31,12,31,12,30,127,31,147,31,207,31,207,30,80,31,73,31,73,30,55,31,185,31,127,31,93,31,241,31,197,31,42,31,192,31,232,31,110,31,195,31,192,31,39,31,113,31,66,31,208,31,251,31,251,30,71,31,71,30,110,31,24,31,24,30,28,31,184,31,145,31,128,31,79,31,6,31,6,30,200,31,230,31,254,31,239,31,222,31,116,31,227,31,213,31,36,31,216,31,60,31,117,31,215,31,179,31,157,31,241,31,36,31,36,30,228,31,25,31,229,31,202,31,79,31,83,31,170,31,236,31,212,31,79,31,194,31,110,31,49,31,227,31,189,31,69,31,69,30,37,31,184,31,206,31,62,31,177,31,177,30,245,31,140,31,140,30,140,29,140,28,197,31,197,30,197,29,196,31,38,31,29,31,147,31,147,30,131,31,115,31,114,31,114,30,114,29,211,31,45,31,12,31,172,31,3,31,223,31,91,31,160,31,246,31,246,30,3,31,17,31,17,30,158,31,94,31,94,30,207,31,7,31,171,31,171,30,194,31,222,31,71,31,71,30,164,31,133,31,133,30,133,29,40,31,196,31,96,31,82,31,227,31,83,31,177,31,34,31,84,31,56,31,98,31,161,31,183,31,183,30,104,31,66,31,66,30,121,31,188,31,180,31,251,31,190,31,190,30,254,31,83,31,204,31,171,31,171,30,156,31,51,31,135,31,207,31,234,31,117,31,90,31,3,31,253,31,253,30,111,31,112,31,112,31,112,30,224,31,224,30,224,29,172,31,37,31,242,31,242,30,19,31,19,30,85,31,74,31,74,30,160,31,255,31,255,30,110,31,175,31,175,30,36,31,138,31,138,30,114,31,5,31,198,31,201,31,57,31,236,31,63,31,33,31,138,31,138,30,14,31,142,31,96,31,179,31,179,30,112,31,73,31,8,31,8,30,64,31,24,31,179,31,128,31,45,31,45,30,126,31,126,30,191,31,17,31,202,31,202,30,202,29,119,31,26,31,145,31,145,30,129,31,220,31,193,31,56,31,56,30,193,31,119,31,255,31,113,31,83,31,64,31,175,31,247,31,167,31,176,31,187,31,187,30,127,31,210,31,109,31,71,31,131,31,54,31,235,31,235,30,7,31,194,31,53,31,79,31,240,31,246,31,57,31,156,31,144,31,43,31,8,31,214,31,214,30,85,31,193,31,239,31,70,31,109,31,190,31,14,31,121,31,26,31,168,31,129,31,214,31,23,31,23,30,220,31,220,30,3,31,105,31,213,31,119,31,36,31,151,31,201,31,201,30,205,31,197,31,197,30,199,31,36,31,21,31,21,30,21,29,142,31,244,31,196,31,162,31,183,31,10,31,155,31,155,30,34,31,214,31,241,31,247,31,139,31,139,30,47,31,47,30,49,31,234,31,200,31,61,31,61,30,61,29,153,31,225,31,32,31,171,31,246,31,90,31,109,31,109,30,150,31,26,31,191,31,232,31,232,30,253,31,59,31,154,31,72,31,185,31,204,31,112,31,48,31,203,31,219,31,85,31,36,31,20,31,166,31,56,31,184,31,140,31,13,31,13,30,188,31,177,31,254,31,43,31,42,31,138,31,246,31,93,31,93,30,87,31,150,31,150,31,32,31,207,31,142,31,142,30,67,31,164,31,59,31,40,31,55,31,43,31,91,31,40,31,40,30,254,31,144,31,143,31,193,31,193,30,203,31,47,31,26,31,55,31,135,31,127,31,165,31,201,31,131,31,183,31,183,30,155,31,222,31,222,30,29,31,124,31,30,31,173,31,173,30,173,29,176,31,25,31,25,30,25,29,238,31,54,31,8,31,108,31,136,31,170,31,170,30,57,31,57,30,158,31,27,31,143,31,143,30,143,29,43,31,43,30,146,31,229,31,187,31,221,31,221,30,221,29,221,28,243,31,243,30,53,31,124,31,89,31,46,31,46,30,46,29,252,31,161,31,39,31,39,30,218,31,233,31,233,30,6,31,34,31,137,31,109,31,60,31,98,31,172,31,229,31,157,31,192,31,46,31,60,31,201,31,7,31,163,31,238,31,221,31,128,31,15,31,186,31,184,31,198,31,125,31,149,31,149,30,149,29,149,28,149,27,248,31,179,31,180,31,94,31,66,31,234,31,207,31,129,31,232,31,232,30,221,31,89,31,243,31,243,30,29,31,250,31,129,31,151,31,190,31,44,31,211,31,221,31,235,31,15,31,36,31,90,31,90,30,170,31,198,31,59,31,59,30,233,31,208,31,208,30,32,31,173,31,98,31,39,31,182,31,182,30,161,31,156,31,39,31,223,31,4,31,243,31,106,31,106,30,19,31,51,31,15,31,107,31,84,31,209,31,152,31,38,31,38,30,190,31,228,31,132,31,132,30,132,29,232,31,232,30,203,31,243,31,244,31,20,31,20,30,20,29,9,31,101,31,115,31,115,30,178,31,162,31,162,30,55,31,55,30,55,31,55,30,187,31,23,31,23,30,163,31,151,31,170,31,73,31,82,31,26,31,26,30,49,31,192,31,192,30,253,31,163,31,16,31,31,31,181,31,117,31,21,31,56,31,251,31,112,31,6,31,6,30,133,31,133,30,7,31,154,31,17,31,17,30,239,31,151,31,18,31,96,31,64,31,80,31,228,31,228,30,73,31,73,30,113,31,228,31,237,31,159,31,60,31,167,31,167,30,167,29,105,31,183,31,183,30,49,31,209,31,132,31,70,31,114,31,191,31,174,31,214,31,214,30,243,31,231,31,231,30,235,31,235,30,235,29,235,28,123,31,4,31,70,31,180,31,212,31,231,31,214,31,90,31,247,31,247,30,48,31,172,31,138,31,163,31,163,30,46,31,46,30,46,29,107,31,29,31,29,30,161,31,161,30,53,31,194,31,194,30,145,31,145,30,244,31,40,31,84,31,78,31,192,31,62,31,62,30,83,31,152,31,152,30,152,29,232,31,232,30,150,31,171,31,48,31,165,31,176,31,176,30,255,31,255,30,139,31,29,31,241,31,159,31,150,31,150,30,94,31,61,31,30,31,207,31,148,31,30,31,140,31,246,31,246,30,71,31,144,31,144,30,144,31,158,31,144,31,147,31,172,31,213,31,2,31,180,31,180,30,152,31,28,31,79,31,26,31,26,30,98,31,98,30,167,31,167,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
