-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 402;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (191,0,0,0,211,0,62,0,40,0,0,0,173,0,28,0,90,0,60,0,0,0,3,0,126,0,225,0,159,0,0,0,179,0,0,0,137,0,34,0,73,0,120,0,5,0,64,0,226,0,234,0,254,0,194,0,0,0,63,0,0,0,48,0,193,0,11,0,111,0,0,0,213,0,12,0,155,0,141,0,100,0,56,0,97,0,0,0,113,0,40,0,134,0,160,0,12,0,0,0,205,0,80,0,255,0,205,0,0,0,0,0,50,0,66,0,175,0,149,0,153,0,179,0,183,0,195,0,145,0,0,0,115,0,206,0,0,0,0,0,0,0,180,0,77,0,49,0,67,0,0,0,0,0,159,0,0,0,123,0,81,0,136,0,204,0,0,0,68,0,209,0,0,0,148,0,212,0,140,0,80,0,0,0,220,0,251,0,214,0,236,0,0,0,213,0,0,0,0,0,180,0,105,0,0,0,7,0,0,0,171,0,0,0,90,0,0,0,124,0,11,0,61,0,43,0,178,0,0,0,230,0,178,0,97,0,175,0,34,0,27,0,211,0,6,0,187,0,146,0,121,0,153,0,192,0,70,0,199,0,105,0,90,0,9,0,141,0,97,0,214,0,0,0,237,0,167,0,35,0,32,0,0,0,103,0,100,0,0,0,195,0,108,0,103,0,110,0,0,0,0,0,180,0,207,0,79,0,159,0,0,0,95,0,71,0,0,0,0,0,55,0,26,0,249,0,246,0,208,0,234,0,0,0,0,0,11,0,223,0,88,0,98,0,130,0,0,0,18,0,136,0,158,0,181,0,124,0,82,0,233,0,93,0,253,0,43,0,22,0,38,0,0,0,168,0,17,0,208,0,136,0,161,0,123,0,129,0,65,0,194,0,29,0,0,0,1,0,0,0,223,0,172,0,134,0,0,0,132,0,0,0,176,0,245,0,188,0,0,0,167,0,0,0,0,0,147,0,123,0,151,0,242,0,129,0,124,0,71,0,0,0,0,0,189,0,224,0,248,0,198,0,0,0,198,0,46,0,90,0,156,0,8,0,220,0,16,0,162,0,3,0,0,0,200,0,82,0,109,0,0,0,0,0,117,0,249,0,109,0,85,0,56,0,224,0,52,0,45,0,201,0,118,0,29,0,0,0,6,0,1,0,0,0,3,0,0,0,241,0,170,0,0,0,60,0,80,0,253,0,21,0,250,0,177,0,159,0,0,0,194,0,105,0,108,0,63,0,140,0,36,0,102,0,47,0,224,0,149,0,139,0,161,0,164,0,118,0,98,0,154,0,194,0,217,0,31,0,19,0,23,0,143,0,70,0,70,0,128,0,219,0,216,0,230,0,0,0,169,0,93,0,112,0,200,0,222,0,4,0,196,0,0,0,0,0,105,0,54,0,0,0,72,0,160,0,107,0,190,0,253,0,76,0,186,0,171,0,111,0,204,0,0,0,243,0,0,0,208,0,203,0,180,0,0,0,21,0,173,0,87,0,24,0,18,0,145,0,77,0,112,0,0,0,24,0,72,0,0,0,0,0,132,0,218,0,214,0,0,0,168,0,133,0,56,0,152,0,189,0,148,0,221,0,0,0,0,0,61,0,148,0,232,0,74,0,164,0,105,0,136,0,0,0,154,0,0,0,95,0,0,0,174,0,116,0,195,0,58,0,190,0,189,0,64,0,6,0,225,0,196,0,12,0,126,0,113,0,180,0,76,0,219,0,23,0,0,0,27,0,82,0,0,0,0,0,178,0,45,0,166,0,249,0,85,0,214,0,105,0,88,0,228,0,0,0,0,0,236,0,56,0,0,0);
signal scenario_full  : scenario_type := (191,31,191,30,211,31,62,31,40,31,40,30,173,31,28,31,90,31,60,31,60,30,3,31,126,31,225,31,159,31,159,30,179,31,179,30,137,31,34,31,73,31,120,31,5,31,64,31,226,31,234,31,254,31,194,31,194,30,63,31,63,30,48,31,193,31,11,31,111,31,111,30,213,31,12,31,155,31,141,31,100,31,56,31,97,31,97,30,113,31,40,31,134,31,160,31,12,31,12,30,205,31,80,31,255,31,205,31,205,30,205,29,50,31,66,31,175,31,149,31,153,31,179,31,183,31,195,31,145,31,145,30,115,31,206,31,206,30,206,29,206,28,180,31,77,31,49,31,67,31,67,30,67,29,159,31,159,30,123,31,81,31,136,31,204,31,204,30,68,31,209,31,209,30,148,31,212,31,140,31,80,31,80,30,220,31,251,31,214,31,236,31,236,30,213,31,213,30,213,29,180,31,105,31,105,30,7,31,7,30,171,31,171,30,90,31,90,30,124,31,11,31,61,31,43,31,178,31,178,30,230,31,178,31,97,31,175,31,34,31,27,31,211,31,6,31,187,31,146,31,121,31,153,31,192,31,70,31,199,31,105,31,90,31,9,31,141,31,97,31,214,31,214,30,237,31,167,31,35,31,32,31,32,30,103,31,100,31,100,30,195,31,108,31,103,31,110,31,110,30,110,29,180,31,207,31,79,31,159,31,159,30,95,31,71,31,71,30,71,29,55,31,26,31,249,31,246,31,208,31,234,31,234,30,234,29,11,31,223,31,88,31,98,31,130,31,130,30,18,31,136,31,158,31,181,31,124,31,82,31,233,31,93,31,253,31,43,31,22,31,38,31,38,30,168,31,17,31,208,31,136,31,161,31,123,31,129,31,65,31,194,31,29,31,29,30,1,31,1,30,223,31,172,31,134,31,134,30,132,31,132,30,176,31,245,31,188,31,188,30,167,31,167,30,167,29,147,31,123,31,151,31,242,31,129,31,124,31,71,31,71,30,71,29,189,31,224,31,248,31,198,31,198,30,198,31,46,31,90,31,156,31,8,31,220,31,16,31,162,31,3,31,3,30,200,31,82,31,109,31,109,30,109,29,117,31,249,31,109,31,85,31,56,31,224,31,52,31,45,31,201,31,118,31,29,31,29,30,6,31,1,31,1,30,3,31,3,30,241,31,170,31,170,30,60,31,80,31,253,31,21,31,250,31,177,31,159,31,159,30,194,31,105,31,108,31,63,31,140,31,36,31,102,31,47,31,224,31,149,31,139,31,161,31,164,31,118,31,98,31,154,31,194,31,217,31,31,31,19,31,23,31,143,31,70,31,70,31,128,31,219,31,216,31,230,31,230,30,169,31,93,31,112,31,200,31,222,31,4,31,196,31,196,30,196,29,105,31,54,31,54,30,72,31,160,31,107,31,190,31,253,31,76,31,186,31,171,31,111,31,204,31,204,30,243,31,243,30,208,31,203,31,180,31,180,30,21,31,173,31,87,31,24,31,18,31,145,31,77,31,112,31,112,30,24,31,72,31,72,30,72,29,132,31,218,31,214,31,214,30,168,31,133,31,56,31,152,31,189,31,148,31,221,31,221,30,221,29,61,31,148,31,232,31,74,31,164,31,105,31,136,31,136,30,154,31,154,30,95,31,95,30,174,31,116,31,195,31,58,31,190,31,189,31,64,31,6,31,225,31,196,31,12,31,126,31,113,31,180,31,76,31,219,31,23,31,23,30,27,31,82,31,82,30,82,29,178,31,45,31,166,31,249,31,85,31,214,31,105,31,88,31,228,31,228,30,228,29,236,31,56,31,56,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
