-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_549 is
end project_tb_549;

architecture project_tb_arch_549 of project_tb_549 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 919;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (218,0,187,0,141,0,163,0,121,0,86,0,196,0,81,0,0,0,0,0,6,0,73,0,249,0,71,0,25,0,223,0,145,0,178,0,129,0,200,0,170,0,7,0,0,0,77,0,22,0,156,0,144,0,175,0,0,0,35,0,97,0,180,0,94,0,103,0,245,0,0,0,2,0,246,0,150,0,212,0,0,0,185,0,152,0,12,0,54,0,0,0,57,0,166,0,51,0,0,0,41,0,215,0,80,0,1,0,6,0,21,0,233,0,251,0,211,0,0,0,26,0,19,0,0,0,207,0,0,0,0,0,246,0,16,0,36,0,99,0,114,0,118,0,185,0,217,0,251,0,219,0,49,0,0,0,88,0,0,0,13,0,19,0,58,0,0,0,225,0,193,0,0,0,174,0,120,0,0,0,0,0,199,0,87,0,135,0,105,0,44,0,217,0,34,0,171,0,75,0,159,0,154,0,255,0,94,0,73,0,5,0,63,0,55,0,0,0,30,0,16,0,67,0,236,0,188,0,196,0,25,0,237,0,101,0,0,0,155,0,79,0,59,0,70,0,63,0,33,0,145,0,57,0,200,0,80,0,0,0,0,0,130,0,0,0,0,0,155,0,142,0,239,0,2,0,0,0,170,0,0,0,197,0,94,0,188,0,28,0,0,0,244,0,200,0,0,0,226,0,59,0,22,0,0,0,216,0,39,0,13,0,0,0,174,0,141,0,84,0,27,0,1,0,51,0,69,0,124,0,224,0,93,0,123,0,0,0,0,0,141,0,9,0,25,0,18,0,4,0,58,0,7,0,155,0,127,0,153,0,62,0,0,0,0,0,0,0,50,0,0,0,0,0,239,0,182,0,0,0,233,0,216,0,15,0,25,0,87,0,241,0,24,0,173,0,246,0,60,0,208,0,204,0,196,0,52,0,22,0,225,0,23,0,225,0,43,0,38,0,120,0,0,0,59,0,68,0,0,0,68,0,195,0,50,0,0,0,41,0,159,0,181,0,100,0,237,0,133,0,200,0,33,0,248,0,101,0,247,0,0,0,30,0,161,0,2,0,123,0,228,0,59,0,0,0,0,0,168,0,83,0,80,0,223,0,0,0,103,0,126,0,0,0,45,0,215,0,123,0,81,0,19,0,217,0,255,0,84,0,26,0,21,0,118,0,42,0,112,0,106,0,199,0,224,0,246,0,175,0,250,0,186,0,201,0,210,0,127,0,0,0,83,0,43,0,0,0,41,0,1,0,52,0,130,0,32,0,0,0,166,0,9,0,57,0,168,0,0,0,91,0,76,0,189,0,0,0,170,0,0,0,230,0,0,0,123,0,178,0,75,0,0,0,187,0,27,0,209,0,28,0,84,0,145,0,0,0,0,0,112,0,65,0,0,0,195,0,170,0,89,0,211,0,0,0,41,0,77,0,140,0,170,0,142,0,48,0,106,0,0,0,6,0,57,0,68,0,9,0,0,0,216,0,0,0,248,0,0,0,51,0,188,0,204,0,153,0,250,0,217,0,0,0,0,0,233,0,242,0,43,0,250,0,0,0,0,0,117,0,177,0,17,0,47,0,62,0,8,0,192,0,225,0,36,0,175,0,230,0,40,0,0,0,186,0,0,0,18,0,0,0,0,0,128,0,174,0,152,0,41,0,229,0,82,0,230,0,0,0,0,0,140,0,0,0,0,0,17,0,4,0,0,0,212,0,239,0,186,0,51,0,4,0,137,0,8,0,94,0,4,0,105,0,163,0,222,0,0,0,0,0,195,0,93,0,162,0,0,0,233,0,74,0,101,0,137,0,220,0,225,0,10,0,109,0,94,0,4,0,134,0,234,0,179,0,12,0,192,0,106,0,7,0,166,0,195,0,0,0,233,0,0,0,108,0,3,0,12,0,0,0,216,0,250,0,155,0,1,0,0,0,96,0,0,0,244,0,113,0,166,0,77,0,106,0,237,0,230,0,7,0,233,0,186,0,54,0,159,0,37,0,23,0,0,0,48,0,121,0,157,0,0,0,169,0,116,0,223,0,255,0,0,0,222,0,130,0,20,0,179,0,13,0,239,0,180,0,0,0,12,0,0,0,176,0,29,0,15,0,0,0,184,0,0,0,0,0,0,0,0,0,54,0,0,0,203,0,71,0,80,0,168,0,53,0,35,0,149,0,157,0,0,0,0,0,242,0,80,0,203,0,23,0,0,0,176,0,208,0,75,0,125,0,0,0,0,0,55,0,207,0,0,0,164,0,160,0,32,0,0,0,103,0,165,0,194,0,0,0,0,0,0,0,100,0,158,0,85,0,228,0,100,0,0,0,0,0,0,0,0,0,27,0,185,0,170,0,122,0,0,0,0,0,93,0,149,0,47,0,210,0,70,0,93,0,0,0,127,0,187,0,0,0,17,0,0,0,161,0,196,0,185,0,0,0,72,0,0,0,136,0,87,0,114,0,120,0,254,0,208,0,0,0,79,0,74,0,128,0,235,0,105,0,44,0,120,0,56,0,23,0,127,0,1,0,0,0,14,0,94,0,0,0,138,0,168,0,216,0,196,0,0,0,247,0,150,0,100,0,217,0,222,0,30,0,195,0,87,0,9,0,0,0,0,0,0,0,0,0,16,0,15,0,0,0,61,0,0,0,220,0,205,0,74,0,0,0,0,0,139,0,245,0,38,0,219,0,110,0,80,0,62,0,81,0,76,0,56,0,0,0,166,0,50,0,0,0,90,0,0,0,0,0,189,0,0,0,81,0,0,0,0,0,135,0,125,0,0,0,21,0,0,0,119,0,247,0,118,0,119,0,101,0,0,0,65,0,56,0,0,0,156,0,189,0,166,0,148,0,44,0,204,0,156,0,95,0,68,0,137,0,0,0,199,0,0,0,127,0,41,0,213,0,58,0,114,0,36,0,64,0,42,0,225,0,0,0,224,0,0,0,106,0,102,0,0,0,0,0,248,0,20,0,0,0,0,0,0,0,198,0,6,0,0,0,82,0,1,0,22,0,0,0,75,0,148,0,13,0,101,0,225,0,212,0,180,0,151,0,125,0,146,0,0,0,220,0,153,0,245,0,131,0,188,0,84,0,23,0,142,0,102,0,126,0,85,0,162,0,113,0,231,0,0,0,0,0,0,0,179,0,188,0,0,0,215,0,169,0,51,0,97,0,173,0,134,0,0,0,0,0,188,0,254,0,33,0,253,0,67,0,226,0,152,0,237,0,102,0,0,0,105,0,24,0,173,0,60,0,221,0,32,0,96,0,207,0,2,0,71,0,61,0,166,0,0,0,0,0,2,0,0,0,0,0,198,0,143,0,150,0,142,0,0,0,197,0,234,0,246,0,60,0,249,0,110,0,208,0,204,0,187,0,39,0,0,0,215,0,10,0,1,0,243,0,0,0,14,0,50,0,0,0,226,0,253,0,0,0,164,0,171,0,0,0,50,0,216,0,221,0,9,0,0,0,65,0,144,0,76,0,97,0,187,0,92,0,145,0,64,0,244,0,227,0,0,0,141,0,28,0,0,0,0,0,255,0,189,0,232,0,19,0,0,0,0,0,49,0,142,0,44,0,109,0,64,0,0,0,235,0,0,0,225,0,22,0,238,0,0,0,222,0,46,0,105,0,0,0,162,0,114,0,209,0,209,0,38,0,187,0,0,0,189,0,0,0,0,0,237,0,0,0,0,0,0,0,162,0,241,0,0,0,9,0,0,0,0,0,109,0,0,0,11,0,98,0,171,0,210,0,0,0,20,0,153,0,0,0,145,0,160,0,90,0,0,0,81,0,0,0,75,0,160,0,100,0,0,0,186,0,162,0,38,0,0,0,32,0,87,0,146,0,170,0,0,0,197,0,182,0,0,0,87,0,0,0,166,0,0,0,133,0,0,0,118,0,79,0,206,0,247,0,94,0,206,0,21,0,3,0,68,0,141,0,164,0,184,0,140,0,145,0,4,0,0,0,51,0,31,0,28,0,247,0,0,0,0,0,226,0,93,0,0,0,36,0,0,0,104,0,0,0,57,0,240,0,79,0,0,0,158,0,218,0,167,0,0,0,102,0,47,0,185,0,215,0,221,0,0,0,255,0,231,0,0,0,112,0,166,0,20,0,3,0,209,0,164,0,199,0,0,0,136,0,0,0);
signal scenario_full  : scenario_type := (218,31,187,31,141,31,163,31,121,31,86,31,196,31,81,31,81,30,81,29,6,31,73,31,249,31,71,31,25,31,223,31,145,31,178,31,129,31,200,31,170,31,7,31,7,30,77,31,22,31,156,31,144,31,175,31,175,30,35,31,97,31,180,31,94,31,103,31,245,31,245,30,2,31,246,31,150,31,212,31,212,30,185,31,152,31,12,31,54,31,54,30,57,31,166,31,51,31,51,30,41,31,215,31,80,31,1,31,6,31,21,31,233,31,251,31,211,31,211,30,26,31,19,31,19,30,207,31,207,30,207,29,246,31,16,31,36,31,99,31,114,31,118,31,185,31,217,31,251,31,219,31,49,31,49,30,88,31,88,30,13,31,19,31,58,31,58,30,225,31,193,31,193,30,174,31,120,31,120,30,120,29,199,31,87,31,135,31,105,31,44,31,217,31,34,31,171,31,75,31,159,31,154,31,255,31,94,31,73,31,5,31,63,31,55,31,55,30,30,31,16,31,67,31,236,31,188,31,196,31,25,31,237,31,101,31,101,30,155,31,79,31,59,31,70,31,63,31,33,31,145,31,57,31,200,31,80,31,80,30,80,29,130,31,130,30,130,29,155,31,142,31,239,31,2,31,2,30,170,31,170,30,197,31,94,31,188,31,28,31,28,30,244,31,200,31,200,30,226,31,59,31,22,31,22,30,216,31,39,31,13,31,13,30,174,31,141,31,84,31,27,31,1,31,51,31,69,31,124,31,224,31,93,31,123,31,123,30,123,29,141,31,9,31,25,31,18,31,4,31,58,31,7,31,155,31,127,31,153,31,62,31,62,30,62,29,62,28,50,31,50,30,50,29,239,31,182,31,182,30,233,31,216,31,15,31,25,31,87,31,241,31,24,31,173,31,246,31,60,31,208,31,204,31,196,31,52,31,22,31,225,31,23,31,225,31,43,31,38,31,120,31,120,30,59,31,68,31,68,30,68,31,195,31,50,31,50,30,41,31,159,31,181,31,100,31,237,31,133,31,200,31,33,31,248,31,101,31,247,31,247,30,30,31,161,31,2,31,123,31,228,31,59,31,59,30,59,29,168,31,83,31,80,31,223,31,223,30,103,31,126,31,126,30,45,31,215,31,123,31,81,31,19,31,217,31,255,31,84,31,26,31,21,31,118,31,42,31,112,31,106,31,199,31,224,31,246,31,175,31,250,31,186,31,201,31,210,31,127,31,127,30,83,31,43,31,43,30,41,31,1,31,52,31,130,31,32,31,32,30,166,31,9,31,57,31,168,31,168,30,91,31,76,31,189,31,189,30,170,31,170,30,230,31,230,30,123,31,178,31,75,31,75,30,187,31,27,31,209,31,28,31,84,31,145,31,145,30,145,29,112,31,65,31,65,30,195,31,170,31,89,31,211,31,211,30,41,31,77,31,140,31,170,31,142,31,48,31,106,31,106,30,6,31,57,31,68,31,9,31,9,30,216,31,216,30,248,31,248,30,51,31,188,31,204,31,153,31,250,31,217,31,217,30,217,29,233,31,242,31,43,31,250,31,250,30,250,29,117,31,177,31,17,31,47,31,62,31,8,31,192,31,225,31,36,31,175,31,230,31,40,31,40,30,186,31,186,30,18,31,18,30,18,29,128,31,174,31,152,31,41,31,229,31,82,31,230,31,230,30,230,29,140,31,140,30,140,29,17,31,4,31,4,30,212,31,239,31,186,31,51,31,4,31,137,31,8,31,94,31,4,31,105,31,163,31,222,31,222,30,222,29,195,31,93,31,162,31,162,30,233,31,74,31,101,31,137,31,220,31,225,31,10,31,109,31,94,31,4,31,134,31,234,31,179,31,12,31,192,31,106,31,7,31,166,31,195,31,195,30,233,31,233,30,108,31,3,31,12,31,12,30,216,31,250,31,155,31,1,31,1,30,96,31,96,30,244,31,113,31,166,31,77,31,106,31,237,31,230,31,7,31,233,31,186,31,54,31,159,31,37,31,23,31,23,30,48,31,121,31,157,31,157,30,169,31,116,31,223,31,255,31,255,30,222,31,130,31,20,31,179,31,13,31,239,31,180,31,180,30,12,31,12,30,176,31,29,31,15,31,15,30,184,31,184,30,184,29,184,28,184,27,54,31,54,30,203,31,71,31,80,31,168,31,53,31,35,31,149,31,157,31,157,30,157,29,242,31,80,31,203,31,23,31,23,30,176,31,208,31,75,31,125,31,125,30,125,29,55,31,207,31,207,30,164,31,160,31,32,31,32,30,103,31,165,31,194,31,194,30,194,29,194,28,100,31,158,31,85,31,228,31,100,31,100,30,100,29,100,28,100,27,27,31,185,31,170,31,122,31,122,30,122,29,93,31,149,31,47,31,210,31,70,31,93,31,93,30,127,31,187,31,187,30,17,31,17,30,161,31,196,31,185,31,185,30,72,31,72,30,136,31,87,31,114,31,120,31,254,31,208,31,208,30,79,31,74,31,128,31,235,31,105,31,44,31,120,31,56,31,23,31,127,31,1,31,1,30,14,31,94,31,94,30,138,31,168,31,216,31,196,31,196,30,247,31,150,31,100,31,217,31,222,31,30,31,195,31,87,31,9,31,9,30,9,29,9,28,9,27,16,31,15,31,15,30,61,31,61,30,220,31,205,31,74,31,74,30,74,29,139,31,245,31,38,31,219,31,110,31,80,31,62,31,81,31,76,31,56,31,56,30,166,31,50,31,50,30,90,31,90,30,90,29,189,31,189,30,81,31,81,30,81,29,135,31,125,31,125,30,21,31,21,30,119,31,247,31,118,31,119,31,101,31,101,30,65,31,56,31,56,30,156,31,189,31,166,31,148,31,44,31,204,31,156,31,95,31,68,31,137,31,137,30,199,31,199,30,127,31,41,31,213,31,58,31,114,31,36,31,64,31,42,31,225,31,225,30,224,31,224,30,106,31,102,31,102,30,102,29,248,31,20,31,20,30,20,29,20,28,198,31,6,31,6,30,82,31,1,31,22,31,22,30,75,31,148,31,13,31,101,31,225,31,212,31,180,31,151,31,125,31,146,31,146,30,220,31,153,31,245,31,131,31,188,31,84,31,23,31,142,31,102,31,126,31,85,31,162,31,113,31,231,31,231,30,231,29,231,28,179,31,188,31,188,30,215,31,169,31,51,31,97,31,173,31,134,31,134,30,134,29,188,31,254,31,33,31,253,31,67,31,226,31,152,31,237,31,102,31,102,30,105,31,24,31,173,31,60,31,221,31,32,31,96,31,207,31,2,31,71,31,61,31,166,31,166,30,166,29,2,31,2,30,2,29,198,31,143,31,150,31,142,31,142,30,197,31,234,31,246,31,60,31,249,31,110,31,208,31,204,31,187,31,39,31,39,30,215,31,10,31,1,31,243,31,243,30,14,31,50,31,50,30,226,31,253,31,253,30,164,31,171,31,171,30,50,31,216,31,221,31,9,31,9,30,65,31,144,31,76,31,97,31,187,31,92,31,145,31,64,31,244,31,227,31,227,30,141,31,28,31,28,30,28,29,255,31,189,31,232,31,19,31,19,30,19,29,49,31,142,31,44,31,109,31,64,31,64,30,235,31,235,30,225,31,22,31,238,31,238,30,222,31,46,31,105,31,105,30,162,31,114,31,209,31,209,31,38,31,187,31,187,30,189,31,189,30,189,29,237,31,237,30,237,29,237,28,162,31,241,31,241,30,9,31,9,30,9,29,109,31,109,30,11,31,98,31,171,31,210,31,210,30,20,31,153,31,153,30,145,31,160,31,90,31,90,30,81,31,81,30,75,31,160,31,100,31,100,30,186,31,162,31,38,31,38,30,32,31,87,31,146,31,170,31,170,30,197,31,182,31,182,30,87,31,87,30,166,31,166,30,133,31,133,30,118,31,79,31,206,31,247,31,94,31,206,31,21,31,3,31,68,31,141,31,164,31,184,31,140,31,145,31,4,31,4,30,51,31,31,31,28,31,247,31,247,30,247,29,226,31,93,31,93,30,36,31,36,30,104,31,104,30,57,31,240,31,79,31,79,30,158,31,218,31,167,31,167,30,102,31,47,31,185,31,215,31,221,31,221,30,255,31,231,31,231,30,112,31,166,31,20,31,3,31,209,31,164,31,199,31,199,30,136,31,136,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
