-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_835 is
end project_tb_835;

architecture project_tb_arch_835 of project_tb_835 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 579;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (178,0,0,0,235,0,236,0,0,0,126,0,142,0,22,0,36,0,0,0,226,0,177,0,94,0,237,0,0,0,41,0,207,0,25,0,214,0,159,0,0,0,46,0,57,0,111,0,9,0,0,0,233,0,25,0,0,0,215,0,0,0,174,0,69,0,138,0,175,0,0,0,151,0,0,0,3,0,49,0,194,0,202,0,11,0,0,0,125,0,61,0,0,0,0,0,2,0,121,0,80,0,0,0,62,0,42,0,110,0,48,0,120,0,67,0,17,0,230,0,249,0,155,0,136,0,0,0,0,0,36,0,150,0,24,0,0,0,202,0,92,0,219,0,144,0,0,0,66,0,147,0,122,0,0,0,239,0,122,0,205,0,0,0,82,0,79,0,106,0,38,0,71,0,26,0,233,0,136,0,252,0,0,0,50,0,6,0,0,0,231,0,158,0,226,0,231,0,39,0,119,0,63,0,20,0,108,0,107,0,39,0,46,0,0,0,162,0,6,0,211,0,95,0,131,0,196,0,253,0,93,0,149,0,72,0,20,0,223,0,227,0,51,0,166,0,94,0,120,0,158,0,67,0,11,0,2,0,26,0,153,0,12,0,0,0,104,0,0,0,4,0,78,0,202,0,0,0,240,0,169,0,0,0,0,0,15,0,81,0,22,0,116,0,22,0,51,0,231,0,0,0,98,0,248,0,107,0,1,0,214,0,0,0,101,0,96,0,154,0,151,0,144,0,251,0,114,0,108,0,194,0,182,0,240,0,99,0,147,0,251,0,174,0,242,0,0,0,52,0,159,0,149,0,0,0,240,0,113,0,116,0,217,0,221,0,20,0,0,0,0,0,35,0,0,0,40,0,220,0,149,0,188,0,184,0,21,0,19,0,0,0,0,0,171,0,0,0,97,0,82,0,30,0,244,0,59,0,225,0,153,0,89,0,234,0,115,0,0,0,0,0,0,0,229,0,147,0,171,0,0,0,69,0,86,0,196,0,70,0,194,0,187,0,165,0,66,0,64,0,76,0,237,0,218,0,0,0,63,0,78,0,134,0,0,0,218,0,248,0,60,0,0,0,77,0,234,0,8,0,18,0,253,0,252,0,0,0,204,0,201,0,105,0,114,0,0,0,144,0,172,0,139,0,219,0,0,0,0,0,128,0,0,0,156,0,0,0,110,0,13,0,114,0,94,0,109,0,0,0,146,0,228,0,248,0,1,0,0,0,61,0,58,0,61,0,9,0,0,0,23,0,0,0,36,0,0,0,6,0,223,0,0,0,109,0,247,0,212,0,129,0,122,0,99,0,73,0,127,0,182,0,0,0,42,0,0,0,100,0,181,0,203,0,218,0,196,0,170,0,221,0,72,0,7,0,114,0,20,0,155,0,32,0,45,0,0,0,217,0,22,0,0,0,91,0,175,0,0,0,74,0,22,0,78,0,70,0,169,0,241,0,0,0,215,0,0,0,76,0,109,0,237,0,78,0,138,0,95,0,223,0,188,0,129,0,95,0,167,0,131,0,0,0,63,0,155,0,0,0,0,0,0,0,146,0,55,0,239,0,94,0,69,0,133,0,0,0,60,0,245,0,151,0,0,0,234,0,0,0,74,0,14,0,105,0,148,0,219,0,154,0,97,0,236,0,220,0,94,0,191,0,0,0,0,0,214,0,0,0,145,0,0,0,100,0,248,0,199,0,155,0,133,0,58,0,85,0,27,0,231,0,2,0,217,0,43,0,39,0,163,0,170,0,0,0,0,0,100,0,148,0,42,0,0,0,0,0,204,0,37,0,235,0,0,0,188,0,0,0,22,0,0,0,0,0,0,0,129,0,10,0,0,0,146,0,225,0,136,0,103,0,0,0,39,0,45,0,0,0,0,0,150,0,0,0,240,0,0,0,37,0,175,0,0,0,206,0,203,0,118,0,214,0,148,0,183,0,44,0,214,0,64,0,44,0,0,0,146,0,155,0,55,0,186,0,0,0,0,0,0,0,73,0,18,0,0,0,88,0,151,0,156,0,84,0,68,0,0,0,98,0,78,0,64,0,104,0,0,0,0,0,179,0,237,0,0,0,99,0,163,0,91,0,38,0,5,0,18,0,0,0,0,0,0,0,46,0,136,0,153,0,107,0,50,0,115,0,97,0,31,0,155,0,40,0,45,0,162,0,0,0,0,0,64,0,0,0,99,0,0,0,30,0,76,0,70,0,37,0,167,0,253,0,55,0,0,0,146,0,29,0,67,0,0,0,93,0,201,0,243,0,184,0,0,0,0,0,128,0,0,0,3,0,247,0,158,0,0,0,228,0,89,0,181,0,239,0,168,0,0,0,199,0,207,0,149,0,0,0,0,0,113,0,203,0,235,0,0,0,111,0,85,0,13,0,230,0,56,0,199,0,5,0,105,0,7,0,120,0,9,0,15,0,208,0,205,0,0,0,42,0,15,0,29,0,238,0,0,0,68,0,177,0,166,0,0,0,214,0,31,0,0,0,157,0,0,0,0,0,181,0,66,0,0,0,199,0,97,0,248,0,198,0,156,0,0,0,197,0,178,0,219,0,0,0,45,0,32,0,252,0,0,0,94,0,86,0,204,0,70,0,89,0,26,0,156,0);
signal scenario_full  : scenario_type := (178,31,178,30,235,31,236,31,236,30,126,31,142,31,22,31,36,31,36,30,226,31,177,31,94,31,237,31,237,30,41,31,207,31,25,31,214,31,159,31,159,30,46,31,57,31,111,31,9,31,9,30,233,31,25,31,25,30,215,31,215,30,174,31,69,31,138,31,175,31,175,30,151,31,151,30,3,31,49,31,194,31,202,31,11,31,11,30,125,31,61,31,61,30,61,29,2,31,121,31,80,31,80,30,62,31,42,31,110,31,48,31,120,31,67,31,17,31,230,31,249,31,155,31,136,31,136,30,136,29,36,31,150,31,24,31,24,30,202,31,92,31,219,31,144,31,144,30,66,31,147,31,122,31,122,30,239,31,122,31,205,31,205,30,82,31,79,31,106,31,38,31,71,31,26,31,233,31,136,31,252,31,252,30,50,31,6,31,6,30,231,31,158,31,226,31,231,31,39,31,119,31,63,31,20,31,108,31,107,31,39,31,46,31,46,30,162,31,6,31,211,31,95,31,131,31,196,31,253,31,93,31,149,31,72,31,20,31,223,31,227,31,51,31,166,31,94,31,120,31,158,31,67,31,11,31,2,31,26,31,153,31,12,31,12,30,104,31,104,30,4,31,78,31,202,31,202,30,240,31,169,31,169,30,169,29,15,31,81,31,22,31,116,31,22,31,51,31,231,31,231,30,98,31,248,31,107,31,1,31,214,31,214,30,101,31,96,31,154,31,151,31,144,31,251,31,114,31,108,31,194,31,182,31,240,31,99,31,147,31,251,31,174,31,242,31,242,30,52,31,159,31,149,31,149,30,240,31,113,31,116,31,217,31,221,31,20,31,20,30,20,29,35,31,35,30,40,31,220,31,149,31,188,31,184,31,21,31,19,31,19,30,19,29,171,31,171,30,97,31,82,31,30,31,244,31,59,31,225,31,153,31,89,31,234,31,115,31,115,30,115,29,115,28,229,31,147,31,171,31,171,30,69,31,86,31,196,31,70,31,194,31,187,31,165,31,66,31,64,31,76,31,237,31,218,31,218,30,63,31,78,31,134,31,134,30,218,31,248,31,60,31,60,30,77,31,234,31,8,31,18,31,253,31,252,31,252,30,204,31,201,31,105,31,114,31,114,30,144,31,172,31,139,31,219,31,219,30,219,29,128,31,128,30,156,31,156,30,110,31,13,31,114,31,94,31,109,31,109,30,146,31,228,31,248,31,1,31,1,30,61,31,58,31,61,31,9,31,9,30,23,31,23,30,36,31,36,30,6,31,223,31,223,30,109,31,247,31,212,31,129,31,122,31,99,31,73,31,127,31,182,31,182,30,42,31,42,30,100,31,181,31,203,31,218,31,196,31,170,31,221,31,72,31,7,31,114,31,20,31,155,31,32,31,45,31,45,30,217,31,22,31,22,30,91,31,175,31,175,30,74,31,22,31,78,31,70,31,169,31,241,31,241,30,215,31,215,30,76,31,109,31,237,31,78,31,138,31,95,31,223,31,188,31,129,31,95,31,167,31,131,31,131,30,63,31,155,31,155,30,155,29,155,28,146,31,55,31,239,31,94,31,69,31,133,31,133,30,60,31,245,31,151,31,151,30,234,31,234,30,74,31,14,31,105,31,148,31,219,31,154,31,97,31,236,31,220,31,94,31,191,31,191,30,191,29,214,31,214,30,145,31,145,30,100,31,248,31,199,31,155,31,133,31,58,31,85,31,27,31,231,31,2,31,217,31,43,31,39,31,163,31,170,31,170,30,170,29,100,31,148,31,42,31,42,30,42,29,204,31,37,31,235,31,235,30,188,31,188,30,22,31,22,30,22,29,22,28,129,31,10,31,10,30,146,31,225,31,136,31,103,31,103,30,39,31,45,31,45,30,45,29,150,31,150,30,240,31,240,30,37,31,175,31,175,30,206,31,203,31,118,31,214,31,148,31,183,31,44,31,214,31,64,31,44,31,44,30,146,31,155,31,55,31,186,31,186,30,186,29,186,28,73,31,18,31,18,30,88,31,151,31,156,31,84,31,68,31,68,30,98,31,78,31,64,31,104,31,104,30,104,29,179,31,237,31,237,30,99,31,163,31,91,31,38,31,5,31,18,31,18,30,18,29,18,28,46,31,136,31,153,31,107,31,50,31,115,31,97,31,31,31,155,31,40,31,45,31,162,31,162,30,162,29,64,31,64,30,99,31,99,30,30,31,76,31,70,31,37,31,167,31,253,31,55,31,55,30,146,31,29,31,67,31,67,30,93,31,201,31,243,31,184,31,184,30,184,29,128,31,128,30,3,31,247,31,158,31,158,30,228,31,89,31,181,31,239,31,168,31,168,30,199,31,207,31,149,31,149,30,149,29,113,31,203,31,235,31,235,30,111,31,85,31,13,31,230,31,56,31,199,31,5,31,105,31,7,31,120,31,9,31,15,31,208,31,205,31,205,30,42,31,15,31,29,31,238,31,238,30,68,31,177,31,166,31,166,30,214,31,31,31,31,30,157,31,157,30,157,29,181,31,66,31,66,30,199,31,97,31,248,31,198,31,156,31,156,30,197,31,178,31,219,31,219,30,45,31,32,31,252,31,252,30,94,31,86,31,204,31,70,31,89,31,26,31,156,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
