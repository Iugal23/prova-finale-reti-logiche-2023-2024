-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_604 is
end project_tb_604;

architecture project_tb_arch_604 of project_tb_604 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 342;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (95,0,203,0,114,0,0,0,232,0,121,0,54,0,0,0,34,0,120,0,1,0,29,0,0,0,0,0,225,0,240,0,49,0,250,0,253,0,134,0,173,0,46,0,95,0,124,0,209,0,0,0,252,0,224,0,115,0,0,0,214,0,147,0,40,0,0,0,204,0,181,0,0,0,83,0,0,0,214,0,83,0,0,0,75,0,231,0,129,0,174,0,105,0,0,0,0,0,228,0,0,0,30,0,5,0,29,0,238,0,88,0,227,0,166,0,155,0,226,0,189,0,188,0,109,0,108,0,143,0,0,0,135,0,251,0,85,0,82,0,91,0,138,0,162,0,238,0,38,0,87,0,219,0,49,0,32,0,175,0,0,0,49,0,109,0,165,0,143,0,100,0,139,0,40,0,0,0,0,0,0,0,0,0,0,0,246,0,0,0,21,0,144,0,73,0,0,0,229,0,129,0,181,0,49,0,0,0,0,0,42,0,255,0,252,0,42,0,45,0,135,0,0,0,253,0,0,0,226,0,130,0,163,0,35,0,28,0,17,0,51,0,205,0,0,0,173,0,235,0,211,0,182,0,172,0,0,0,236,0,152,0,93,0,93,0,0,0,96,0,0,0,128,0,194,0,0,0,134,0,131,0,124,0,196,0,53,0,189,0,125,0,81,0,87,0,212,0,191,0,70,0,89,0,203,0,0,0,104,0,0,0,153,0,47,0,131,0,170,0,54,0,0,0,229,0,226,0,209,0,236,0,249,0,42,0,143,0,0,0,102,0,39,0,34,0,235,0,207,0,0,0,0,0,0,0,229,0,187,0,0,0,111,0,25,0,148,0,80,0,154,0,20,0,147,0,51,0,44,0,238,0,18,0,146,0,73,0,220,0,20,0,0,0,94,0,86,0,161,0,175,0,0,0,131,0,79,0,0,0,214,0,249,0,0,0,10,0,200,0,0,0,126,0,0,0,0,0,0,0,188,0,162,0,30,0,210,0,216,0,115,0,208,0,26,0,184,0,166,0,0,0,250,0,204,0,0,0,244,0,0,0,0,0,0,0,133,0,64,0,0,0,49,0,0,0,99,0,212,0,137,0,188,0,246,0,79,0,59,0,241,0,9,0,0,0,33,0,0,0,182,0,150,0,192,0,49,0,0,0,185,0,0,0,0,0,142,0,121,0,234,0,84,0,240,0,24,0,153,0,225,0,130,0,182,0,45,0,165,0,223,0,153,0,130,0,76,0,0,0,131,0,161,0,219,0,151,0,221,0,96,0,185,0,0,0,0,0,0,0,164,0,69,0,207,0,43,0,121,0,138,0,101,0,55,0,196,0,172,0,46,0,0,0,185,0,106,0,148,0,48,0,0,0,246,0,222,0,25,0,37,0,40,0,0,0,65,0,65,0,0,0,96,0,209,0,0,0,0,0,0,0,126,0,79,0,155,0,85,0,0,0,0,0,196,0,0,0,236,0,0,0,98,0,78,0,15,0,204,0,84,0,199,0,0,0,125,0,57,0,48,0,0,0,0,0,251,0,0,0,203,0,183,0);
signal scenario_full  : scenario_type := (95,31,203,31,114,31,114,30,232,31,121,31,54,31,54,30,34,31,120,31,1,31,29,31,29,30,29,29,225,31,240,31,49,31,250,31,253,31,134,31,173,31,46,31,95,31,124,31,209,31,209,30,252,31,224,31,115,31,115,30,214,31,147,31,40,31,40,30,204,31,181,31,181,30,83,31,83,30,214,31,83,31,83,30,75,31,231,31,129,31,174,31,105,31,105,30,105,29,228,31,228,30,30,31,5,31,29,31,238,31,88,31,227,31,166,31,155,31,226,31,189,31,188,31,109,31,108,31,143,31,143,30,135,31,251,31,85,31,82,31,91,31,138,31,162,31,238,31,38,31,87,31,219,31,49,31,32,31,175,31,175,30,49,31,109,31,165,31,143,31,100,31,139,31,40,31,40,30,40,29,40,28,40,27,40,26,246,31,246,30,21,31,144,31,73,31,73,30,229,31,129,31,181,31,49,31,49,30,49,29,42,31,255,31,252,31,42,31,45,31,135,31,135,30,253,31,253,30,226,31,130,31,163,31,35,31,28,31,17,31,51,31,205,31,205,30,173,31,235,31,211,31,182,31,172,31,172,30,236,31,152,31,93,31,93,31,93,30,96,31,96,30,128,31,194,31,194,30,134,31,131,31,124,31,196,31,53,31,189,31,125,31,81,31,87,31,212,31,191,31,70,31,89,31,203,31,203,30,104,31,104,30,153,31,47,31,131,31,170,31,54,31,54,30,229,31,226,31,209,31,236,31,249,31,42,31,143,31,143,30,102,31,39,31,34,31,235,31,207,31,207,30,207,29,207,28,229,31,187,31,187,30,111,31,25,31,148,31,80,31,154,31,20,31,147,31,51,31,44,31,238,31,18,31,146,31,73,31,220,31,20,31,20,30,94,31,86,31,161,31,175,31,175,30,131,31,79,31,79,30,214,31,249,31,249,30,10,31,200,31,200,30,126,31,126,30,126,29,126,28,188,31,162,31,30,31,210,31,216,31,115,31,208,31,26,31,184,31,166,31,166,30,250,31,204,31,204,30,244,31,244,30,244,29,244,28,133,31,64,31,64,30,49,31,49,30,99,31,212,31,137,31,188,31,246,31,79,31,59,31,241,31,9,31,9,30,33,31,33,30,182,31,150,31,192,31,49,31,49,30,185,31,185,30,185,29,142,31,121,31,234,31,84,31,240,31,24,31,153,31,225,31,130,31,182,31,45,31,165,31,223,31,153,31,130,31,76,31,76,30,131,31,161,31,219,31,151,31,221,31,96,31,185,31,185,30,185,29,185,28,164,31,69,31,207,31,43,31,121,31,138,31,101,31,55,31,196,31,172,31,46,31,46,30,185,31,106,31,148,31,48,31,48,30,246,31,222,31,25,31,37,31,40,31,40,30,65,31,65,31,65,30,96,31,209,31,209,30,209,29,209,28,126,31,79,31,155,31,85,31,85,30,85,29,196,31,196,30,236,31,236,30,98,31,78,31,15,31,204,31,84,31,199,31,199,30,125,31,57,31,48,31,48,30,48,29,251,31,251,30,203,31,183,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
