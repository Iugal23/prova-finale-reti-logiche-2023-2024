-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_484 is
end project_tb_484;

architecture project_tb_arch_484 of project_tb_484 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 683;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (36,0,14,0,25,0,0,0,0,0,0,0,0,0,0,0,152,0,32,0,0,0,45,0,0,0,77,0,30,0,122,0,0,0,62,0,62,0,5,0,0,0,0,0,0,0,255,0,193,0,60,0,19,0,100,0,146,0,0,0,3,0,79,0,220,0,152,0,87,0,0,0,55,0,0,0,254,0,87,0,107,0,0,0,85,0,191,0,185,0,0,0,173,0,208,0,37,0,176,0,210,0,31,0,5,0,105,0,0,0,0,0,209,0,55,0,36,0,0,0,34,0,67,0,23,0,0,0,0,0,201,0,40,0,0,0,221,0,54,0,216,0,0,0,178,0,98,0,102,0,0,0,0,0,110,0,0,0,103,0,142,0,221,0,0,0,153,0,164,0,190,0,0,0,191,0,0,0,0,0,0,0,13,0,76,0,153,0,0,0,68,0,7,0,46,0,247,0,145,0,0,0,159,0,0,0,0,0,138,0,0,0,244,0,0,0,55,0,179,0,224,0,215,0,0,0,62,0,64,0,167,0,138,0,63,0,113,0,14,0,19,0,95,0,60,0,0,0,214,0,0,0,45,0,0,0,146,0,0,0,66,0,77,0,126,0,102,0,241,0,1,0,198,0,0,0,140,0,243,0,7,0,193,0,0,0,231,0,23,0,0,0,162,0,0,0,9,0,38,0,189,0,173,0,5,0,66,0,128,0,0,0,0,0,16,0,12,0,0,0,241,0,83,0,100,0,0,0,0,0,245,0,247,0,126,0,122,0,199,0,11,0,99,0,59,0,0,0,96,0,122,0,0,0,28,0,243,0,17,0,202,0,227,0,78,0,0,0,168,0,234,0,227,0,72,0,191,0,27,0,0,0,137,0,95,0,130,0,0,0,111,0,0,0,120,0,0,0,0,0,9,0,106,0,0,0,16,0,0,0,201,0,179,0,165,0,111,0,248,0,162,0,0,0,175,0,194,0,75,0,246,0,125,0,152,0,165,0,0,0,175,0,0,0,201,0,0,0,117,0,131,0,201,0,0,0,35,0,44,0,0,0,170,0,248,0,113,0,103,0,128,0,0,0,216,0,230,0,0,0,57,0,19,0,110,0,110,0,74,0,0,0,240,0,40,0,255,0,162,0,163,0,68,0,0,0,0,0,155,0,3,0,141,0,0,0,85,0,58,0,97,0,201,0,214,0,25,0,165,0,203,0,63,0,98,0,164,0,173,0,83,0,13,0,202,0,87,0,166,0,137,0,48,0,144,0,190,0,101,0,0,0,111,0,34,0,29,0,9,0,174,0,115,0,51,0,85,0,44,0,193,0,80,0,64,0,66,0,62,0,202,0,0,0,238,0,68,0,235,0,15,0,228,0,0,0,157,0,17,0,198,0,203,0,249,0,44,0,191,0,230,0,80,0,0,0,110,0,208,0,250,0,56,0,0,0,240,0,0,0,61,0,0,0,61,0,221,0,175,0,218,0,87,0,57,0,136,0,0,0,54,0,44,0,228,0,210,0,251,0,0,0,0,0,176,0,0,0,64,0,47,0,120,0,0,0,18,0,0,0,132,0,13,0,48,0,51,0,71,0,148,0,217,0,172,0,87,0,221,0,0,0,161,0,74,0,4,0,197,0,0,0,1,0,0,0,0,0,164,0,95,0,0,0,0,0,55,0,95,0,65,0,116,0,176,0,52,0,0,0,249,0,53,0,177,0,15,0,243,0,124,0,10,0,0,0,96,0,50,0,191,0,236,0,142,0,188,0,0,0,164,0,95,0,69,0,84,0,86,0,0,0,253,0,154,0,114,0,71,0,121,0,83,0,181,0,88,0,192,0,65,0,17,0,41,0,79,0,106,0,107,0,0,0,47,0,86,0,94,0,46,0,253,0,86,0,34,0,248,0,244,0,0,0,27,0,87,0,58,0,17,0,207,0,0,0,210,0,145,0,86,0,173,0,200,0,145,0,0,0,174,0,123,0,243,0,0,0,50,0,178,0,39,0,0,0,0,0,144,0,209,0,34,0,117,0,0,0,128,0,118,0,104,0,127,0,0,0,0,0,51,0,45,0,105,0,208,0,3,0,101,0,0,0,75,0,0,0,0,0,78,0,148,0,0,0,0,0,46,0,126,0,198,0,121,0,142,0,199,0,90,0,141,0,0,0,26,0,31,0,38,0,0,0,46,0,226,0,93,0,0,0,0,0,184,0,0,0,58,0,244,0,122,0,0,0,64,0,0,0,105,0,0,0,106,0,53,0,70,0,114,0,235,0,0,0,0,0,33,0,32,0,84,0,97,0,0,0,128,0,182,0,150,0,126,0,128,0,214,0,181,0,46,0,44,0,148,0,137,0,0,0,147,0,170,0,0,0,0,0,160,0,0,0,57,0,73,0,108,0,205,0,107,0,0,0,0,0,177,0,0,0,0,0,3,0,103,0,70,0,74,0,191,0,0,0,121,0,0,0,0,0,247,0,0,0,47,0,244,0,178,0,162,0,246,0,0,0,0,0,22,0,64,0,237,0,1,0,0,0,207,0,123,0,205,0,0,0,210,0,146,0,76,0,5,0,15,0,154,0,0,0,130,0,245,0,62,0,108,0,100,0,0,0,49,0,117,0,0,0,7,0,132,0,252,0,192,0,69,0,0,0,230,0,169,0,31,0,48,0,0,0,109,0,183,0,216,0,110,0,233,0,84,0,113,0,32,0,0,0,0,0,0,0,0,0,46,0,105,0,0,0,255,0,238,0,107,0,242,0,0,0,228,0,246,0,240,0,192,0,0,0,226,0,0,0,43,0,183,0,207,0,250,0,55,0,109,0,166,0,0,0,175,0,49,0,149,0,14,0,57,0,110,0,32,0,163,0,173,0,0,0,0,0,207,0,225,0,99,0,0,0,0,0,127,0,119,0,1,0,129,0,69,0,97,0,53,0,11,0,233,0,0,0,107,0,144,0,132,0,106,0,21,0,86,0,41,0,173,0,56,0,128,0,51,0,9,0,139,0,16,0,148,0,208,0,137,0,126,0,249,0,150,0,0,0,114,0,163,0,188,0,1,0,0,0,97,0,162,0,0,0,79,0,177,0);
signal scenario_full  : scenario_type := (36,31,14,31,25,31,25,30,25,29,25,28,25,27,25,26,152,31,32,31,32,30,45,31,45,30,77,31,30,31,122,31,122,30,62,31,62,31,5,31,5,30,5,29,5,28,255,31,193,31,60,31,19,31,100,31,146,31,146,30,3,31,79,31,220,31,152,31,87,31,87,30,55,31,55,30,254,31,87,31,107,31,107,30,85,31,191,31,185,31,185,30,173,31,208,31,37,31,176,31,210,31,31,31,5,31,105,31,105,30,105,29,209,31,55,31,36,31,36,30,34,31,67,31,23,31,23,30,23,29,201,31,40,31,40,30,221,31,54,31,216,31,216,30,178,31,98,31,102,31,102,30,102,29,110,31,110,30,103,31,142,31,221,31,221,30,153,31,164,31,190,31,190,30,191,31,191,30,191,29,191,28,13,31,76,31,153,31,153,30,68,31,7,31,46,31,247,31,145,31,145,30,159,31,159,30,159,29,138,31,138,30,244,31,244,30,55,31,179,31,224,31,215,31,215,30,62,31,64,31,167,31,138,31,63,31,113,31,14,31,19,31,95,31,60,31,60,30,214,31,214,30,45,31,45,30,146,31,146,30,66,31,77,31,126,31,102,31,241,31,1,31,198,31,198,30,140,31,243,31,7,31,193,31,193,30,231,31,23,31,23,30,162,31,162,30,9,31,38,31,189,31,173,31,5,31,66,31,128,31,128,30,128,29,16,31,12,31,12,30,241,31,83,31,100,31,100,30,100,29,245,31,247,31,126,31,122,31,199,31,11,31,99,31,59,31,59,30,96,31,122,31,122,30,28,31,243,31,17,31,202,31,227,31,78,31,78,30,168,31,234,31,227,31,72,31,191,31,27,31,27,30,137,31,95,31,130,31,130,30,111,31,111,30,120,31,120,30,120,29,9,31,106,31,106,30,16,31,16,30,201,31,179,31,165,31,111,31,248,31,162,31,162,30,175,31,194,31,75,31,246,31,125,31,152,31,165,31,165,30,175,31,175,30,201,31,201,30,117,31,131,31,201,31,201,30,35,31,44,31,44,30,170,31,248,31,113,31,103,31,128,31,128,30,216,31,230,31,230,30,57,31,19,31,110,31,110,31,74,31,74,30,240,31,40,31,255,31,162,31,163,31,68,31,68,30,68,29,155,31,3,31,141,31,141,30,85,31,58,31,97,31,201,31,214,31,25,31,165,31,203,31,63,31,98,31,164,31,173,31,83,31,13,31,202,31,87,31,166,31,137,31,48,31,144,31,190,31,101,31,101,30,111,31,34,31,29,31,9,31,174,31,115,31,51,31,85,31,44,31,193,31,80,31,64,31,66,31,62,31,202,31,202,30,238,31,68,31,235,31,15,31,228,31,228,30,157,31,17,31,198,31,203,31,249,31,44,31,191,31,230,31,80,31,80,30,110,31,208,31,250,31,56,31,56,30,240,31,240,30,61,31,61,30,61,31,221,31,175,31,218,31,87,31,57,31,136,31,136,30,54,31,44,31,228,31,210,31,251,31,251,30,251,29,176,31,176,30,64,31,47,31,120,31,120,30,18,31,18,30,132,31,13,31,48,31,51,31,71,31,148,31,217,31,172,31,87,31,221,31,221,30,161,31,74,31,4,31,197,31,197,30,1,31,1,30,1,29,164,31,95,31,95,30,95,29,55,31,95,31,65,31,116,31,176,31,52,31,52,30,249,31,53,31,177,31,15,31,243,31,124,31,10,31,10,30,96,31,50,31,191,31,236,31,142,31,188,31,188,30,164,31,95,31,69,31,84,31,86,31,86,30,253,31,154,31,114,31,71,31,121,31,83,31,181,31,88,31,192,31,65,31,17,31,41,31,79,31,106,31,107,31,107,30,47,31,86,31,94,31,46,31,253,31,86,31,34,31,248,31,244,31,244,30,27,31,87,31,58,31,17,31,207,31,207,30,210,31,145,31,86,31,173,31,200,31,145,31,145,30,174,31,123,31,243,31,243,30,50,31,178,31,39,31,39,30,39,29,144,31,209,31,34,31,117,31,117,30,128,31,118,31,104,31,127,31,127,30,127,29,51,31,45,31,105,31,208,31,3,31,101,31,101,30,75,31,75,30,75,29,78,31,148,31,148,30,148,29,46,31,126,31,198,31,121,31,142,31,199,31,90,31,141,31,141,30,26,31,31,31,38,31,38,30,46,31,226,31,93,31,93,30,93,29,184,31,184,30,58,31,244,31,122,31,122,30,64,31,64,30,105,31,105,30,106,31,53,31,70,31,114,31,235,31,235,30,235,29,33,31,32,31,84,31,97,31,97,30,128,31,182,31,150,31,126,31,128,31,214,31,181,31,46,31,44,31,148,31,137,31,137,30,147,31,170,31,170,30,170,29,160,31,160,30,57,31,73,31,108,31,205,31,107,31,107,30,107,29,177,31,177,30,177,29,3,31,103,31,70,31,74,31,191,31,191,30,121,31,121,30,121,29,247,31,247,30,47,31,244,31,178,31,162,31,246,31,246,30,246,29,22,31,64,31,237,31,1,31,1,30,207,31,123,31,205,31,205,30,210,31,146,31,76,31,5,31,15,31,154,31,154,30,130,31,245,31,62,31,108,31,100,31,100,30,49,31,117,31,117,30,7,31,132,31,252,31,192,31,69,31,69,30,230,31,169,31,31,31,48,31,48,30,109,31,183,31,216,31,110,31,233,31,84,31,113,31,32,31,32,30,32,29,32,28,32,27,46,31,105,31,105,30,255,31,238,31,107,31,242,31,242,30,228,31,246,31,240,31,192,31,192,30,226,31,226,30,43,31,183,31,207,31,250,31,55,31,109,31,166,31,166,30,175,31,49,31,149,31,14,31,57,31,110,31,32,31,163,31,173,31,173,30,173,29,207,31,225,31,99,31,99,30,99,29,127,31,119,31,1,31,129,31,69,31,97,31,53,31,11,31,233,31,233,30,107,31,144,31,132,31,106,31,21,31,86,31,41,31,173,31,56,31,128,31,51,31,9,31,139,31,16,31,148,31,208,31,137,31,126,31,249,31,150,31,150,30,114,31,163,31,188,31,1,31,1,30,97,31,162,31,162,30,79,31,177,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
