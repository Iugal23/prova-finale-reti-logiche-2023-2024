-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_946 is
end project_tb_946;

architecture project_tb_arch_946 of project_tb_946 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 200;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (89,0,0,0,247,0,0,0,0,0,76,0,215,0,158,0,1,0,92,0,169,0,215,0,0,0,92,0,0,0,4,0,152,0,3,0,0,0,0,0,55,0,101,0,181,0,19,0,6,0,222,0,79,0,0,0,0,0,177,0,145,0,212,0,248,0,0,0,146,0,200,0,93,0,0,0,0,0,8,0,0,0,111,0,212,0,246,0,174,0,171,0,6,0,241,0,39,0,186,0,71,0,10,0,74,0,206,0,132,0,9,0,143,0,32,0,35,0,169,0,0,0,48,0,52,0,145,0,72,0,129,0,0,0,88,0,166,0,182,0,92,0,64,0,0,0,162,0,154,0,8,0,0,0,17,0,0,0,83,0,122,0,241,0,123,0,144,0,28,0,50,0,220,0,34,0,135,0,134,0,66,0,82,0,136,0,161,0,33,0,46,0,88,0,48,0,0,0,80,0,152,0,28,0,148,0,64,0,191,0,41,0,243,0,25,0,39,0,210,0,0,0,220,0,0,0,48,0,6,0,23,0,113,0,82,0,63,0,121,0,154,0,0,0,127,0,0,0,0,0,190,0,182,0,24,0,1,0,115,0,149,0,139,0,59,0,249,0,90,0,141,0,0,0,176,0,57,0,151,0,0,0,229,0,127,0,0,0,0,0,242,0,102,0,86,0,37,0,20,0,159,0,0,0,157,0,0,0,13,0,236,0,0,0,64,0,19,0,231,0,0,0,131,0,112,0,181,0,206,0,72,0,37,0,0,0,7,0,203,0,169,0,29,0,119,0,0,0,0,0,128,0,0,0,185,0,51,0,34,0,0,0,107,0,16,0,0,0,0,0,141,0,228,0,191,0,162,0,0,0,178,0,35,0,0,0,51,0,0,0,22,0,122,0,129,0,184,0,169,0);
signal scenario_full  : scenario_type := (89,31,89,30,247,31,247,30,247,29,76,31,215,31,158,31,1,31,92,31,169,31,215,31,215,30,92,31,92,30,4,31,152,31,3,31,3,30,3,29,55,31,101,31,181,31,19,31,6,31,222,31,79,31,79,30,79,29,177,31,145,31,212,31,248,31,248,30,146,31,200,31,93,31,93,30,93,29,8,31,8,30,111,31,212,31,246,31,174,31,171,31,6,31,241,31,39,31,186,31,71,31,10,31,74,31,206,31,132,31,9,31,143,31,32,31,35,31,169,31,169,30,48,31,52,31,145,31,72,31,129,31,129,30,88,31,166,31,182,31,92,31,64,31,64,30,162,31,154,31,8,31,8,30,17,31,17,30,83,31,122,31,241,31,123,31,144,31,28,31,50,31,220,31,34,31,135,31,134,31,66,31,82,31,136,31,161,31,33,31,46,31,88,31,48,31,48,30,80,31,152,31,28,31,148,31,64,31,191,31,41,31,243,31,25,31,39,31,210,31,210,30,220,31,220,30,48,31,6,31,23,31,113,31,82,31,63,31,121,31,154,31,154,30,127,31,127,30,127,29,190,31,182,31,24,31,1,31,115,31,149,31,139,31,59,31,249,31,90,31,141,31,141,30,176,31,57,31,151,31,151,30,229,31,127,31,127,30,127,29,242,31,102,31,86,31,37,31,20,31,159,31,159,30,157,31,157,30,13,31,236,31,236,30,64,31,19,31,231,31,231,30,131,31,112,31,181,31,206,31,72,31,37,31,37,30,7,31,203,31,169,31,29,31,119,31,119,30,119,29,128,31,128,30,185,31,51,31,34,31,34,30,107,31,16,31,16,30,16,29,141,31,228,31,191,31,162,31,162,30,178,31,35,31,35,30,51,31,51,30,22,31,122,31,129,31,184,31,169,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
