-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_331 is
end project_tb_331;

architecture project_tb_arch_331 of project_tb_331 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 206;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (129,0,236,0,0,0,0,0,249,0,0,0,230,0,151,0,24,0,214,0,47,0,148,0,67,0,174,0,253,0,16,0,167,0,61,0,0,0,237,0,0,0,83,0,142,0,95,0,168,0,151,0,208,0,197,0,78,0,16,0,0,0,118,0,0,0,0,0,98,0,223,0,48,0,0,0,161,0,197,0,128,0,0,0,0,0,72,0,225,0,186,0,139,0,207,0,65,0,0,0,27,0,179,0,0,0,190,0,0,0,0,0,0,0,105,0,240,0,41,0,185,0,129,0,47,0,0,0,234,0,93,0,87,0,152,0,6,0,0,0,0,0,84,0,61,0,200,0,138,0,52,0,29,0,116,0,0,0,181,0,197,0,212,0,134,0,0,0,57,0,60,0,124,0,0,0,4,0,0,0,0,0,1,0,253,0,1,0,0,0,43,0,82,0,142,0,36,0,140,0,202,0,0,0,0,0,157,0,122,0,153,0,66,0,36,0,47,0,128,0,0,0,132,0,205,0,43,0,93,0,0,0,206,0,225,0,111,0,52,0,87,0,0,0,133,0,147,0,94,0,217,0,0,0,136,0,244,0,191,0,1,0,223,0,73,0,149,0,0,0,0,0,108,0,46,0,93,0,0,0,147,0,221,0,95,0,103,0,33,0,154,0,0,0,224,0,125,0,230,0,41,0,0,0,0,0,220,0,8,0,234,0,0,0,43,0,93,0,122,0,171,0,55,0,0,0,132,0,0,0,142,0,114,0,77,0,0,0,44,0,0,0,0,0,224,0,2,0,0,0,0,0,0,0,57,0,0,0,0,0,251,0,0,0,70,0,237,0,0,0,152,0,44,0,27,0,0,0,116,0,192,0,218,0,0,0,177,0,252,0,232,0,249,0,156,0,93,0,155,0,0,0,7,0,182,0,98,0,50,0,0,0);
signal scenario_full  : scenario_type := (129,31,236,31,236,30,236,29,249,31,249,30,230,31,151,31,24,31,214,31,47,31,148,31,67,31,174,31,253,31,16,31,167,31,61,31,61,30,237,31,237,30,83,31,142,31,95,31,168,31,151,31,208,31,197,31,78,31,16,31,16,30,118,31,118,30,118,29,98,31,223,31,48,31,48,30,161,31,197,31,128,31,128,30,128,29,72,31,225,31,186,31,139,31,207,31,65,31,65,30,27,31,179,31,179,30,190,31,190,30,190,29,190,28,105,31,240,31,41,31,185,31,129,31,47,31,47,30,234,31,93,31,87,31,152,31,6,31,6,30,6,29,84,31,61,31,200,31,138,31,52,31,29,31,116,31,116,30,181,31,197,31,212,31,134,31,134,30,57,31,60,31,124,31,124,30,4,31,4,30,4,29,1,31,253,31,1,31,1,30,43,31,82,31,142,31,36,31,140,31,202,31,202,30,202,29,157,31,122,31,153,31,66,31,36,31,47,31,128,31,128,30,132,31,205,31,43,31,93,31,93,30,206,31,225,31,111,31,52,31,87,31,87,30,133,31,147,31,94,31,217,31,217,30,136,31,244,31,191,31,1,31,223,31,73,31,149,31,149,30,149,29,108,31,46,31,93,31,93,30,147,31,221,31,95,31,103,31,33,31,154,31,154,30,224,31,125,31,230,31,41,31,41,30,41,29,220,31,8,31,234,31,234,30,43,31,93,31,122,31,171,31,55,31,55,30,132,31,132,30,142,31,114,31,77,31,77,30,44,31,44,30,44,29,224,31,2,31,2,30,2,29,2,28,57,31,57,30,57,29,251,31,251,30,70,31,237,31,237,30,152,31,44,31,27,31,27,30,116,31,192,31,218,31,218,30,177,31,252,31,232,31,249,31,156,31,93,31,155,31,155,30,7,31,182,31,98,31,50,31,50,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
