-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 750;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (218,0,0,0,0,0,0,0,39,0,40,0,221,0,34,0,0,0,151,0,0,0,52,0,60,0,192,0,251,0,147,0,0,0,97,0,189,0,143,0,219,0,185,0,7,0,86,0,226,0,245,0,49,0,161,0,120,0,169,0,0,0,210,0,238,0,192,0,196,0,106,0,0,0,30,0,132,0,220,0,52,0,97,0,244,0,0,0,126,0,174,0,0,0,173,0,33,0,116,0,0,0,0,0,47,0,108,0,97,0,209,0,232,0,0,0,0,0,204,0,36,0,0,0,71,0,205,0,0,0,208,0,71,0,2,0,0,0,0,0,249,0,154,0,132,0,108,0,156,0,189,0,225,0,106,0,66,0,193,0,0,0,179,0,77,0,252,0,120,0,232,0,14,0,16,0,159,0,0,0,117,0,17,0,138,0,155,0,228,0,0,0,143,0,177,0,163,0,145,0,186,0,37,0,110,0,125,0,50,0,107,0,145,0,0,0,137,0,19,0,59,0,190,0,76,0,33,0,92,0,65,0,51,0,0,0,0,0,49,0,53,0,166,0,119,0,113,0,235,0,0,0,2,0,96,0,147,0,0,0,78,0,179,0,247,0,29,0,0,0,0,0,0,0,0,0,0,0,76,0,131,0,123,0,0,0,166,0,188,0,8,0,98,0,0,0,35,0,0,0,156,0,106,0,58,0,148,0,146,0,0,0,54,0,226,0,13,0,231,0,94,0,0,0,210,0,106,0,178,0,0,0,59,0,232,0,107,0,77,0,38,0,60,0,236,0,20,0,128,0,47,0,0,0,188,0,0,0,174,0,182,0,33,0,236,0,254,0,146,0,37,0,187,0,128,0,35,0,0,0,0,0,0,0,85,0,123,0,109,0,0,0,189,0,0,0,152,0,52,0,131,0,242,0,221,0,0,0,0,0,243,0,142,0,136,0,165,0,108,0,70,0,230,0,4,0,147,0,0,0,62,0,13,0,230,0,89,0,110,0,107,0,19,0,253,0,160,0,0,0,21,0,156,0,253,0,21,0,219,0,175,0,144,0,107,0,3,0,145,0,0,0,48,0,95,0,121,0,105,0,0,0,131,0,234,0,247,0,118,0,159,0,250,0,178,0,40,0,174,0,68,0,0,0,254,0,174,0,242,0,106,0,36,0,18,0,177,0,241,0,0,0,187,0,78,0,161,0,0,0,71,0,78,0,0,0,0,0,0,0,138,0,18,0,42,0,209,0,250,0,0,0,109,0,170,0,121,0,56,0,117,0,141,0,51,0,0,0,230,0,0,0,250,0,150,0,0,0,242,0,10,0,252,0,85,0,0,0,192,0,241,0,227,0,93,0,20,0,60,0,49,0,36,0,251,0,113,0,37,0,168,0,77,0,216,0,0,0,55,0,194,0,16,0,130,0,139,0,0,0,227,0,181,0,0,0,221,0,252,0,217,0,179,0,243,0,192,0,14,0,7,0,5,0,146,0,130,0,0,0,80,0,0,0,0,0,75,0,182,0,41,0,0,0,73,0,222,0,140,0,199,0,185,0,168,0,49,0,28,0,204,0,0,0,0,0,142,0,103,0,0,0,38,0,249,0,15,0,238,0,156,0,199,0,1,0,0,0,100,0,237,0,0,0,131,0,34,0,104,0,121,0,250,0,236,0,0,0,183,0,0,0,211,0,49,0,0,0,233,0,218,0,58,0,0,0,204,0,123,0,213,0,253,0,3,0,56,0,59,0,5,0,10,0,82,0,41,0,193,0,0,0,92,0,188,0,0,0,226,0,14,0,39,0,48,0,0,0,210,0,173,0,234,0,0,0,237,0,0,0,197,0,81,0,238,0,240,0,187,0,152,0,152,0,63,0,148,0,153,0,0,0,0,0,78,0,224,0,213,0,0,0,6,0,113,0,218,0,176,0,199,0,0,0,211,0,187,0,73,0,236,0,135,0,250,0,3,0,91,0,47,0,0,0,15,0,36,0,0,0,180,0,153,0,0,0,173,0,106,0,240,0,0,0,163,0,9,0,251,0,120,0,0,0,0,0,235,0,149,0,197,0,5,0,75,0,0,0,0,0,53,0,0,0,223,0,0,0,33,0,167,0,111,0,105,0,159,0,102,0,0,0,0,0,0,0,204,0,0,0,226,0,34,0,131,0,210,0,0,0,0,0,182,0,98,0,0,0,0,0,108,0,218,0,71,0,145,0,208,0,94,0,159,0,0,0,0,0,4,0,0,0,81,0,152,0,228,0,250,0,0,0,161,0,87,0,8,0,0,0,0,0,0,0,226,0,47,0,152,0,169,0,108,0,0,0,0,0,145,0,70,0,0,0,50,0,0,0,0,0,188,0,17,0,93,0,0,0,239,0,254,0,178,0,0,0,195,0,210,0,190,0,157,0,0,0,44,0,0,0,108,0,97,0,42,0,230,0,166,0,5,0,90,0,253,0,162,0,137,0,185,0,186,0,220,0,235,0,219,0,19,0,112,0,195,0,150,0,154,0,0,0,30,0,167,0,247,0,233,0,127,0,8,0,0,0,192,0,122,0,126,0,66,0,135,0,0,0,234,0,65,0,157,0,83,0,208,0,94,0,174,0,172,0,219,0,127,0,196,0,158,0,81,0,80,0,0,0,83,0,51,0,231,0,96,0,0,0,130,0,15,0,245,0,182,0,208,0,196,0,0,0,205,0,129,0,165,0,0,0,175,0,0,0,0,0,0,0,50,0,84,0,159,0,0,0,150,0,156,0,191,0,204,0,143,0,174,0,183,0,49,0,188,0,38,0,0,0,183,0,110,0,214,0,155,0,123,0,176,0,57,0,102,0,219,0,181,0,172,0,208,0,171,0,0,0,6,0,137,0,25,0,0,0,144,0,19,0,27,0,129,0,181,0,52,0,163,0,25,0,0,0,0,0,77,0,255,0,0,0,170,0,23,0,33,0,150,0,38,0,91,0,118,0,211,0,179,0,0,0,226,0,5,0,210,0,0,0,31,0,56,0,0,0,223,0,184,0,245,0,0,0,143,0,103,0,0,0,191,0,87,0,137,0,200,0,201,0,136,0,120,0,215,0,158,0,45,0,214,0,30,0,0,0,0,0,97,0,9,0,129,0,232,0,190,0,89,0,199,0,24,0,22,0,68,0,0,0,190,0,137,0,118,0,18,0,237,0,74,0,173,0,75,0,156,0,120,0,13,0,191,0,104,0,220,0,200,0,176,0,101,0,62,0,223,0,232,0,227,0,0,0,163,0,181,0,0,0,0,0,156,0,139,0,124,0,0,0,86,0,0,0,238,0,0,0,142,0,95,0,212,0,93,0,61,0,0,0,234,0,176,0,131,0,144,0,24,0,107,0,0,0,161,0,107,0,117,0,167,0);
signal scenario_full  : scenario_type := (218,31,218,30,218,29,218,28,39,31,40,31,221,31,34,31,34,30,151,31,151,30,52,31,60,31,192,31,251,31,147,31,147,30,97,31,189,31,143,31,219,31,185,31,7,31,86,31,226,31,245,31,49,31,161,31,120,31,169,31,169,30,210,31,238,31,192,31,196,31,106,31,106,30,30,31,132,31,220,31,52,31,97,31,244,31,244,30,126,31,174,31,174,30,173,31,33,31,116,31,116,30,116,29,47,31,108,31,97,31,209,31,232,31,232,30,232,29,204,31,36,31,36,30,71,31,205,31,205,30,208,31,71,31,2,31,2,30,2,29,249,31,154,31,132,31,108,31,156,31,189,31,225,31,106,31,66,31,193,31,193,30,179,31,77,31,252,31,120,31,232,31,14,31,16,31,159,31,159,30,117,31,17,31,138,31,155,31,228,31,228,30,143,31,177,31,163,31,145,31,186,31,37,31,110,31,125,31,50,31,107,31,145,31,145,30,137,31,19,31,59,31,190,31,76,31,33,31,92,31,65,31,51,31,51,30,51,29,49,31,53,31,166,31,119,31,113,31,235,31,235,30,2,31,96,31,147,31,147,30,78,31,179,31,247,31,29,31,29,30,29,29,29,28,29,27,29,26,76,31,131,31,123,31,123,30,166,31,188,31,8,31,98,31,98,30,35,31,35,30,156,31,106,31,58,31,148,31,146,31,146,30,54,31,226,31,13,31,231,31,94,31,94,30,210,31,106,31,178,31,178,30,59,31,232,31,107,31,77,31,38,31,60,31,236,31,20,31,128,31,47,31,47,30,188,31,188,30,174,31,182,31,33,31,236,31,254,31,146,31,37,31,187,31,128,31,35,31,35,30,35,29,35,28,85,31,123,31,109,31,109,30,189,31,189,30,152,31,52,31,131,31,242,31,221,31,221,30,221,29,243,31,142,31,136,31,165,31,108,31,70,31,230,31,4,31,147,31,147,30,62,31,13,31,230,31,89,31,110,31,107,31,19,31,253,31,160,31,160,30,21,31,156,31,253,31,21,31,219,31,175,31,144,31,107,31,3,31,145,31,145,30,48,31,95,31,121,31,105,31,105,30,131,31,234,31,247,31,118,31,159,31,250,31,178,31,40,31,174,31,68,31,68,30,254,31,174,31,242,31,106,31,36,31,18,31,177,31,241,31,241,30,187,31,78,31,161,31,161,30,71,31,78,31,78,30,78,29,78,28,138,31,18,31,42,31,209,31,250,31,250,30,109,31,170,31,121,31,56,31,117,31,141,31,51,31,51,30,230,31,230,30,250,31,150,31,150,30,242,31,10,31,252,31,85,31,85,30,192,31,241,31,227,31,93,31,20,31,60,31,49,31,36,31,251,31,113,31,37,31,168,31,77,31,216,31,216,30,55,31,194,31,16,31,130,31,139,31,139,30,227,31,181,31,181,30,221,31,252,31,217,31,179,31,243,31,192,31,14,31,7,31,5,31,146,31,130,31,130,30,80,31,80,30,80,29,75,31,182,31,41,31,41,30,73,31,222,31,140,31,199,31,185,31,168,31,49,31,28,31,204,31,204,30,204,29,142,31,103,31,103,30,38,31,249,31,15,31,238,31,156,31,199,31,1,31,1,30,100,31,237,31,237,30,131,31,34,31,104,31,121,31,250,31,236,31,236,30,183,31,183,30,211,31,49,31,49,30,233,31,218,31,58,31,58,30,204,31,123,31,213,31,253,31,3,31,56,31,59,31,5,31,10,31,82,31,41,31,193,31,193,30,92,31,188,31,188,30,226,31,14,31,39,31,48,31,48,30,210,31,173,31,234,31,234,30,237,31,237,30,197,31,81,31,238,31,240,31,187,31,152,31,152,31,63,31,148,31,153,31,153,30,153,29,78,31,224,31,213,31,213,30,6,31,113,31,218,31,176,31,199,31,199,30,211,31,187,31,73,31,236,31,135,31,250,31,3,31,91,31,47,31,47,30,15,31,36,31,36,30,180,31,153,31,153,30,173,31,106,31,240,31,240,30,163,31,9,31,251,31,120,31,120,30,120,29,235,31,149,31,197,31,5,31,75,31,75,30,75,29,53,31,53,30,223,31,223,30,33,31,167,31,111,31,105,31,159,31,102,31,102,30,102,29,102,28,204,31,204,30,226,31,34,31,131,31,210,31,210,30,210,29,182,31,98,31,98,30,98,29,108,31,218,31,71,31,145,31,208,31,94,31,159,31,159,30,159,29,4,31,4,30,81,31,152,31,228,31,250,31,250,30,161,31,87,31,8,31,8,30,8,29,8,28,226,31,47,31,152,31,169,31,108,31,108,30,108,29,145,31,70,31,70,30,50,31,50,30,50,29,188,31,17,31,93,31,93,30,239,31,254,31,178,31,178,30,195,31,210,31,190,31,157,31,157,30,44,31,44,30,108,31,97,31,42,31,230,31,166,31,5,31,90,31,253,31,162,31,137,31,185,31,186,31,220,31,235,31,219,31,19,31,112,31,195,31,150,31,154,31,154,30,30,31,167,31,247,31,233,31,127,31,8,31,8,30,192,31,122,31,126,31,66,31,135,31,135,30,234,31,65,31,157,31,83,31,208,31,94,31,174,31,172,31,219,31,127,31,196,31,158,31,81,31,80,31,80,30,83,31,51,31,231,31,96,31,96,30,130,31,15,31,245,31,182,31,208,31,196,31,196,30,205,31,129,31,165,31,165,30,175,31,175,30,175,29,175,28,50,31,84,31,159,31,159,30,150,31,156,31,191,31,204,31,143,31,174,31,183,31,49,31,188,31,38,31,38,30,183,31,110,31,214,31,155,31,123,31,176,31,57,31,102,31,219,31,181,31,172,31,208,31,171,31,171,30,6,31,137,31,25,31,25,30,144,31,19,31,27,31,129,31,181,31,52,31,163,31,25,31,25,30,25,29,77,31,255,31,255,30,170,31,23,31,33,31,150,31,38,31,91,31,118,31,211,31,179,31,179,30,226,31,5,31,210,31,210,30,31,31,56,31,56,30,223,31,184,31,245,31,245,30,143,31,103,31,103,30,191,31,87,31,137,31,200,31,201,31,136,31,120,31,215,31,158,31,45,31,214,31,30,31,30,30,30,29,97,31,9,31,129,31,232,31,190,31,89,31,199,31,24,31,22,31,68,31,68,30,190,31,137,31,118,31,18,31,237,31,74,31,173,31,75,31,156,31,120,31,13,31,191,31,104,31,220,31,200,31,176,31,101,31,62,31,223,31,232,31,227,31,227,30,163,31,181,31,181,30,181,29,156,31,139,31,124,31,124,30,86,31,86,30,238,31,238,30,142,31,95,31,212,31,93,31,61,31,61,30,234,31,176,31,131,31,144,31,24,31,107,31,107,30,161,31,107,31,117,31,167,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
