-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 456;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (21,0,151,0,0,0,18,0,158,0,160,0,0,0,0,0,0,0,222,0,175,0,116,0,192,0,228,0,143,0,0,0,116,0,96,0,203,0,176,0,85,0,0,0,245,0,215,0,205,0,78,0,109,0,81,0,0,0,116,0,242,0,2,0,62,0,154,0,65,0,36,0,144,0,0,0,22,0,60,0,129,0,253,0,38,0,227,0,96,0,18,0,175,0,152,0,0,0,165,0,174,0,0,0,213,0,127,0,171,0,213,0,202,0,0,0,44,0,239,0,42,0,198,0,201,0,157,0,79,0,219,0,0,0,71,0,0,0,51,0,133,0,245,0,145,0,54,0,0,0,24,0,210,0,0,0,143,0,68,0,182,0,0,0,80,0,147,0,75,0,0,0,165,0,43,0,40,0,75,0,148,0,30,0,0,0,18,0,149,0,216,0,133,0,0,0,32,0,165,0,0,0,39,0,238,0,21,0,110,0,249,0,214,0,184,0,134,0,61,0,90,0,0,0,0,0,0,0,209,0,228,0,40,0,0,0,0,0,91,0,78,0,238,0,249,0,42,0,59,0,139,0,253,0,0,0,250,0,33,0,206,0,71,0,189,0,42,0,83,0,0,0,28,0,207,0,92,0,0,0,29,0,162,0,189,0,50,0,0,0,0,0,148,0,238,0,226,0,138,0,196,0,179,0,0,0,9,0,218,0,0,0,91,0,238,0,198,0,253,0,46,0,16,0,157,0,215,0,0,0,86,0,19,0,215,0,0,0,103,0,125,0,29,0,96,0,0,0,58,0,151,0,143,0,231,0,150,0,226,0,193,0,205,0,183,0,92,0,13,0,216,0,242,0,0,0,226,0,0,0,207,0,0,0,84,0,17,0,252,0,0,0,10,0,47,0,78,0,237,0,228,0,155,0,202,0,154,0,0,0,0,0,90,0,0,0,153,0,192,0,178,0,34,0,48,0,221,0,87,0,0,0,212,0,230,0,175,0,220,0,220,0,0,0,6,0,241,0,32,0,0,0,69,0,147,0,31,0,0,0,43,0,139,0,145,0,0,0,215,0,21,0,38,0,37,0,250,0,74,0,109,0,183,0,25,0,59,0,246,0,127,0,231,0,163,0,43,0,30,0,0,0,28,0,144,0,219,0,162,0,22,0,245,0,105,0,215,0,226,0,237,0,78,0,0,0,0,0,111,0,92,0,0,0,242,0,227,0,13,0,220,0,218,0,56,0,0,0,68,0,0,0,54,0,241,0,69,0,61,0,35,0,69,0,140,0,34,0,163,0,198,0,0,0,98,0,37,0,200,0,96,0,22,0,166,0,154,0,58,0,128,0,17,0,33,0,193,0,0,0,185,0,0,0,220,0,7,0,211,0,42,0,74,0,142,0,0,0,49,0,208,0,208,0,95,0,53,0,41,0,134,0,57,0,41,0,0,0,61,0,38,0,121,0,165,0,139,0,50,0,76,0,0,0,0,0,53,0,71,0,95,0,73,0,0,0,0,0,128,0,157,0,13,0,0,0,41,0,117,0,165,0,237,0,179,0,0,0,196,0,114,0,204,0,114,0,0,0,0,0,5,0,145,0,124,0,5,0,197,0,33,0,151,0,146,0,247,0,87,0,0,0,96,0,80,0,164,0,64,0,46,0,19,0,0,0,92,0,17,0,0,0,0,0,112,0,227,0,136,0,0,0,218,0,101,0,162,0,0,0,161,0,232,0,77,0,29,0,134,0,0,0,66,0,0,0,229,0,32,0,8,0,166,0,118,0,131,0,233,0,79,0,0,0,0,0,75,0,9,0,25,0,147,0,77,0,174,0,176,0,89,0,101,0,0,0,137,0,0,0,109,0,97,0,61,0,138,0,155,0,134,0,7,0,151,0,0,0,165,0,163,0,0,0,249,0,132,0,19,0,120,0,35,0,68,0,0,0,124,0,204,0,246,0,116,0,0,0,214,0,64,0,14,0,0,0,0,0,249,0,0,0,203,0,37,0,128,0,157,0,96,0,0,0,0,0,139,0,0,0,236,0,204,0,0,0,131,0,221,0,0,0);
signal scenario_full  : scenario_type := (21,31,151,31,151,30,18,31,158,31,160,31,160,30,160,29,160,28,222,31,175,31,116,31,192,31,228,31,143,31,143,30,116,31,96,31,203,31,176,31,85,31,85,30,245,31,215,31,205,31,78,31,109,31,81,31,81,30,116,31,242,31,2,31,62,31,154,31,65,31,36,31,144,31,144,30,22,31,60,31,129,31,253,31,38,31,227,31,96,31,18,31,175,31,152,31,152,30,165,31,174,31,174,30,213,31,127,31,171,31,213,31,202,31,202,30,44,31,239,31,42,31,198,31,201,31,157,31,79,31,219,31,219,30,71,31,71,30,51,31,133,31,245,31,145,31,54,31,54,30,24,31,210,31,210,30,143,31,68,31,182,31,182,30,80,31,147,31,75,31,75,30,165,31,43,31,40,31,75,31,148,31,30,31,30,30,18,31,149,31,216,31,133,31,133,30,32,31,165,31,165,30,39,31,238,31,21,31,110,31,249,31,214,31,184,31,134,31,61,31,90,31,90,30,90,29,90,28,209,31,228,31,40,31,40,30,40,29,91,31,78,31,238,31,249,31,42,31,59,31,139,31,253,31,253,30,250,31,33,31,206,31,71,31,189,31,42,31,83,31,83,30,28,31,207,31,92,31,92,30,29,31,162,31,189,31,50,31,50,30,50,29,148,31,238,31,226,31,138,31,196,31,179,31,179,30,9,31,218,31,218,30,91,31,238,31,198,31,253,31,46,31,16,31,157,31,215,31,215,30,86,31,19,31,215,31,215,30,103,31,125,31,29,31,96,31,96,30,58,31,151,31,143,31,231,31,150,31,226,31,193,31,205,31,183,31,92,31,13,31,216,31,242,31,242,30,226,31,226,30,207,31,207,30,84,31,17,31,252,31,252,30,10,31,47,31,78,31,237,31,228,31,155,31,202,31,154,31,154,30,154,29,90,31,90,30,153,31,192,31,178,31,34,31,48,31,221,31,87,31,87,30,212,31,230,31,175,31,220,31,220,31,220,30,6,31,241,31,32,31,32,30,69,31,147,31,31,31,31,30,43,31,139,31,145,31,145,30,215,31,21,31,38,31,37,31,250,31,74,31,109,31,183,31,25,31,59,31,246,31,127,31,231,31,163,31,43,31,30,31,30,30,28,31,144,31,219,31,162,31,22,31,245,31,105,31,215,31,226,31,237,31,78,31,78,30,78,29,111,31,92,31,92,30,242,31,227,31,13,31,220,31,218,31,56,31,56,30,68,31,68,30,54,31,241,31,69,31,61,31,35,31,69,31,140,31,34,31,163,31,198,31,198,30,98,31,37,31,200,31,96,31,22,31,166,31,154,31,58,31,128,31,17,31,33,31,193,31,193,30,185,31,185,30,220,31,7,31,211,31,42,31,74,31,142,31,142,30,49,31,208,31,208,31,95,31,53,31,41,31,134,31,57,31,41,31,41,30,61,31,38,31,121,31,165,31,139,31,50,31,76,31,76,30,76,29,53,31,71,31,95,31,73,31,73,30,73,29,128,31,157,31,13,31,13,30,41,31,117,31,165,31,237,31,179,31,179,30,196,31,114,31,204,31,114,31,114,30,114,29,5,31,145,31,124,31,5,31,197,31,33,31,151,31,146,31,247,31,87,31,87,30,96,31,80,31,164,31,64,31,46,31,19,31,19,30,92,31,17,31,17,30,17,29,112,31,227,31,136,31,136,30,218,31,101,31,162,31,162,30,161,31,232,31,77,31,29,31,134,31,134,30,66,31,66,30,229,31,32,31,8,31,166,31,118,31,131,31,233,31,79,31,79,30,79,29,75,31,9,31,25,31,147,31,77,31,174,31,176,31,89,31,101,31,101,30,137,31,137,30,109,31,97,31,61,31,138,31,155,31,134,31,7,31,151,31,151,30,165,31,163,31,163,30,249,31,132,31,19,31,120,31,35,31,68,31,68,30,124,31,204,31,246,31,116,31,116,30,214,31,64,31,14,31,14,30,14,29,249,31,249,30,203,31,37,31,128,31,157,31,96,31,96,30,96,29,139,31,139,30,236,31,204,31,204,30,131,31,221,31,221,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
