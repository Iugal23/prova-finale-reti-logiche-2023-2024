-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_678 is
end project_tb_678;

architecture project_tb_arch_678 of project_tb_678 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 718;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (149,0,30,0,6,0,173,0,255,0,0,0,92,0,111,0,87,0,96,0,17,0,31,0,233,0,0,0,201,0,80,0,132,0,130,0,40,0,183,0,65,0,208,0,0,0,175,0,120,0,249,0,224,0,17,0,175,0,148,0,219,0,0,0,69,0,119,0,0,0,0,0,93,0,140,0,0,0,160,0,33,0,111,0,0,0,98,0,61,0,163,0,213,0,21,0,51,0,0,0,87,0,137,0,210,0,0,0,17,0,126,0,78,0,0,0,68,0,151,0,196,0,138,0,122,0,230,0,123,0,203,0,143,0,55,0,10,0,6,0,138,0,116,0,101,0,231,0,0,0,193,0,192,0,221,0,0,0,0,0,233,0,26,0,106,0,169,0,127,0,125,0,183,0,0,0,0,0,224,0,38,0,0,0,217,0,212,0,167,0,0,0,25,0,226,0,0,0,211,0,0,0,81,0,162,0,135,0,140,0,0,0,175,0,4,0,0,0,210,0,0,0,0,0,145,0,178,0,227,0,0,0,221,0,95,0,230,0,110,0,0,0,0,0,0,0,221,0,124,0,101,0,246,0,144,0,0,0,29,0,7,0,98,0,36,0,0,0,124,0,0,0,146,0,251,0,0,0,123,0,179,0,105,0,30,0,144,0,24,0,89,0,168,0,40,0,100,0,150,0,207,0,0,0,62,0,27,0,222,0,157,0,26,0,171,0,221,0,48,0,202,0,5,0,224,0,0,0,114,0,151,0,0,0,178,0,128,0,219,0,208,0,156,0,59,0,0,0,199,0,170,0,0,0,67,0,0,0,50,0,19,0,199,0,0,0,0,0,7,0,87,0,0,0,226,0,85,0,0,0,86,0,242,0,56,0,89,0,83,0,0,0,188,0,117,0,118,0,64,0,0,0,56,0,113,0,144,0,142,0,88,0,0,0,70,0,81,0,195,0,0,0,106,0,4,0,239,0,0,0,140,0,238,0,247,0,50,0,144,0,0,0,233,0,33,0,188,0,21,0,0,0,187,0,34,0,0,0,0,0,95,0,184,0,211,0,120,0,0,0,66,0,137,0,12,0,237,0,164,0,44,0,115,0,126,0,94,0,150,0,228,0,201,0,163,0,48,0,109,0,177,0,90,0,0,0,117,0,0,0,0,0,224,0,166,0,0,0,66,0,143,0,76,0,41,0,233,0,86,0,183,0,57,0,43,0,16,0,147,0,0,0,8,0,113,0,221,0,79,0,0,0,0,0,130,0,174,0,104,0,0,0,165,0,30,0,235,0,188,0,0,0,110,0,53,0,0,0,5,0,0,0,67,0,53,0,127,0,166,0,139,0,192,0,175,0,73,0,91,0,52,0,146,0,54,0,29,0,224,0,60,0,39,0,118,0,173,0,9,0,206,0,181,0,168,0,14,0,0,0,56,0,91,0,210,0,183,0,80,0,185,0,164,0,168,0,65,0,179,0,207,0,171,0,37,0,155,0,39,0,190,0,86,0,146,0,0,0,207,0,0,0,105,0,124,0,164,0,224,0,200,0,187,0,99,0,244,0,73,0,128,0,0,0,60,0,34,0,13,0,37,0,99,0,33,0,175,0,75,0,0,0,10,0,12,0,72,0,0,0,178,0,213,0,196,0,232,0,156,0,244,0,187,0,113,0,0,0,102,0,240,0,0,0,0,0,140,0,0,0,172,0,200,0,0,0,11,0,17,0,231,0,35,0,246,0,194,0,132,0,60,0,68,0,122,0,170,0,101,0,106,0,79,0,11,0,0,0,151,0,151,0,5,0,143,0,38,0,156,0,0,0,196,0,171,0,221,0,0,0,192,0,7,0,63,0,0,0,106,0,104,0,234,0,63,0,202,0,0,0,61,0,240,0,141,0,130,0,80,0,209,0,110,0,248,0,164,0,0,0,83,0,165,0,29,0,83,0,213,0,0,0,169,0,164,0,84,0,46,0,74,0,92,0,119,0,62,0,250,0,11,0,20,0,218,0,89,0,220,0,144,0,215,0,0,0,61,0,9,0,193,0,161,0,155,0,62,0,215,0,174,0,12,0,22,0,114,0,213,0,0,0,221,0,162,0,10,0,0,0,23,0,13,0,175,0,209,0,6,0,223,0,168,0,0,0,243,0,165,0,162,0,179,0,245,0,200,0,187,0,156,0,0,0,0,0,246,0,0,0,153,0,17,0,240,0,44,0,58,0,135,0,72,0,229,0,254,0,63,0,36,0,31,0,122,0,68,0,248,0,147,0,111,0,10,0,145,0,226,0,171,0,205,0,0,0,172,0,0,0,36,0,181,0,151,0,105,0,0,0,93,0,0,0,152,0,122,0,251,0,67,0,0,0,83,0,0,0,160,0,88,0,251,0,172,0,212,0,68,0,107,0,59,0,158,0,77,0,0,0,51,0,133,0,252,0,237,0,190,0,0,0,0,0,93,0,228,0,52,0,233,0,111,0,200,0,218,0,236,0,11,0,0,0,179,0,0,0,29,0,219,0,118,0,0,0,0,0,170,0,0,0,229,0,16,0,0,0,135,0,25,0,196,0,0,0,67,0,33,0,86,0,207,0,201,0,71,0,0,0,207,0,181,0,32,0,220,0,153,0,224,0,203,0,137,0,190,0,12,0,80,0,244,0,42,0,238,0,0,0,177,0,234,0,153,0,0,0,175,0,99,0,158,0,224,0,205,0,0,0,103,0,58,0,204,0,0,0,0,0,224,0,242,0,0,0,0,0,0,0,173,0,103,0,36,0,226,0,116,0,125,0,0,0,0,0,241,0,0,0,37,0,54,0,83,0,16,0,149,0,100,0,151,0,86,0,124,0,244,0,122,0,175,0,49,0,10,0,68,0,38,0,65,0,153,0,203,0,84,0,0,0,166,0,254,0,25,0,79,0,82,0,177,0,92,0,0,0,170,0,80,0,40,0,102,0,106,0,177,0,0,0,144,0,0,0,115,0,0,0,0,0,4,0,123,0,0,0,0,0,75,0,157,0,0,0,60,0,28,0,11,0,0,0,0,0,32,0,77,0,7,0,134,0,198,0,0,0,154,0,43,0,250,0,31,0,183,0,219,0,136,0,135,0,64,0,59,0,0,0,89,0,39,0,15,0,10,0,0,0,45,0,255,0,251,0,109,0,178,0,0,0,9,0,0,0,59,0,0,0,45,0,0,0,0,0,0,0,164,0,162,0,68,0,0,0,248,0,136,0,121,0,10,0,147,0);
signal scenario_full  : scenario_type := (149,31,30,31,6,31,173,31,255,31,255,30,92,31,111,31,87,31,96,31,17,31,31,31,233,31,233,30,201,31,80,31,132,31,130,31,40,31,183,31,65,31,208,31,208,30,175,31,120,31,249,31,224,31,17,31,175,31,148,31,219,31,219,30,69,31,119,31,119,30,119,29,93,31,140,31,140,30,160,31,33,31,111,31,111,30,98,31,61,31,163,31,213,31,21,31,51,31,51,30,87,31,137,31,210,31,210,30,17,31,126,31,78,31,78,30,68,31,151,31,196,31,138,31,122,31,230,31,123,31,203,31,143,31,55,31,10,31,6,31,138,31,116,31,101,31,231,31,231,30,193,31,192,31,221,31,221,30,221,29,233,31,26,31,106,31,169,31,127,31,125,31,183,31,183,30,183,29,224,31,38,31,38,30,217,31,212,31,167,31,167,30,25,31,226,31,226,30,211,31,211,30,81,31,162,31,135,31,140,31,140,30,175,31,4,31,4,30,210,31,210,30,210,29,145,31,178,31,227,31,227,30,221,31,95,31,230,31,110,31,110,30,110,29,110,28,221,31,124,31,101,31,246,31,144,31,144,30,29,31,7,31,98,31,36,31,36,30,124,31,124,30,146,31,251,31,251,30,123,31,179,31,105,31,30,31,144,31,24,31,89,31,168,31,40,31,100,31,150,31,207,31,207,30,62,31,27,31,222,31,157,31,26,31,171,31,221,31,48,31,202,31,5,31,224,31,224,30,114,31,151,31,151,30,178,31,128,31,219,31,208,31,156,31,59,31,59,30,199,31,170,31,170,30,67,31,67,30,50,31,19,31,199,31,199,30,199,29,7,31,87,31,87,30,226,31,85,31,85,30,86,31,242,31,56,31,89,31,83,31,83,30,188,31,117,31,118,31,64,31,64,30,56,31,113,31,144,31,142,31,88,31,88,30,70,31,81,31,195,31,195,30,106,31,4,31,239,31,239,30,140,31,238,31,247,31,50,31,144,31,144,30,233,31,33,31,188,31,21,31,21,30,187,31,34,31,34,30,34,29,95,31,184,31,211,31,120,31,120,30,66,31,137,31,12,31,237,31,164,31,44,31,115,31,126,31,94,31,150,31,228,31,201,31,163,31,48,31,109,31,177,31,90,31,90,30,117,31,117,30,117,29,224,31,166,31,166,30,66,31,143,31,76,31,41,31,233,31,86,31,183,31,57,31,43,31,16,31,147,31,147,30,8,31,113,31,221,31,79,31,79,30,79,29,130,31,174,31,104,31,104,30,165,31,30,31,235,31,188,31,188,30,110,31,53,31,53,30,5,31,5,30,67,31,53,31,127,31,166,31,139,31,192,31,175,31,73,31,91,31,52,31,146,31,54,31,29,31,224,31,60,31,39,31,118,31,173,31,9,31,206,31,181,31,168,31,14,31,14,30,56,31,91,31,210,31,183,31,80,31,185,31,164,31,168,31,65,31,179,31,207,31,171,31,37,31,155,31,39,31,190,31,86,31,146,31,146,30,207,31,207,30,105,31,124,31,164,31,224,31,200,31,187,31,99,31,244,31,73,31,128,31,128,30,60,31,34,31,13,31,37,31,99,31,33,31,175,31,75,31,75,30,10,31,12,31,72,31,72,30,178,31,213,31,196,31,232,31,156,31,244,31,187,31,113,31,113,30,102,31,240,31,240,30,240,29,140,31,140,30,172,31,200,31,200,30,11,31,17,31,231,31,35,31,246,31,194,31,132,31,60,31,68,31,122,31,170,31,101,31,106,31,79,31,11,31,11,30,151,31,151,31,5,31,143,31,38,31,156,31,156,30,196,31,171,31,221,31,221,30,192,31,7,31,63,31,63,30,106,31,104,31,234,31,63,31,202,31,202,30,61,31,240,31,141,31,130,31,80,31,209,31,110,31,248,31,164,31,164,30,83,31,165,31,29,31,83,31,213,31,213,30,169,31,164,31,84,31,46,31,74,31,92,31,119,31,62,31,250,31,11,31,20,31,218,31,89,31,220,31,144,31,215,31,215,30,61,31,9,31,193,31,161,31,155,31,62,31,215,31,174,31,12,31,22,31,114,31,213,31,213,30,221,31,162,31,10,31,10,30,23,31,13,31,175,31,209,31,6,31,223,31,168,31,168,30,243,31,165,31,162,31,179,31,245,31,200,31,187,31,156,31,156,30,156,29,246,31,246,30,153,31,17,31,240,31,44,31,58,31,135,31,72,31,229,31,254,31,63,31,36,31,31,31,122,31,68,31,248,31,147,31,111,31,10,31,145,31,226,31,171,31,205,31,205,30,172,31,172,30,36,31,181,31,151,31,105,31,105,30,93,31,93,30,152,31,122,31,251,31,67,31,67,30,83,31,83,30,160,31,88,31,251,31,172,31,212,31,68,31,107,31,59,31,158,31,77,31,77,30,51,31,133,31,252,31,237,31,190,31,190,30,190,29,93,31,228,31,52,31,233,31,111,31,200,31,218,31,236,31,11,31,11,30,179,31,179,30,29,31,219,31,118,31,118,30,118,29,170,31,170,30,229,31,16,31,16,30,135,31,25,31,196,31,196,30,67,31,33,31,86,31,207,31,201,31,71,31,71,30,207,31,181,31,32,31,220,31,153,31,224,31,203,31,137,31,190,31,12,31,80,31,244,31,42,31,238,31,238,30,177,31,234,31,153,31,153,30,175,31,99,31,158,31,224,31,205,31,205,30,103,31,58,31,204,31,204,30,204,29,224,31,242,31,242,30,242,29,242,28,173,31,103,31,36,31,226,31,116,31,125,31,125,30,125,29,241,31,241,30,37,31,54,31,83,31,16,31,149,31,100,31,151,31,86,31,124,31,244,31,122,31,175,31,49,31,10,31,68,31,38,31,65,31,153,31,203,31,84,31,84,30,166,31,254,31,25,31,79,31,82,31,177,31,92,31,92,30,170,31,80,31,40,31,102,31,106,31,177,31,177,30,144,31,144,30,115,31,115,30,115,29,4,31,123,31,123,30,123,29,75,31,157,31,157,30,60,31,28,31,11,31,11,30,11,29,32,31,77,31,7,31,134,31,198,31,198,30,154,31,43,31,250,31,31,31,183,31,219,31,136,31,135,31,64,31,59,31,59,30,89,31,39,31,15,31,10,31,10,30,45,31,255,31,251,31,109,31,178,31,178,30,9,31,9,30,59,31,59,30,45,31,45,30,45,29,45,28,164,31,162,31,68,31,68,30,248,31,136,31,121,31,10,31,147,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
