-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_822 is
end project_tb_822;

architecture project_tb_arch_822 of project_tb_822 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 675;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (178,0,91,0,234,0,92,0,192,0,89,0,0,0,0,0,101,0,132,0,73,0,103,0,142,0,239,0,87,0,180,0,0,0,109,0,159,0,0,0,209,0,0,0,0,0,0,0,26,0,3,0,0,0,185,0,101,0,11,0,0,0,0,0,35,0,64,0,232,0,19,0,14,0,181,0,60,0,51,0,110,0,222,0,213,0,0,0,245,0,93,0,117,0,0,0,196,0,86,0,0,0,38,0,0,0,0,0,1,0,141,0,197,0,172,0,0,0,2,0,219,0,53,0,79,0,185,0,81,0,66,0,131,0,72,0,213,0,240,0,190,0,125,0,36,0,0,0,158,0,170,0,0,0,251,0,76,0,17,0,9,0,40,0,115,0,43,0,148,0,230,0,43,0,0,0,0,0,146,0,143,0,0,0,225,0,239,0,18,0,0,0,146,0,228,0,135,0,56,0,52,0,164,0,169,0,0,0,53,0,120,0,48,0,137,0,222,0,53,0,64,0,122,0,0,0,0,0,58,0,241,0,47,0,11,0,27,0,0,0,244,0,152,0,227,0,10,0,103,0,0,0,147,0,195,0,136,0,149,0,56,0,0,0,0,0,0,0,251,0,198,0,219,0,207,0,249,0,89,0,0,0,40,0,144,0,232,0,0,0,142,0,0,0,83,0,255,0,72,0,246,0,37,0,26,0,24,0,179,0,156,0,107,0,105,0,16,0,193,0,183,0,152,0,129,0,198,0,0,0,241,0,129,0,82,0,238,0,186,0,0,0,151,0,63,0,211,0,240,0,140,0,0,0,226,0,0,0,202,0,221,0,0,0,253,0,138,0,201,0,0,0,170,0,229,0,16,0,113,0,208,0,0,0,229,0,56,0,0,0,209,0,58,0,31,0,92,0,212,0,16,0,74,0,211,0,222,0,233,0,75,0,106,0,29,0,0,0,82,0,0,0,136,0,42,0,93,0,227,0,126,0,0,0,240,0,201,0,63,0,120,0,95,0,71,0,210,0,89,0,0,0,24,0,143,0,0,0,140,0,104,0,220,0,5,0,27,0,69,0,194,0,183,0,0,0,145,0,79,0,168,0,234,0,201,0,0,0,121,0,190,0,0,0,247,0,28,0,119,0,226,0,71,0,111,0,173,0,61,0,4,0,233,0,248,0,169,0,117,0,0,0,247,0,0,0,0,0,134,0,0,0,116,0,24,0,126,0,103,0,0,0,0,0,133,0,74,0,0,0,157,0,206,0,0,0,253,0,95,0,184,0,169,0,0,0,0,0,185,0,50,0,162,0,97,0,0,0,171,0,42,0,26,0,186,0,225,0,37,0,165,0,160,0,224,0,121,0,114,0,224,0,0,0,205,0,0,0,207,0,127,0,143,0,247,0,0,0,18,0,228,0,142,0,117,0,37,0,0,0,156,0,239,0,19,0,112,0,15,0,14,0,35,0,107,0,171,0,0,0,106,0,109,0,20,0,143,0,0,0,236,0,93,0,0,0,241,0,109,0,0,0,0,0,67,0,192,0,145,0,3,0,226,0,161,0,167,0,70,0,43,0,51,0,110,0,209,0,0,0,135,0,72,0,147,0,44,0,109,0,58,0,42,0,91,0,86,0,5,0,153,0,141,0,249,0,198,0,222,0,0,0,159,0,0,0,68,0,55,0,187,0,4,0,78,0,0,0,82,0,0,0,51,0,182,0,170,0,213,0,224,0,229,0,22,0,243,0,179,0,100,0,91,0,254,0,0,0,0,0,75,0,207,0,137,0,0,0,83,0,134,0,162,0,103,0,172,0,0,0,203,0,188,0,81,0,254,0,15,0,179,0,80,0,43,0,189,0,215,0,0,0,6,0,0,0,0,0,0,0,205,0,144,0,10,0,71,0,120,0,170,0,215,0,145,0,160,0,43,0,132,0,58,0,114,0,20,0,169,0,0,0,91,0,48,0,197,0,86,0,121,0,168,0,253,0,249,0,100,0,176,0,161,0,0,0,0,0,0,0,57,0,0,0,0,0,0,0,73,0,167,0,0,0,0,0,0,0,30,0,157,0,239,0,89,0,83,0,0,0,154,0,211,0,140,0,68,0,153,0,97,0,228,0,126,0,67,0,0,0,106,0,66,0,148,0,0,0,44,0,147,0,63,0,94,0,114,0,225,0,125,0,74,0,114,0,179,0,166,0,126,0,126,0,65,0,0,0,48,0,22,0,219,0,240,0,249,0,0,0,71,0,41,0,229,0,38,0,81,0,61,0,240,0,4,0,0,0,3,0,127,0,146,0,144,0,152,0,179,0,113,0,0,0,52,0,0,0,1,0,242,0,65,0,242,0,143,0,3,0,39,0,170,0,100,0,213,0,44,0,203,0,112,0,154,0,202,0,0,0,65,0,68,0,0,0,95,0,159,0,164,0,0,0,251,0,146,0,30,0,0,0,134,0,212,0,0,0,22,0,129,0,0,0,0,0,20,0,34,0,153,0,237,0,170,0,88,0,255,0,37,0,253,0,184,0,233,0,228,0,81,0,90,0,106,0,31,0,202,0,178,0,128,0,125,0,206,0,4,0,33,0,204,0,118,0,128,0,244,0,0,0,154,0,92,0,0,0,62,0,202,0,199,0,187,0,3,0,36,0,8,0,62,0,51,0,124,0,185,0,0,0,0,0,0,0,0,0,158,0,0,0,0,0,0,0,195,0,6,0,89,0,42,0,177,0,0,0,0,0,65,0,95,0,0,0,235,0,0,0,95,0,0,0,216,0,0,0,105,0,149,0,0,0,85,0,184,0,145,0,229,0,134,0,0,0,0,0,0,0,96,0,164,0,33,0,9,0,0,0,11,0,153,0,0,0,19,0,245,0,0,0,237,0,195,0,12,0,0,0,204,0,172,0,0,0,252,0,74,0,14,0,71,0,11,0,0,0,169,0,97,0,171,0,231,0,160,0,87,0,160,0,7,0,113,0,181,0,34,0,22,0,83,0,0,0,135,0,92,0,102,0,201,0,119,0,55,0,87,0,72,0,0,0,143,0,0,0,0,0);
signal scenario_full  : scenario_type := (178,31,91,31,234,31,92,31,192,31,89,31,89,30,89,29,101,31,132,31,73,31,103,31,142,31,239,31,87,31,180,31,180,30,109,31,159,31,159,30,209,31,209,30,209,29,209,28,26,31,3,31,3,30,185,31,101,31,11,31,11,30,11,29,35,31,64,31,232,31,19,31,14,31,181,31,60,31,51,31,110,31,222,31,213,31,213,30,245,31,93,31,117,31,117,30,196,31,86,31,86,30,38,31,38,30,38,29,1,31,141,31,197,31,172,31,172,30,2,31,219,31,53,31,79,31,185,31,81,31,66,31,131,31,72,31,213,31,240,31,190,31,125,31,36,31,36,30,158,31,170,31,170,30,251,31,76,31,17,31,9,31,40,31,115,31,43,31,148,31,230,31,43,31,43,30,43,29,146,31,143,31,143,30,225,31,239,31,18,31,18,30,146,31,228,31,135,31,56,31,52,31,164,31,169,31,169,30,53,31,120,31,48,31,137,31,222,31,53,31,64,31,122,31,122,30,122,29,58,31,241,31,47,31,11,31,27,31,27,30,244,31,152,31,227,31,10,31,103,31,103,30,147,31,195,31,136,31,149,31,56,31,56,30,56,29,56,28,251,31,198,31,219,31,207,31,249,31,89,31,89,30,40,31,144,31,232,31,232,30,142,31,142,30,83,31,255,31,72,31,246,31,37,31,26,31,24,31,179,31,156,31,107,31,105,31,16,31,193,31,183,31,152,31,129,31,198,31,198,30,241,31,129,31,82,31,238,31,186,31,186,30,151,31,63,31,211,31,240,31,140,31,140,30,226,31,226,30,202,31,221,31,221,30,253,31,138,31,201,31,201,30,170,31,229,31,16,31,113,31,208,31,208,30,229,31,56,31,56,30,209,31,58,31,31,31,92,31,212,31,16,31,74,31,211,31,222,31,233,31,75,31,106,31,29,31,29,30,82,31,82,30,136,31,42,31,93,31,227,31,126,31,126,30,240,31,201,31,63,31,120,31,95,31,71,31,210,31,89,31,89,30,24,31,143,31,143,30,140,31,104,31,220,31,5,31,27,31,69,31,194,31,183,31,183,30,145,31,79,31,168,31,234,31,201,31,201,30,121,31,190,31,190,30,247,31,28,31,119,31,226,31,71,31,111,31,173,31,61,31,4,31,233,31,248,31,169,31,117,31,117,30,247,31,247,30,247,29,134,31,134,30,116,31,24,31,126,31,103,31,103,30,103,29,133,31,74,31,74,30,157,31,206,31,206,30,253,31,95,31,184,31,169,31,169,30,169,29,185,31,50,31,162,31,97,31,97,30,171,31,42,31,26,31,186,31,225,31,37,31,165,31,160,31,224,31,121,31,114,31,224,31,224,30,205,31,205,30,207,31,127,31,143,31,247,31,247,30,18,31,228,31,142,31,117,31,37,31,37,30,156,31,239,31,19,31,112,31,15,31,14,31,35,31,107,31,171,31,171,30,106,31,109,31,20,31,143,31,143,30,236,31,93,31,93,30,241,31,109,31,109,30,109,29,67,31,192,31,145,31,3,31,226,31,161,31,167,31,70,31,43,31,51,31,110,31,209,31,209,30,135,31,72,31,147,31,44,31,109,31,58,31,42,31,91,31,86,31,5,31,153,31,141,31,249,31,198,31,222,31,222,30,159,31,159,30,68,31,55,31,187,31,4,31,78,31,78,30,82,31,82,30,51,31,182,31,170,31,213,31,224,31,229,31,22,31,243,31,179,31,100,31,91,31,254,31,254,30,254,29,75,31,207,31,137,31,137,30,83,31,134,31,162,31,103,31,172,31,172,30,203,31,188,31,81,31,254,31,15,31,179,31,80,31,43,31,189,31,215,31,215,30,6,31,6,30,6,29,6,28,205,31,144,31,10,31,71,31,120,31,170,31,215,31,145,31,160,31,43,31,132,31,58,31,114,31,20,31,169,31,169,30,91,31,48,31,197,31,86,31,121,31,168,31,253,31,249,31,100,31,176,31,161,31,161,30,161,29,161,28,57,31,57,30,57,29,57,28,73,31,167,31,167,30,167,29,167,28,30,31,157,31,239,31,89,31,83,31,83,30,154,31,211,31,140,31,68,31,153,31,97,31,228,31,126,31,67,31,67,30,106,31,66,31,148,31,148,30,44,31,147,31,63,31,94,31,114,31,225,31,125,31,74,31,114,31,179,31,166,31,126,31,126,31,65,31,65,30,48,31,22,31,219,31,240,31,249,31,249,30,71,31,41,31,229,31,38,31,81,31,61,31,240,31,4,31,4,30,3,31,127,31,146,31,144,31,152,31,179,31,113,31,113,30,52,31,52,30,1,31,242,31,65,31,242,31,143,31,3,31,39,31,170,31,100,31,213,31,44,31,203,31,112,31,154,31,202,31,202,30,65,31,68,31,68,30,95,31,159,31,164,31,164,30,251,31,146,31,30,31,30,30,134,31,212,31,212,30,22,31,129,31,129,30,129,29,20,31,34,31,153,31,237,31,170,31,88,31,255,31,37,31,253,31,184,31,233,31,228,31,81,31,90,31,106,31,31,31,202,31,178,31,128,31,125,31,206,31,4,31,33,31,204,31,118,31,128,31,244,31,244,30,154,31,92,31,92,30,62,31,202,31,199,31,187,31,3,31,36,31,8,31,62,31,51,31,124,31,185,31,185,30,185,29,185,28,185,27,158,31,158,30,158,29,158,28,195,31,6,31,89,31,42,31,177,31,177,30,177,29,65,31,95,31,95,30,235,31,235,30,95,31,95,30,216,31,216,30,105,31,149,31,149,30,85,31,184,31,145,31,229,31,134,31,134,30,134,29,134,28,96,31,164,31,33,31,9,31,9,30,11,31,153,31,153,30,19,31,245,31,245,30,237,31,195,31,12,31,12,30,204,31,172,31,172,30,252,31,74,31,14,31,71,31,11,31,11,30,169,31,97,31,171,31,231,31,160,31,87,31,160,31,7,31,113,31,181,31,34,31,22,31,83,31,83,30,135,31,92,31,102,31,201,31,119,31,55,31,87,31,72,31,72,30,143,31,143,30,143,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
