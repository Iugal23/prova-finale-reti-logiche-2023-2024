-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_60 is
end project_tb_60;

architecture project_tb_arch_60 of project_tb_60 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1001;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (109,0,61,0,142,0,181,0,242,0,0,0,203,0,0,0,122,0,0,0,193,0,107,0,0,0,122,0,0,0,89,0,41,0,239,0,56,0,82,0,26,0,0,0,29,0,0,0,250,0,232,0,77,0,152,0,161,0,129,0,107,0,218,0,253,0,80,0,0,0,104,0,28,0,206,0,28,0,156,0,0,0,90,0,228,0,0,0,78,0,233,0,174,0,143,0,38,0,0,0,173,0,0,0,0,0,147,0,160,0,56,0,243,0,0,0,0,0,67,0,135,0,70,0,37,0,148,0,199,0,135,0,135,0,28,0,178,0,8,0,0,0,25,0,0,0,74,0,20,0,0,0,215,0,0,0,0,0,213,0,32,0,100,0,0,0,151,0,222,0,248,0,0,0,0,0,165,0,0,0,160,0,0,0,12,0,21,0,82,0,233,0,113,0,233,0,240,0,185,0,76,0,67,0,40,0,62,0,234,0,0,0,126,0,49,0,0,0,0,0,0,0,135,0,0,0,158,0,198,0,28,0,167,0,68,0,0,0,226,0,171,0,187,0,203,0,45,0,56,0,217,0,226,0,47,0,203,0,43,0,174,0,188,0,0,0,125,0,191,0,254,0,182,0,33,0,231,0,201,0,113,0,0,0,117,0,80,0,0,0,146,0,194,0,219,0,0,0,192,0,174,0,72,0,0,0,96,0,62,0,232,0,104,0,145,0,137,0,37,0,63,0,61,0,56,0,83,0,147,0,147,0,74,0,212,0,105,0,78,0,103,0,0,0,23,0,242,0,232,0,253,0,0,0,12,0,19,0,114,0,0,0,244,0,146,0,105,0,96,0,54,0,157,0,109,0,100,0,0,0,228,0,16,0,82,0,79,0,115,0,0,0,0,0,141,0,60,0,57,0,216,0,217,0,210,0,131,0,217,0,63,0,88,0,168,0,146,0,35,0,0,0,29,0,138,0,222,0,129,0,17,0,211,0,139,0,243,0,27,0,101,0,71,0,212,0,0,0,193,0,152,0,0,0,109,0,207,0,172,0,140,0,99,0,28,0,191,0,65,0,128,0,138,0,41,0,239,0,0,0,152,0,81,0,121,0,0,0,200,0,37,0,21,0,32,0,61,0,85,0,213,0,0,0,0,0,0,0,86,0,144,0,101,0,146,0,153,0,0,0,0,0,6,0,51,0,0,0,6,0,137,0,11,0,0,0,134,0,201,0,103,0,132,0,247,0,131,0,208,0,76,0,225,0,198,0,114,0,107,0,0,0,164,0,8,0,39,0,188,0,219,0,185,0,140,0,141,0,0,0,0,0,0,0,93,0,231,0,48,0,138,0,119,0,177,0,220,0,77,0,0,0,0,0,200,0,0,0,0,0,222,0,169,0,47,0,23,0,147,0,0,0,0,0,44,0,69,0,221,0,161,0,0,0,117,0,35,0,96,0,242,0,23,0,253,0,151,0,0,0,234,0,52,0,35,0,68,0,0,0,0,0,132,0,232,0,0,0,129,0,177,0,176,0,251,0,226,0,175,0,103,0,115,0,108,0,239,0,117,0,101,0,251,0,230,0,230,0,0,0,0,0,0,0,151,0,178,0,196,0,6,0,165,0,94,0,231,0,213,0,129,0,23,0,0,0,19,0,192,0,95,0,215,0,233,0,84,0,25,0,151,0,130,0,0,0,27,0,32,0,24,0,173,0,17,0,250,0,56,0,238,0,69,0,0,0,126,0,13,0,131,0,0,0,16,0,8,0,34,0,0,0,0,0,123,0,189,0,119,0,176,0,175,0,151,0,93,0,198,0,27,0,79,0,30,0,255,0,0,0,97,0,236,0,25,0,23,0,0,0,140,0,117,0,0,0,0,0,74,0,0,0,29,0,2,0,7,0,8,0,180,0,37,0,124,0,168,0,0,0,0,0,0,0,57,0,226,0,223,0,181,0,130,0,224,0,39,0,97,0,0,0,156,0,51,0,198,0,0,0,153,0,111,0,247,0,0,0,218,0,14,0,142,0,238,0,57,0,4,0,173,0,101,0,147,0,57,0,0,0,53,0,22,0,0,0,0,0,241,0,0,0,47,0,195,0,117,0,231,0,43,0,5,0,60,0,144,0,105,0,133,0,230,0,247,0,70,0,139,0,87,0,200,0,226,0,0,0,0,0,54,0,175,0,99,0,39,0,0,0,0,0,129,0,220,0,0,0,148,0,36,0,0,0,222,0,249,0,126,0,66,0,158,0,147,0,0,0,143,0,78,0,241,0,131,0,72,0,218,0,14,0,175,0,214,0,52,0,104,0,169,0,239,0,0,0,0,0,6,0,240,0,129,0,0,0,71,0,152,0,55,0,46,0,62,0,0,0,192,0,37,0,0,0,131,0,193,0,0,0,0,0,129,0,128,0,206,0,0,0,181,0,53,0,202,0,188,0,81,0,243,0,83,0,30,0,247,0,0,0,167,0,20,0,151,0,118,0,6,0,0,0,0,0,145,0,16,0,231,0,4,0,63,0,21,0,248,0,128,0,187,0,137,0,100,0,0,0,0,0,201,0,90,0,71,0,130,0,43,0,28,0,0,0,4,0,175,0,86,0,0,0,178,0,42,0,44,0,0,0,83,0,0,0,67,0,255,0,220,0,210,0,171,0,205,0,0,0,142,0,251,0,57,0,247,0,0,0,177,0,0,0,179,0,0,0,136,0,14,0,204,0,165,0,163,0,115,0,0,0,62,0,174,0,0,0,211,0,89,0,140,0,7,0,150,0,203,0,181,0,0,0,74,0,60,0,65,0,0,0,68,0,83,0,225,0,41,0,119,0,15,0,108,0,24,0,0,0,0,0,240,0,92,0,70,0,185,0,236,0,0,0,104,0,121,0,87,0,193,0,141,0,7,0,10,0,125,0,74,0,100,0,0,0,215,0,86,0,69,0,205,0,158,0,132,0,40,0,0,0,0,0,0,0,144,0,82,0,116,0,94,0,220,0,139,0,56,0,43,0,176,0,225,0,0,0,70,0,40,0,100,0,0,0,127,0,0,0,126,0,143,0,126,0,98,0,54,0,165,0,0,0,39,0,78,0,165,0,0,0,49,0,0,0,125,0,0,0,72,0,19,0,116,0,0,0,0,0,79,0,0,0,207,0,0,0,118,0,187,0,0,0,0,0,123,0,230,0,112,0,108,0,173,0,101,0,3,0,150,0,100,0,36,0,0,0,0,0,229,0,0,0,162,0,16,0,135,0,49,0,0,0,179,0,16,0,0,0,137,0,8,0,184,0,0,0,185,0,153,0,222,0,79,0,84,0,163,0,180,0,202,0,179,0,68,0,103,0,0,0,133,0,33,0,245,0,158,0,248,0,98,0,77,0,108,0,143,0,5,0,0,0,0,0,142,0,200,0,63,0,126,0,0,0,14,0,192,0,185,0,48,0,151,0,254,0,0,0,220,0,232,0,162,0,177,0,212,0,202,0,61,0,0,0,198,0,0,0,19,0,0,0,201,0,41,0,32,0,60,0,103,0,135,0,164,0,181,0,153,0,54,0,50,0,49,0,14,0,128,0,79,0,141,0,68,0,0,0,201,0,134,0,48,0,0,0,199,0,223,0,110,0,66,0,0,0,120,0,118,0,117,0,209,0,25,0,96,0,172,0,119,0,31,0,75,0,97,0,83,0,1,0,226,0,0,0,166,0,94,0,24,0,80,0,129,0,120,0,199,0,41,0,234,0,23,0,141,0,173,0,94,0,72,0,235,0,143,0,163,0,124,0,183,0,222,0,112,0,130,0,127,0,107,0,0,0,3,0,141,0,208,0,125,0,28,0,51,0,242,0,81,0,214,0,38,0,94,0,211,0,123,0,7,0,0,0,44,0,0,0,0,0,46,0,133,0,254,0,247,0,122,0,62,0,249,0,116,0,172,0,159,0,182,0,247,0,120,0,21,0,163,0,0,0,228,0,27,0,64,0,136,0,211,0,167,0,77,0,247,0,39,0,37,0,196,0,0,0,129,0,8,0,19,0,126,0,192,0,66,0,103,0,154,0,162,0,166,0,176,0,0,0,202,0,124,0,90,0,81,0,142,0,249,0,253,0,132,0,3,0,9,0,101,0,0,0,0,0,219,0,0,0,61,0,0,0,46,0,220,0,255,0,201,0,137,0,98,0,237,0,190,0,68,0,71,0,73,0,60,0,131,0,0,0,157,0,162,0,0,0,155,0,140,0,0,0,0,0,236,0,146,0,85,0,120,0,79,0,212,0,231,0,89,0,75,0,62,0,254,0,13,0,18,0,177,0,236,0,171,0,7,0,208,0,136,0,149,0,172,0,12,0,0,0,11,0,82,0,193,0,67,0,88,0,114,0,32,0,0,0,164,0,54,0,136,0,0,0,255,0,81,0,29,0,133,0,189,0,247,0,0,0,90,0,0,0,0,0,0,0,72,0,132,0,59,0,14,0,0,0,91,0,196,0,0,0,1,0,101,0,215,0,82,0,0,0,110,0,226,0,0,0);
signal scenario_full  : scenario_type := (109,31,61,31,142,31,181,31,242,31,242,30,203,31,203,30,122,31,122,30,193,31,107,31,107,30,122,31,122,30,89,31,41,31,239,31,56,31,82,31,26,31,26,30,29,31,29,30,250,31,232,31,77,31,152,31,161,31,129,31,107,31,218,31,253,31,80,31,80,30,104,31,28,31,206,31,28,31,156,31,156,30,90,31,228,31,228,30,78,31,233,31,174,31,143,31,38,31,38,30,173,31,173,30,173,29,147,31,160,31,56,31,243,31,243,30,243,29,67,31,135,31,70,31,37,31,148,31,199,31,135,31,135,31,28,31,178,31,8,31,8,30,25,31,25,30,74,31,20,31,20,30,215,31,215,30,215,29,213,31,32,31,100,31,100,30,151,31,222,31,248,31,248,30,248,29,165,31,165,30,160,31,160,30,12,31,21,31,82,31,233,31,113,31,233,31,240,31,185,31,76,31,67,31,40,31,62,31,234,31,234,30,126,31,49,31,49,30,49,29,49,28,135,31,135,30,158,31,198,31,28,31,167,31,68,31,68,30,226,31,171,31,187,31,203,31,45,31,56,31,217,31,226,31,47,31,203,31,43,31,174,31,188,31,188,30,125,31,191,31,254,31,182,31,33,31,231,31,201,31,113,31,113,30,117,31,80,31,80,30,146,31,194,31,219,31,219,30,192,31,174,31,72,31,72,30,96,31,62,31,232,31,104,31,145,31,137,31,37,31,63,31,61,31,56,31,83,31,147,31,147,31,74,31,212,31,105,31,78,31,103,31,103,30,23,31,242,31,232,31,253,31,253,30,12,31,19,31,114,31,114,30,244,31,146,31,105,31,96,31,54,31,157,31,109,31,100,31,100,30,228,31,16,31,82,31,79,31,115,31,115,30,115,29,141,31,60,31,57,31,216,31,217,31,210,31,131,31,217,31,63,31,88,31,168,31,146,31,35,31,35,30,29,31,138,31,222,31,129,31,17,31,211,31,139,31,243,31,27,31,101,31,71,31,212,31,212,30,193,31,152,31,152,30,109,31,207,31,172,31,140,31,99,31,28,31,191,31,65,31,128,31,138,31,41,31,239,31,239,30,152,31,81,31,121,31,121,30,200,31,37,31,21,31,32,31,61,31,85,31,213,31,213,30,213,29,213,28,86,31,144,31,101,31,146,31,153,31,153,30,153,29,6,31,51,31,51,30,6,31,137,31,11,31,11,30,134,31,201,31,103,31,132,31,247,31,131,31,208,31,76,31,225,31,198,31,114,31,107,31,107,30,164,31,8,31,39,31,188,31,219,31,185,31,140,31,141,31,141,30,141,29,141,28,93,31,231,31,48,31,138,31,119,31,177,31,220,31,77,31,77,30,77,29,200,31,200,30,200,29,222,31,169,31,47,31,23,31,147,31,147,30,147,29,44,31,69,31,221,31,161,31,161,30,117,31,35,31,96,31,242,31,23,31,253,31,151,31,151,30,234,31,52,31,35,31,68,31,68,30,68,29,132,31,232,31,232,30,129,31,177,31,176,31,251,31,226,31,175,31,103,31,115,31,108,31,239,31,117,31,101,31,251,31,230,31,230,31,230,30,230,29,230,28,151,31,178,31,196,31,6,31,165,31,94,31,231,31,213,31,129,31,23,31,23,30,19,31,192,31,95,31,215,31,233,31,84,31,25,31,151,31,130,31,130,30,27,31,32,31,24,31,173,31,17,31,250,31,56,31,238,31,69,31,69,30,126,31,13,31,131,31,131,30,16,31,8,31,34,31,34,30,34,29,123,31,189,31,119,31,176,31,175,31,151,31,93,31,198,31,27,31,79,31,30,31,255,31,255,30,97,31,236,31,25,31,23,31,23,30,140,31,117,31,117,30,117,29,74,31,74,30,29,31,2,31,7,31,8,31,180,31,37,31,124,31,168,31,168,30,168,29,168,28,57,31,226,31,223,31,181,31,130,31,224,31,39,31,97,31,97,30,156,31,51,31,198,31,198,30,153,31,111,31,247,31,247,30,218,31,14,31,142,31,238,31,57,31,4,31,173,31,101,31,147,31,57,31,57,30,53,31,22,31,22,30,22,29,241,31,241,30,47,31,195,31,117,31,231,31,43,31,5,31,60,31,144,31,105,31,133,31,230,31,247,31,70,31,139,31,87,31,200,31,226,31,226,30,226,29,54,31,175,31,99,31,39,31,39,30,39,29,129,31,220,31,220,30,148,31,36,31,36,30,222,31,249,31,126,31,66,31,158,31,147,31,147,30,143,31,78,31,241,31,131,31,72,31,218,31,14,31,175,31,214,31,52,31,104,31,169,31,239,31,239,30,239,29,6,31,240,31,129,31,129,30,71,31,152,31,55,31,46,31,62,31,62,30,192,31,37,31,37,30,131,31,193,31,193,30,193,29,129,31,128,31,206,31,206,30,181,31,53,31,202,31,188,31,81,31,243,31,83,31,30,31,247,31,247,30,167,31,20,31,151,31,118,31,6,31,6,30,6,29,145,31,16,31,231,31,4,31,63,31,21,31,248,31,128,31,187,31,137,31,100,31,100,30,100,29,201,31,90,31,71,31,130,31,43,31,28,31,28,30,4,31,175,31,86,31,86,30,178,31,42,31,44,31,44,30,83,31,83,30,67,31,255,31,220,31,210,31,171,31,205,31,205,30,142,31,251,31,57,31,247,31,247,30,177,31,177,30,179,31,179,30,136,31,14,31,204,31,165,31,163,31,115,31,115,30,62,31,174,31,174,30,211,31,89,31,140,31,7,31,150,31,203,31,181,31,181,30,74,31,60,31,65,31,65,30,68,31,83,31,225,31,41,31,119,31,15,31,108,31,24,31,24,30,24,29,240,31,92,31,70,31,185,31,236,31,236,30,104,31,121,31,87,31,193,31,141,31,7,31,10,31,125,31,74,31,100,31,100,30,215,31,86,31,69,31,205,31,158,31,132,31,40,31,40,30,40,29,40,28,144,31,82,31,116,31,94,31,220,31,139,31,56,31,43,31,176,31,225,31,225,30,70,31,40,31,100,31,100,30,127,31,127,30,126,31,143,31,126,31,98,31,54,31,165,31,165,30,39,31,78,31,165,31,165,30,49,31,49,30,125,31,125,30,72,31,19,31,116,31,116,30,116,29,79,31,79,30,207,31,207,30,118,31,187,31,187,30,187,29,123,31,230,31,112,31,108,31,173,31,101,31,3,31,150,31,100,31,36,31,36,30,36,29,229,31,229,30,162,31,16,31,135,31,49,31,49,30,179,31,16,31,16,30,137,31,8,31,184,31,184,30,185,31,153,31,222,31,79,31,84,31,163,31,180,31,202,31,179,31,68,31,103,31,103,30,133,31,33,31,245,31,158,31,248,31,98,31,77,31,108,31,143,31,5,31,5,30,5,29,142,31,200,31,63,31,126,31,126,30,14,31,192,31,185,31,48,31,151,31,254,31,254,30,220,31,232,31,162,31,177,31,212,31,202,31,61,31,61,30,198,31,198,30,19,31,19,30,201,31,41,31,32,31,60,31,103,31,135,31,164,31,181,31,153,31,54,31,50,31,49,31,14,31,128,31,79,31,141,31,68,31,68,30,201,31,134,31,48,31,48,30,199,31,223,31,110,31,66,31,66,30,120,31,118,31,117,31,209,31,25,31,96,31,172,31,119,31,31,31,75,31,97,31,83,31,1,31,226,31,226,30,166,31,94,31,24,31,80,31,129,31,120,31,199,31,41,31,234,31,23,31,141,31,173,31,94,31,72,31,235,31,143,31,163,31,124,31,183,31,222,31,112,31,130,31,127,31,107,31,107,30,3,31,141,31,208,31,125,31,28,31,51,31,242,31,81,31,214,31,38,31,94,31,211,31,123,31,7,31,7,30,44,31,44,30,44,29,46,31,133,31,254,31,247,31,122,31,62,31,249,31,116,31,172,31,159,31,182,31,247,31,120,31,21,31,163,31,163,30,228,31,27,31,64,31,136,31,211,31,167,31,77,31,247,31,39,31,37,31,196,31,196,30,129,31,8,31,19,31,126,31,192,31,66,31,103,31,154,31,162,31,166,31,176,31,176,30,202,31,124,31,90,31,81,31,142,31,249,31,253,31,132,31,3,31,9,31,101,31,101,30,101,29,219,31,219,30,61,31,61,30,46,31,220,31,255,31,201,31,137,31,98,31,237,31,190,31,68,31,71,31,73,31,60,31,131,31,131,30,157,31,162,31,162,30,155,31,140,31,140,30,140,29,236,31,146,31,85,31,120,31,79,31,212,31,231,31,89,31,75,31,62,31,254,31,13,31,18,31,177,31,236,31,171,31,7,31,208,31,136,31,149,31,172,31,12,31,12,30,11,31,82,31,193,31,67,31,88,31,114,31,32,31,32,30,164,31,54,31,136,31,136,30,255,31,81,31,29,31,133,31,189,31,247,31,247,30,90,31,90,30,90,29,90,28,72,31,132,31,59,31,14,31,14,30,91,31,196,31,196,30,1,31,101,31,215,31,82,31,82,30,110,31,226,31,226,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
