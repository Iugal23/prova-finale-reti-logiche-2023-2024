-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_263 is
end project_tb_263;

architecture project_tb_arch_263 of project_tb_263 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 667;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (140,0,124,0,113,0,34,0,73,0,0,0,135,0,193,0,36,0,192,0,92,0,170,0,0,0,60,0,189,0,140,0,207,0,238,0,50,0,203,0,103,0,0,0,21,0,71,0,234,0,46,0,25,0,0,0,95,0,56,0,226,0,140,0,216,0,141,0,0,0,151,0,155,0,74,0,114,0,255,0,16,0,221,0,182,0,62,0,0,0,54,0,245,0,154,0,228,0,13,0,204,0,34,0,117,0,71,0,0,0,110,0,0,0,180,0,35,0,117,0,246,0,177,0,198,0,125,0,128,0,103,0,73,0,82,0,0,0,219,0,80,0,224,0,0,0,0,0,251,0,0,0,128,0,180,0,93,0,18,0,68,0,116,0,36,0,27,0,185,0,87,0,74,0,0,0,229,0,0,0,29,0,238,0,4,0,222,0,195,0,38,0,158,0,187,0,158,0,0,0,229,0,35,0,234,0,194,0,0,0,48,0,34,0,221,0,150,0,0,0,0,0,119,0,0,0,190,0,152,0,0,0,241,0,144,0,73,0,40,0,50,0,78,0,116,0,52,0,0,0,107,0,0,0,127,0,195,0,0,0,158,0,152,0,39,0,150,0,217,0,222,0,160,0,199,0,0,0,0,0,29,0,80,0,167,0,201,0,86,0,40,0,16,0,138,0,237,0,115,0,0,0,169,0,0,0,5,0,46,0,39,0,182,0,30,0,253,0,158,0,20,0,46,0,246,0,149,0,244,0,79,0,57,0,28,0,1,0,5,0,0,0,240,0,21,0,45,0,147,0,0,0,198,0,198,0,191,0,144,0,174,0,165,0,81,0,55,0,248,0,0,0,147,0,159,0,240,0,219,0,0,0,152,0,0,0,194,0,228,0,13,0,158,0,214,0,17,0,8,0,122,0,160,0,64,0,0,0,230,0,191,0,11,0,216,0,82,0,96,0,78,0,117,0,172,0,214,0,3,0,21,0,180,0,221,0,0,0,240,0,97,0,60,0,114,0,239,0,0,0,141,0,196,0,0,0,0,0,72,0,234,0,0,0,98,0,32,0,0,0,145,0,252,0,223,0,0,0,174,0,246,0,210,0,19,0,148,0,0,0,91,0,39,0,0,0,213,0,52,0,245,0,50,0,144,0,213,0,254,0,197,0,16,0,6,0,66,0,0,0,0,0,181,0,104,0,142,0,132,0,229,0,214,0,137,0,52,0,0,0,54,0,189,0,0,0,33,0,126,0,0,0,119,0,0,0,215,0,0,0,226,0,64,0,159,0,62,0,0,0,145,0,0,0,121,0,82,0,206,0,128,0,128,0,47,0,72,0,53,0,227,0,0,0,226,0,0,0,0,0,89,0,118,0,249,0,183,0,66,0,199,0,40,0,0,0,55,0,63,0,0,0,0,0,153,0,21,0,139,0,0,0,0,0,255,0,0,0,214,0,109,0,0,0,240,0,56,0,0,0,179,0,8,0,240,0,85,0,46,0,240,0,54,0,118,0,231,0,37,0,105,0,0,0,236,0,251,0,107,0,85,0,218,0,227,0,31,0,72,0,249,0,0,0,95,0,124,0,0,0,6,0,119,0,0,0,39,0,26,0,0,0,237,0,0,0,0,0,144,0,57,0,22,0,106,0,117,0,0,0,0,0,72,0,129,0,197,0,143,0,0,0,195,0,71,0,206,0,0,0,247,0,43,0,66,0,59,0,0,0,248,0,78,0,245,0,151,0,197,0,18,0,0,0,86,0,43,0,240,0,17,0,10,0,186,0,221,0,93,0,0,0,102,0,66,0,82,0,208,0,0,0,216,0,205,0,236,0,97,0,0,0,76,0,0,0,0,0,89,0,189,0,230,0,214,0,48,0,80,0,142,0,0,0,64,0,0,0,0,0,19,0,241,0,72,0,63,0,93,0,25,0,0,0,204,0,213,0,147,0,153,0,0,0,180,0,134,0,234,0,0,0,74,0,0,0,253,0,9,0,0,0,70,0,222,0,0,0,0,0,136,0,39,0,0,0,51,0,0,0,241,0,126,0,104,0,217,0,0,0,73,0,68,0,156,0,198,0,117,0,11,0,160,0,0,0,20,0,158,0,19,0,126,0,22,0,0,0,225,0,17,0,84,0,35,0,99,0,203,0,10,0,101,0,133,0,184,0,43,0,162,0,217,0,187,0,60,0,214,0,48,0,210,0,201,0,109,0,197,0,174,0,35,0,65,0,65,0,0,0,11,0,227,0,0,0,0,0,67,0,235,0,32,0,206,0,0,0,60,0,104,0,234,0,251,0,13,0,255,0,66,0,210,0,0,0,235,0,148,0,0,0,212,0,1,0,29,0,1,0,0,0,86,0,91,0,0,0,119,0,212,0,105,0,0,0,164,0,100,0,0,0,71,0,0,0,144,0,164,0,228,0,132,0,0,0,56,0,0,0,196,0,175,0,200,0,109,0,166,0,252,0,87,0,153,0,16,0,89,0,84,0,0,0,126,0,41,0,185,0,221,0,0,0,82,0,168,0,50,0,155,0,0,0,240,0,91,0,206,0,80,0,42,0,80,0,75,0,151,0,218,0,15,0,0,0,103,0,183,0,0,0,171,0,0,0,0,0,141,0,57,0,129,0,0,0,85,0,72,0,28,0,141,0,123,0,253,0,140,0,123,0,0,0,131,0,0,0,250,0,71,0,206,0,134,0,210,0,181,0,255,0,24,0,222,0,207,0,44,0,98,0,134,0,91,0,4,0,0,0,208,0,50,0,255,0,108,0,196,0,0,0,16,0,62,0,152,0,121,0,214,0,0,0,192,0,192,0,61,0,0,0,35,0,244,0,183,0,231,0,41,0,17,0,110,0,164,0,174,0,184,0,219,0,0,0,249,0,26,0,0,0,233,0,22,0,58,0,45,0,118,0,131,0,99,0,16,0,245,0,0,0,207,0,232,0,0,0,52,0,93,0,0,0,0,0,224,0,251,0,97,0,220,0,145,0,78,0,118,0,38,0,0,0);
signal scenario_full  : scenario_type := (140,31,124,31,113,31,34,31,73,31,73,30,135,31,193,31,36,31,192,31,92,31,170,31,170,30,60,31,189,31,140,31,207,31,238,31,50,31,203,31,103,31,103,30,21,31,71,31,234,31,46,31,25,31,25,30,95,31,56,31,226,31,140,31,216,31,141,31,141,30,151,31,155,31,74,31,114,31,255,31,16,31,221,31,182,31,62,31,62,30,54,31,245,31,154,31,228,31,13,31,204,31,34,31,117,31,71,31,71,30,110,31,110,30,180,31,35,31,117,31,246,31,177,31,198,31,125,31,128,31,103,31,73,31,82,31,82,30,219,31,80,31,224,31,224,30,224,29,251,31,251,30,128,31,180,31,93,31,18,31,68,31,116,31,36,31,27,31,185,31,87,31,74,31,74,30,229,31,229,30,29,31,238,31,4,31,222,31,195,31,38,31,158,31,187,31,158,31,158,30,229,31,35,31,234,31,194,31,194,30,48,31,34,31,221,31,150,31,150,30,150,29,119,31,119,30,190,31,152,31,152,30,241,31,144,31,73,31,40,31,50,31,78,31,116,31,52,31,52,30,107,31,107,30,127,31,195,31,195,30,158,31,152,31,39,31,150,31,217,31,222,31,160,31,199,31,199,30,199,29,29,31,80,31,167,31,201,31,86,31,40,31,16,31,138,31,237,31,115,31,115,30,169,31,169,30,5,31,46,31,39,31,182,31,30,31,253,31,158,31,20,31,46,31,246,31,149,31,244,31,79,31,57,31,28,31,1,31,5,31,5,30,240,31,21,31,45,31,147,31,147,30,198,31,198,31,191,31,144,31,174,31,165,31,81,31,55,31,248,31,248,30,147,31,159,31,240,31,219,31,219,30,152,31,152,30,194,31,228,31,13,31,158,31,214,31,17,31,8,31,122,31,160,31,64,31,64,30,230,31,191,31,11,31,216,31,82,31,96,31,78,31,117,31,172,31,214,31,3,31,21,31,180,31,221,31,221,30,240,31,97,31,60,31,114,31,239,31,239,30,141,31,196,31,196,30,196,29,72,31,234,31,234,30,98,31,32,31,32,30,145,31,252,31,223,31,223,30,174,31,246,31,210,31,19,31,148,31,148,30,91,31,39,31,39,30,213,31,52,31,245,31,50,31,144,31,213,31,254,31,197,31,16,31,6,31,66,31,66,30,66,29,181,31,104,31,142,31,132,31,229,31,214,31,137,31,52,31,52,30,54,31,189,31,189,30,33,31,126,31,126,30,119,31,119,30,215,31,215,30,226,31,64,31,159,31,62,31,62,30,145,31,145,30,121,31,82,31,206,31,128,31,128,31,47,31,72,31,53,31,227,31,227,30,226,31,226,30,226,29,89,31,118,31,249,31,183,31,66,31,199,31,40,31,40,30,55,31,63,31,63,30,63,29,153,31,21,31,139,31,139,30,139,29,255,31,255,30,214,31,109,31,109,30,240,31,56,31,56,30,179,31,8,31,240,31,85,31,46,31,240,31,54,31,118,31,231,31,37,31,105,31,105,30,236,31,251,31,107,31,85,31,218,31,227,31,31,31,72,31,249,31,249,30,95,31,124,31,124,30,6,31,119,31,119,30,39,31,26,31,26,30,237,31,237,30,237,29,144,31,57,31,22,31,106,31,117,31,117,30,117,29,72,31,129,31,197,31,143,31,143,30,195,31,71,31,206,31,206,30,247,31,43,31,66,31,59,31,59,30,248,31,78,31,245,31,151,31,197,31,18,31,18,30,86,31,43,31,240,31,17,31,10,31,186,31,221,31,93,31,93,30,102,31,66,31,82,31,208,31,208,30,216,31,205,31,236,31,97,31,97,30,76,31,76,30,76,29,89,31,189,31,230,31,214,31,48,31,80,31,142,31,142,30,64,31,64,30,64,29,19,31,241,31,72,31,63,31,93,31,25,31,25,30,204,31,213,31,147,31,153,31,153,30,180,31,134,31,234,31,234,30,74,31,74,30,253,31,9,31,9,30,70,31,222,31,222,30,222,29,136,31,39,31,39,30,51,31,51,30,241,31,126,31,104,31,217,31,217,30,73,31,68,31,156,31,198,31,117,31,11,31,160,31,160,30,20,31,158,31,19,31,126,31,22,31,22,30,225,31,17,31,84,31,35,31,99,31,203,31,10,31,101,31,133,31,184,31,43,31,162,31,217,31,187,31,60,31,214,31,48,31,210,31,201,31,109,31,197,31,174,31,35,31,65,31,65,31,65,30,11,31,227,31,227,30,227,29,67,31,235,31,32,31,206,31,206,30,60,31,104,31,234,31,251,31,13,31,255,31,66,31,210,31,210,30,235,31,148,31,148,30,212,31,1,31,29,31,1,31,1,30,86,31,91,31,91,30,119,31,212,31,105,31,105,30,164,31,100,31,100,30,71,31,71,30,144,31,164,31,228,31,132,31,132,30,56,31,56,30,196,31,175,31,200,31,109,31,166,31,252,31,87,31,153,31,16,31,89,31,84,31,84,30,126,31,41,31,185,31,221,31,221,30,82,31,168,31,50,31,155,31,155,30,240,31,91,31,206,31,80,31,42,31,80,31,75,31,151,31,218,31,15,31,15,30,103,31,183,31,183,30,171,31,171,30,171,29,141,31,57,31,129,31,129,30,85,31,72,31,28,31,141,31,123,31,253,31,140,31,123,31,123,30,131,31,131,30,250,31,71,31,206,31,134,31,210,31,181,31,255,31,24,31,222,31,207,31,44,31,98,31,134,31,91,31,4,31,4,30,208,31,50,31,255,31,108,31,196,31,196,30,16,31,62,31,152,31,121,31,214,31,214,30,192,31,192,31,61,31,61,30,35,31,244,31,183,31,231,31,41,31,17,31,110,31,164,31,174,31,184,31,219,31,219,30,249,31,26,31,26,30,233,31,22,31,58,31,45,31,118,31,131,31,99,31,16,31,245,31,245,30,207,31,232,31,232,30,52,31,93,31,93,30,93,29,224,31,251,31,97,31,220,31,145,31,78,31,118,31,38,31,38,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
