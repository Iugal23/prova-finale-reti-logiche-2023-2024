-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_934 is
end project_tb_934;

architecture project_tb_arch_934 of project_tb_934 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 801;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (211,0,164,0,188,0,88,0,0,0,214,0,176,0,32,0,0,0,32,0,164,0,97,0,147,0,0,0,230,0,101,0,110,0,248,0,154,0,122,0,67,0,8,0,217,0,0,0,111,0,203,0,240,0,119,0,92,0,109,0,73,0,180,0,94,0,171,0,0,0,40,0,169,0,182,0,191,0,104,0,67,0,103,0,62,0,59,0,37,0,198,0,145,0,91,0,78,0,146,0,0,0,0,0,70,0,0,0,138,0,242,0,36,0,199,0,81,0,245,0,237,0,120,0,61,0,181,0,235,0,67,0,97,0,0,0,0,0,191,0,27,0,16,0,0,0,0,0,0,0,173,0,15,0,180,0,3,0,0,0,50,0,198,0,55,0,129,0,98,0,89,0,115,0,0,0,0,0,109,0,246,0,167,0,161,0,18,0,195,0,64,0,253,0,0,0,51,0,12,0,58,0,43,0,10,0,39,0,0,0,0,0,104,0,82,0,0,0,151,0,0,0,251,0,249,0,225,0,72,0,190,0,0,0,117,0,197,0,0,0,133,0,53,0,0,0,68,0,117,0,59,0,135,0,159,0,106,0,242,0,138,0,167,0,241,0,151,0,80,0,241,0,246,0,156,0,229,0,9,0,46,0,61,0,49,0,10,0,174,0,36,0,17,0,179,0,166,0,148,0,4,0,137,0,254,0,116,0,226,0,44,0,62,0,0,0,0,0,178,0,109,0,82,0,21,0,0,0,0,0,79,0,72,0,164,0,176,0,74,0,228,0,177,0,230,0,148,0,0,0,247,0,213,0,226,0,132,0,136,0,188,0,112,0,138,0,132,0,0,0,168,0,0,0,135,0,176,0,0,0,28,0,200,0,63,0,252,0,133,0,77,0,223,0,10,0,178,0,91,0,0,0,0,0,137,0,72,0,41,0,217,0,27,0,232,0,79,0,101,0,95,0,241,0,0,0,195,0,99,0,223,0,174,0,171,0,197,0,0,0,18,0,198,0,0,0,174,0,90,0,198,0,0,0,90,0,239,0,69,0,95,0,30,0,37,0,0,0,54,0,236,0,62,0,137,0,0,0,86,0,35,0,103,0,0,0,0,0,0,0,150,0,0,0,0,0,36,0,99,0,229,0,94,0,58,0,0,0,48,0,222,0,0,0,0,0,80,0,218,0,51,0,0,0,230,0,104,0,127,0,251,0,236,0,0,0,5,0,144,0,187,0,56,0,235,0,81,0,0,0,179,0,114,0,0,0,247,0,0,0,11,0,85,0,240,0,68,0,3,0,142,0,158,0,89,0,108,0,0,0,151,0,0,0,0,0,137,0,95,0,183,0,146,0,36,0,82,0,86,0,193,0,10,0,242,0,39,0,202,0,47,0,0,0,0,0,172,0,0,0,246,0,0,0,59,0,71,0,227,0,179,0,22,0,167,0,60,0,242,0,41,0,145,0,11,0,134,0,0,0,57,0,74,0,80,0,0,0,182,0,22,0,98,0,0,0,164,0,128,0,44,0,63,0,213,0,225,0,0,0,0,0,127,0,0,0,182,0,0,0,34,0,0,0,0,0,182,0,42,0,185,0,163,0,0,0,181,0,64,0,134,0,0,0,57,0,9,0,233,0,0,0,212,0,236,0,0,0,207,0,8,0,2,0,136,0,255,0,40,0,133,0,167,0,31,0,146,0,50,0,119,0,233,0,247,0,0,0,28,0,0,0,33,0,231,0,72,0,0,0,0,0,0,0,0,0,127,0,0,0,76,0,124,0,39,0,52,0,72,0,0,0,145,0,18,0,17,0,8,0,168,0,82,0,238,0,86,0,0,0,171,0,0,0,0,0,66,0,138,0,59,0,204,0,21,0,42,0,0,0,150,0,0,0,57,0,228,0,100,0,0,0,41,0,78,0,10,0,141,0,0,0,152,0,98,0,0,0,157,0,92,0,0,0,82,0,0,0,129,0,81,0,31,0,255,0,29,0,62,0,0,0,57,0,0,0,212,0,149,0,67,0,0,0,0,0,141,0,0,0,130,0,42,0,63,0,134,0,83,0,0,0,153,0,47,0,59,0,19,0,175,0,221,0,95,0,87,0,12,0,168,0,233,0,58,0,36,0,135,0,71,0,217,0,63,0,83,0,241,0,13,0,112,0,80,0,39,0,43,0,0,0,0,0,130,0,124,0,0,0,209,0,112,0,56,0,0,0,189,0,0,0,240,0,116,0,0,0,16,0,0,0,158,0,0,0,0,0,78,0,86,0,229,0,0,0,223,0,232,0,0,0,186,0,0,0,106,0,0,0,131,0,0,0,205,0,0,0,0,0,0,0,190,0,0,0,0,0,45,0,0,0,127,0,161,0,71,0,0,0,199,0,0,0,0,0,5,0,107,0,124,0,3,0,7,0,62,0,2,0,105,0,12,0,241,0,56,0,82,0,214,0,48,0,66,0,11,0,56,0,0,0,0,0,0,0,147,0,151,0,128,0,42,0,226,0,110,0,120,0,202,0,207,0,194,0,0,0,105,0,168,0,232,0,233,0,55,0,0,0,56,0,132,0,247,0,139,0,199,0,210,0,197,0,97,0,0,0,116,0,3,0,28,0,245,0,134,0,38,0,148,0,179,0,105,0,197,0,0,0,35,0,176,0,157,0,102,0,187,0,159,0,183,0,0,0,40,0,238,0,212,0,0,0,0,0,231,0,158,0,112,0,6,0,11,0,92,0,0,0,81,0,175,0,148,0,87,0,141,0,88,0,96,0,193,0,115,0,133,0,21,0,22,0,208,0,151,0,122,0,0,0,4,0,0,0,221,0,0,0,155,0,46,0,0,0,113,0,67,0,252,0,4,0,228,0,196,0,70,0,24,0,85,0,0,0,11,0,136,0,190,0,71,0,0,0,172,0,0,0,0,0,237,0,0,0,38,0,106,0,57,0,229,0,0,0,0,0,0,0,254,0,31,0,220,0,122,0,2,0,151,0,0,0,0,0,131,0,208,0,92,0,157,0,166,0,17,0,0,0,244,0,30,0,2,0,0,0,224,0,0,0,82,0,0,0,158,0,0,0,150,0,11,0,0,0,91,0,142,0,193,0,210,0,154,0,157,0,189,0,0,0,84,0,78,0,30,0,200,0,0,0,0,0,227,0,0,0,214,0,245,0,48,0,121,0,11,0,199,0,0,0,247,0,0,0,127,0,0,0,80,0,227,0,20,0,130,0,42,0,0,0,156,0,97,0,111,0,35,0,213,0,0,0,148,0,35,0,97,0,0,0,176,0,0,0,147,0,0,0,160,0,254,0,34,0,103,0,243,0,133,0,0,0,121,0,148,0,30,0,107,0,40,0,19,0,0,0,0,0,0,0,60,0,252,0,170,0,254,0,81,0,26,0,0,0,0,0,6,0,0,0,65,0,54,0,38,0,0,0,244,0,2,0,248,0,227,0,0,0,81,0,161,0,0,0,0,0,0,0,93,0,228,0,134,0,223,0,255,0,245,0,83,0,83,0,11,0,13,0,247,0,0,0,106,0,0,0,0,0,76,0,160,0,45,0,51,0,124,0,32,0,163,0,121,0,88,0,0,0,115,0,39,0,121,0,205,0,76,0,169,0);
signal scenario_full  : scenario_type := (211,31,164,31,188,31,88,31,88,30,214,31,176,31,32,31,32,30,32,31,164,31,97,31,147,31,147,30,230,31,101,31,110,31,248,31,154,31,122,31,67,31,8,31,217,31,217,30,111,31,203,31,240,31,119,31,92,31,109,31,73,31,180,31,94,31,171,31,171,30,40,31,169,31,182,31,191,31,104,31,67,31,103,31,62,31,59,31,37,31,198,31,145,31,91,31,78,31,146,31,146,30,146,29,70,31,70,30,138,31,242,31,36,31,199,31,81,31,245,31,237,31,120,31,61,31,181,31,235,31,67,31,97,31,97,30,97,29,191,31,27,31,16,31,16,30,16,29,16,28,173,31,15,31,180,31,3,31,3,30,50,31,198,31,55,31,129,31,98,31,89,31,115,31,115,30,115,29,109,31,246,31,167,31,161,31,18,31,195,31,64,31,253,31,253,30,51,31,12,31,58,31,43,31,10,31,39,31,39,30,39,29,104,31,82,31,82,30,151,31,151,30,251,31,249,31,225,31,72,31,190,31,190,30,117,31,197,31,197,30,133,31,53,31,53,30,68,31,117,31,59,31,135,31,159,31,106,31,242,31,138,31,167,31,241,31,151,31,80,31,241,31,246,31,156,31,229,31,9,31,46,31,61,31,49,31,10,31,174,31,36,31,17,31,179,31,166,31,148,31,4,31,137,31,254,31,116,31,226,31,44,31,62,31,62,30,62,29,178,31,109,31,82,31,21,31,21,30,21,29,79,31,72,31,164,31,176,31,74,31,228,31,177,31,230,31,148,31,148,30,247,31,213,31,226,31,132,31,136,31,188,31,112,31,138,31,132,31,132,30,168,31,168,30,135,31,176,31,176,30,28,31,200,31,63,31,252,31,133,31,77,31,223,31,10,31,178,31,91,31,91,30,91,29,137,31,72,31,41,31,217,31,27,31,232,31,79,31,101,31,95,31,241,31,241,30,195,31,99,31,223,31,174,31,171,31,197,31,197,30,18,31,198,31,198,30,174,31,90,31,198,31,198,30,90,31,239,31,69,31,95,31,30,31,37,31,37,30,54,31,236,31,62,31,137,31,137,30,86,31,35,31,103,31,103,30,103,29,103,28,150,31,150,30,150,29,36,31,99,31,229,31,94,31,58,31,58,30,48,31,222,31,222,30,222,29,80,31,218,31,51,31,51,30,230,31,104,31,127,31,251,31,236,31,236,30,5,31,144,31,187,31,56,31,235,31,81,31,81,30,179,31,114,31,114,30,247,31,247,30,11,31,85,31,240,31,68,31,3,31,142,31,158,31,89,31,108,31,108,30,151,31,151,30,151,29,137,31,95,31,183,31,146,31,36,31,82,31,86,31,193,31,10,31,242,31,39,31,202,31,47,31,47,30,47,29,172,31,172,30,246,31,246,30,59,31,71,31,227,31,179,31,22,31,167,31,60,31,242,31,41,31,145,31,11,31,134,31,134,30,57,31,74,31,80,31,80,30,182,31,22,31,98,31,98,30,164,31,128,31,44,31,63,31,213,31,225,31,225,30,225,29,127,31,127,30,182,31,182,30,34,31,34,30,34,29,182,31,42,31,185,31,163,31,163,30,181,31,64,31,134,31,134,30,57,31,9,31,233,31,233,30,212,31,236,31,236,30,207,31,8,31,2,31,136,31,255,31,40,31,133,31,167,31,31,31,146,31,50,31,119,31,233,31,247,31,247,30,28,31,28,30,33,31,231,31,72,31,72,30,72,29,72,28,72,27,127,31,127,30,76,31,124,31,39,31,52,31,72,31,72,30,145,31,18,31,17,31,8,31,168,31,82,31,238,31,86,31,86,30,171,31,171,30,171,29,66,31,138,31,59,31,204,31,21,31,42,31,42,30,150,31,150,30,57,31,228,31,100,31,100,30,41,31,78,31,10,31,141,31,141,30,152,31,98,31,98,30,157,31,92,31,92,30,82,31,82,30,129,31,81,31,31,31,255,31,29,31,62,31,62,30,57,31,57,30,212,31,149,31,67,31,67,30,67,29,141,31,141,30,130,31,42,31,63,31,134,31,83,31,83,30,153,31,47,31,59,31,19,31,175,31,221,31,95,31,87,31,12,31,168,31,233,31,58,31,36,31,135,31,71,31,217,31,63,31,83,31,241,31,13,31,112,31,80,31,39,31,43,31,43,30,43,29,130,31,124,31,124,30,209,31,112,31,56,31,56,30,189,31,189,30,240,31,116,31,116,30,16,31,16,30,158,31,158,30,158,29,78,31,86,31,229,31,229,30,223,31,232,31,232,30,186,31,186,30,106,31,106,30,131,31,131,30,205,31,205,30,205,29,205,28,190,31,190,30,190,29,45,31,45,30,127,31,161,31,71,31,71,30,199,31,199,30,199,29,5,31,107,31,124,31,3,31,7,31,62,31,2,31,105,31,12,31,241,31,56,31,82,31,214,31,48,31,66,31,11,31,56,31,56,30,56,29,56,28,147,31,151,31,128,31,42,31,226,31,110,31,120,31,202,31,207,31,194,31,194,30,105,31,168,31,232,31,233,31,55,31,55,30,56,31,132,31,247,31,139,31,199,31,210,31,197,31,97,31,97,30,116,31,3,31,28,31,245,31,134,31,38,31,148,31,179,31,105,31,197,31,197,30,35,31,176,31,157,31,102,31,187,31,159,31,183,31,183,30,40,31,238,31,212,31,212,30,212,29,231,31,158,31,112,31,6,31,11,31,92,31,92,30,81,31,175,31,148,31,87,31,141,31,88,31,96,31,193,31,115,31,133,31,21,31,22,31,208,31,151,31,122,31,122,30,4,31,4,30,221,31,221,30,155,31,46,31,46,30,113,31,67,31,252,31,4,31,228,31,196,31,70,31,24,31,85,31,85,30,11,31,136,31,190,31,71,31,71,30,172,31,172,30,172,29,237,31,237,30,38,31,106,31,57,31,229,31,229,30,229,29,229,28,254,31,31,31,220,31,122,31,2,31,151,31,151,30,151,29,131,31,208,31,92,31,157,31,166,31,17,31,17,30,244,31,30,31,2,31,2,30,224,31,224,30,82,31,82,30,158,31,158,30,150,31,11,31,11,30,91,31,142,31,193,31,210,31,154,31,157,31,189,31,189,30,84,31,78,31,30,31,200,31,200,30,200,29,227,31,227,30,214,31,245,31,48,31,121,31,11,31,199,31,199,30,247,31,247,30,127,31,127,30,80,31,227,31,20,31,130,31,42,31,42,30,156,31,97,31,111,31,35,31,213,31,213,30,148,31,35,31,97,31,97,30,176,31,176,30,147,31,147,30,160,31,254,31,34,31,103,31,243,31,133,31,133,30,121,31,148,31,30,31,107,31,40,31,19,31,19,30,19,29,19,28,60,31,252,31,170,31,254,31,81,31,26,31,26,30,26,29,6,31,6,30,65,31,54,31,38,31,38,30,244,31,2,31,248,31,227,31,227,30,81,31,161,31,161,30,161,29,161,28,93,31,228,31,134,31,223,31,255,31,245,31,83,31,83,31,11,31,13,31,247,31,247,30,106,31,106,30,106,29,76,31,160,31,45,31,51,31,124,31,32,31,163,31,121,31,88,31,88,30,115,31,39,31,121,31,205,31,76,31,169,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
