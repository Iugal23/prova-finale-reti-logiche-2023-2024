-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 361;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (148,0,33,0,0,0,62,0,124,0,158,0,253,0,242,0,153,0,0,0,12,0,197,0,195,0,91,0,0,0,223,0,0,0,56,0,176,0,0,0,41,0,0,0,85,0,85,0,85,0,225,0,191,0,179,0,21,0,216,0,51,0,0,0,151,0,236,0,141,0,48,0,0,0,112,0,235,0,114,0,0,0,65,0,61,0,253,0,206,0,0,0,47,0,0,0,57,0,84,0,39,0,0,0,225,0,86,0,108,0,18,0,0,0,94,0,167,0,192,0,103,0,45,0,76,0,86,0,43,0,13,0,86,0,95,0,0,0,226,0,0,0,215,0,65,0,0,0,0,0,20,0,156,0,0,0,0,0,14,0,0,0,47,0,149,0,25,0,155,0,66,0,0,0,245,0,234,0,218,0,30,0,59,0,168,0,0,0,128,0,0,0,4,0,109,0,120,0,0,0,0,0,121,0,129,0,203,0,138,0,0,0,248,0,107,0,62,0,116,0,93,0,207,0,96,0,180,0,183,0,174,0,92,0,116,0,20,0,118,0,104,0,151,0,0,0,188,0,0,0,176,0,0,0,210,0,10,0,4,0,54,0,27,0,11,0,10,0,48,0,162,0,48,0,0,0,54,0,173,0,86,0,51,0,0,0,89,0,136,0,20,0,62,0,0,0,66,0,27,0,182,0,204,0,56,0,219,0,165,0,0,0,243,0,92,0,241,0,159,0,0,0,188,0,0,0,201,0,77,0,185,0,145,0,203,0,169,0,231,0,32,0,222,0,0,0,110,0,112,0,77,0,16,0,0,0,203,0,0,0,213,0,236,0,249,0,197,0,232,0,160,0,245,0,217,0,120,0,89,0,112,0,0,0,208,0,91,0,119,0,81,0,83,0,136,0,190,0,104,0,67,0,223,0,165,0,45,0,218,0,29,0,120,0,56,0,58,0,11,0,226,0,150,0,232,0,18,0,201,0,177,0,55,0,0,0,0,0,212,0,243,0,249,0,0,0,0,0,212,0,0,0,135,0,0,0,163,0,251,0,0,0,206,0,183,0,6,0,44,0,0,0,194,0,240,0,137,0,120,0,0,0,215,0,0,0,18,0,179,0,0,0,215,0,183,0,0,0,11,0,10,0,202,0,46,0,0,0,88,0,122,0,177,0,154,0,198,0,123,0,230,0,175,0,232,0,1,0,0,0,74,0,20,0,0,0,135,0,238,0,159,0,61,0,0,0,0,0,90,0,63,0,75,0,240,0,192,0,118,0,0,0,49,0,66,0,130,0,249,0,157,0,0,0,60,0,0,0,191,0,103,0,0,0,59,0,0,0,55,0,113,0,244,0,176,0,136,0,204,0,225,0,0,0,40,0,156,0,96,0,31,0,225,0,0,0,196,0,168,0,182,0,0,0,0,0,98,0,154,0,0,0,3,0,252,0,222,0,0,0,197,0,0,0,204,0,229,0,145,0,0,0,40,0,0,0,0,0,87,0,209,0,177,0,0,0,184,0,22,0,71,0,5,0,21,0,154,0,246,0,30,0,0,0,0,0,0,0,0,0,69,0,161,0,0,0,0,0,146,0,0,0,184,0,0,0,162,0,66,0,135,0,148,0,43,0,172,0,0,0,33,0);
signal scenario_full  : scenario_type := (148,31,33,31,33,30,62,31,124,31,158,31,253,31,242,31,153,31,153,30,12,31,197,31,195,31,91,31,91,30,223,31,223,30,56,31,176,31,176,30,41,31,41,30,85,31,85,31,85,31,225,31,191,31,179,31,21,31,216,31,51,31,51,30,151,31,236,31,141,31,48,31,48,30,112,31,235,31,114,31,114,30,65,31,61,31,253,31,206,31,206,30,47,31,47,30,57,31,84,31,39,31,39,30,225,31,86,31,108,31,18,31,18,30,94,31,167,31,192,31,103,31,45,31,76,31,86,31,43,31,13,31,86,31,95,31,95,30,226,31,226,30,215,31,65,31,65,30,65,29,20,31,156,31,156,30,156,29,14,31,14,30,47,31,149,31,25,31,155,31,66,31,66,30,245,31,234,31,218,31,30,31,59,31,168,31,168,30,128,31,128,30,4,31,109,31,120,31,120,30,120,29,121,31,129,31,203,31,138,31,138,30,248,31,107,31,62,31,116,31,93,31,207,31,96,31,180,31,183,31,174,31,92,31,116,31,20,31,118,31,104,31,151,31,151,30,188,31,188,30,176,31,176,30,210,31,10,31,4,31,54,31,27,31,11,31,10,31,48,31,162,31,48,31,48,30,54,31,173,31,86,31,51,31,51,30,89,31,136,31,20,31,62,31,62,30,66,31,27,31,182,31,204,31,56,31,219,31,165,31,165,30,243,31,92,31,241,31,159,31,159,30,188,31,188,30,201,31,77,31,185,31,145,31,203,31,169,31,231,31,32,31,222,31,222,30,110,31,112,31,77,31,16,31,16,30,203,31,203,30,213,31,236,31,249,31,197,31,232,31,160,31,245,31,217,31,120,31,89,31,112,31,112,30,208,31,91,31,119,31,81,31,83,31,136,31,190,31,104,31,67,31,223,31,165,31,45,31,218,31,29,31,120,31,56,31,58,31,11,31,226,31,150,31,232,31,18,31,201,31,177,31,55,31,55,30,55,29,212,31,243,31,249,31,249,30,249,29,212,31,212,30,135,31,135,30,163,31,251,31,251,30,206,31,183,31,6,31,44,31,44,30,194,31,240,31,137,31,120,31,120,30,215,31,215,30,18,31,179,31,179,30,215,31,183,31,183,30,11,31,10,31,202,31,46,31,46,30,88,31,122,31,177,31,154,31,198,31,123,31,230,31,175,31,232,31,1,31,1,30,74,31,20,31,20,30,135,31,238,31,159,31,61,31,61,30,61,29,90,31,63,31,75,31,240,31,192,31,118,31,118,30,49,31,66,31,130,31,249,31,157,31,157,30,60,31,60,30,191,31,103,31,103,30,59,31,59,30,55,31,113,31,244,31,176,31,136,31,204,31,225,31,225,30,40,31,156,31,96,31,31,31,225,31,225,30,196,31,168,31,182,31,182,30,182,29,98,31,154,31,154,30,3,31,252,31,222,31,222,30,197,31,197,30,204,31,229,31,145,31,145,30,40,31,40,30,40,29,87,31,209,31,177,31,177,30,184,31,22,31,71,31,5,31,21,31,154,31,246,31,30,31,30,30,30,29,30,28,30,27,69,31,161,31,161,30,161,29,146,31,146,30,184,31,184,30,162,31,66,31,135,31,148,31,43,31,172,31,172,30,33,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
