-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_201 is
end project_tb_201;

architecture project_tb_arch_201 of project_tb_201 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 295;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (160,0,33,0,193,0,107,0,77,0,136,0,253,0,163,0,171,0,227,0,169,0,161,0,53,0,0,0,0,0,7,0,167,0,198,0,205,0,35,0,88,0,207,0,0,0,185,0,85,0,0,0,180,0,48,0,218,0,74,0,149,0,0,0,59,0,163,0,186,0,114,0,0,0,0,0,5,0,0,0,112,0,152,0,146,0,197,0,40,0,173,0,0,0,92,0,64,0,86,0,255,0,0,0,194,0,26,0,0,0,208,0,0,0,71,0,226,0,58,0,0,0,0,0,243,0,248,0,178,0,0,0,243,0,236,0,7,0,151,0,192,0,109,0,80,0,0,0,204,0,171,0,190,0,0,0,214,0,178,0,68,0,215,0,148,0,35,0,46,0,88,0,217,0,28,0,54,0,243,0,221,0,41,0,199,0,68,0,127,0,0,0,0,0,210,0,226,0,152,0,43,0,157,0,2,0,0,0,25,0,21,0,135,0,0,0,222,0,39,0,85,0,15,0,3,0,95,0,5,0,216,0,0,0,70,0,248,0,102,0,218,0,178,0,27,0,143,0,68,0,0,0,85,0,134,0,255,0,0,0,228,0,238,0,159,0,71,0,186,0,9,0,121,0,0,0,138,0,22,0,187,0,64,0,146,0,102,0,176,0,132,0,4,0,0,0,35,0,230,0,177,0,58,0,108,0,225,0,233,0,162,0,0,0,230,0,230,0,136,0,18,0,81,0,50,0,231,0,196,0,211,0,122,0,21,0,82,0,194,0,187,0,216,0,0,0,236,0,0,0,0,0,194,0,11,0,16,0,0,0,43,0,203,0,100,0,235,0,123,0,85,0,122,0,193,0,0,0,0,0,222,0,0,0,94,0,209,0,98,0,72,0,240,0,49,0,137,0,178,0,0,0,154,0,252,0,13,0,110,0,3,0,0,0,71,0,30,0,245,0,199,0,234,0,148,0,153,0,100,0,149,0,202,0,246,0,47,0,119,0,119,0,226,0,251,0,0,0,234,0,95,0,0,0,241,0,158,0,177,0,0,0,119,0,0,0,5,0,169,0,133,0,21,0,0,0,0,0,64,0,214,0,0,0,61,0,221,0,130,0,85,0,160,0,102,0,167,0,239,0,122,0,183,0,211,0,170,0,87,0,215,0,0,0,172,0,207,0,16,0,171,0,28,0,242,0,217,0,72,0,109,0,26,0,28,0,71,0,0,0,125,0,158,0,176,0,120,0,140,0,142,0,139,0,232,0,5,0,0,0,59,0,0,0,0,0,0,0,116,0,38,0,0,0,16,0,125,0,135,0,0,0,24,0,6,0,35,0,53,0);
signal scenario_full  : scenario_type := (160,31,33,31,193,31,107,31,77,31,136,31,253,31,163,31,171,31,227,31,169,31,161,31,53,31,53,30,53,29,7,31,167,31,198,31,205,31,35,31,88,31,207,31,207,30,185,31,85,31,85,30,180,31,48,31,218,31,74,31,149,31,149,30,59,31,163,31,186,31,114,31,114,30,114,29,5,31,5,30,112,31,152,31,146,31,197,31,40,31,173,31,173,30,92,31,64,31,86,31,255,31,255,30,194,31,26,31,26,30,208,31,208,30,71,31,226,31,58,31,58,30,58,29,243,31,248,31,178,31,178,30,243,31,236,31,7,31,151,31,192,31,109,31,80,31,80,30,204,31,171,31,190,31,190,30,214,31,178,31,68,31,215,31,148,31,35,31,46,31,88,31,217,31,28,31,54,31,243,31,221,31,41,31,199,31,68,31,127,31,127,30,127,29,210,31,226,31,152,31,43,31,157,31,2,31,2,30,25,31,21,31,135,31,135,30,222,31,39,31,85,31,15,31,3,31,95,31,5,31,216,31,216,30,70,31,248,31,102,31,218,31,178,31,27,31,143,31,68,31,68,30,85,31,134,31,255,31,255,30,228,31,238,31,159,31,71,31,186,31,9,31,121,31,121,30,138,31,22,31,187,31,64,31,146,31,102,31,176,31,132,31,4,31,4,30,35,31,230,31,177,31,58,31,108,31,225,31,233,31,162,31,162,30,230,31,230,31,136,31,18,31,81,31,50,31,231,31,196,31,211,31,122,31,21,31,82,31,194,31,187,31,216,31,216,30,236,31,236,30,236,29,194,31,11,31,16,31,16,30,43,31,203,31,100,31,235,31,123,31,85,31,122,31,193,31,193,30,193,29,222,31,222,30,94,31,209,31,98,31,72,31,240,31,49,31,137,31,178,31,178,30,154,31,252,31,13,31,110,31,3,31,3,30,71,31,30,31,245,31,199,31,234,31,148,31,153,31,100,31,149,31,202,31,246,31,47,31,119,31,119,31,226,31,251,31,251,30,234,31,95,31,95,30,241,31,158,31,177,31,177,30,119,31,119,30,5,31,169,31,133,31,21,31,21,30,21,29,64,31,214,31,214,30,61,31,221,31,130,31,85,31,160,31,102,31,167,31,239,31,122,31,183,31,211,31,170,31,87,31,215,31,215,30,172,31,207,31,16,31,171,31,28,31,242,31,217,31,72,31,109,31,26,31,28,31,71,31,71,30,125,31,158,31,176,31,120,31,140,31,142,31,139,31,232,31,5,31,5,30,59,31,59,30,59,29,59,28,116,31,38,31,38,30,16,31,125,31,135,31,135,30,24,31,6,31,35,31,53,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
