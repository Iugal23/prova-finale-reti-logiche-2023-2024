-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_912 is
end project_tb_912;

architecture project_tb_arch_912 of project_tb_912 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 821;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (11,0,30,0,84,0,8,0,4,0,18,0,75,0,18,0,75,0,80,0,167,0,74,0,0,0,122,0,220,0,46,0,203,0,82,0,172,0,196,0,145,0,142,0,92,0,59,0,130,0,247,0,5,0,108,0,34,0,157,0,99,0,0,0,158,0,0,0,0,0,207,0,53,0,0,0,0,0,0,0,0,0,200,0,175,0,142,0,158,0,0,0,0,0,78,0,243,0,191,0,5,0,121,0,216,0,46,0,0,0,35,0,0,0,155,0,230,0,0,0,209,0,10,0,208,0,117,0,64,0,155,0,0,0,220,0,234,0,0,0,11,0,220,0,144,0,83,0,235,0,18,0,53,0,37,0,249,0,195,0,143,0,0,0,179,0,0,0,6,0,147,0,231,0,150,0,224,0,212,0,0,0,111,0,56,0,200,0,0,0,124,0,223,0,230,0,0,0,248,0,0,0,147,0,130,0,188,0,113,0,171,0,0,0,157,0,216,0,0,0,236,0,164,0,0,0,168,0,0,0,119,0,96,0,33,0,133,0,0,0,0,0,0,0,113,0,154,0,59,0,0,0,204,0,15,0,251,0,109,0,38,0,15,0,92,0,0,0,241,0,123,0,217,0,177,0,0,0,0,0,176,0,27,0,220,0,136,0,2,0,0,0,113,0,229,0,155,0,252,0,229,0,156,0,48,0,113,0,99,0,77,0,231,0,123,0,20,0,78,0,25,0,0,0,241,0,0,0,0,0,198,0,0,0,140,0,47,0,12,0,24,0,0,0,86,0,56,0,0,0,13,0,146,0,77,0,192,0,129,0,26,0,202,0,217,0,26,0,80,0,149,0,2,0,0,0,26,0,41,0,141,0,148,0,196,0,132,0,198,0,77,0,199,0,0,0,178,0,214,0,143,0,0,0,122,0,0,0,37,0,0,0,117,0,210,0,0,0,245,0,240,0,161,0,242,0,251,0,14,0,56,0,141,0,0,0,35,0,13,0,79,0,15,0,92,0,243,0,100,0,192,0,225,0,8,0,6,0,121,0,38,0,0,0,0,0,0,0,202,0,29,0,213,0,0,0,255,0,0,0,0,0,213,0,0,0,60,0,213,0,184,0,48,0,0,0,0,0,0,0,0,0,0,0,242,0,90,0,0,0,0,0,164,0,12,0,0,0,120,0,107,0,0,0,109,0,60,0,0,0,0,0,3,0,241,0,35,0,0,0,0,0,70,0,70,0,230,0,19,0,0,0,104,0,247,0,176,0,25,0,0,0,128,0,139,0,132,0,0,0,239,0,76,0,200,0,0,0,210,0,139,0,51,0,0,0,242,0,60,0,103,0,142,0,114,0,105,0,17,0,226,0,87,0,114,0,141,0,0,0,38,0,174,0,167,0,93,0,90,0,130,0,53,0,35,0,135,0,133,0,0,0,3,0,168,0,164,0,43,0,208,0,120,0,231,0,79,0,230,0,16,0,0,0,211,0,230,0,64,0,111,0,8,0,0,0,204,0,138,0,78,0,0,0,200,0,28,0,144,0,89,0,0,0,70,0,193,0,77,0,196,0,38,0,0,0,109,0,217,0,76,0,0,0,33,0,197,0,70,0,36,0,80,0,194,0,50,0,244,0,0,0,39,0,0,0,20,0,40,0,83,0,114,0,130,0,0,0,194,0,39,0,203,0,0,0,0,0,4,0,0,0,0,0,147,0,223,0,0,0,0,0,10,0,49,0,0,0,247,0,93,0,11,0,117,0,239,0,197,0,241,0,219,0,0,0,185,0,0,0,165,0,0,0,72,0,0,0,213,0,61,0,0,0,123,0,83,0,103,0,96,0,33,0,0,0,0,0,94,0,14,0,239,0,159,0,0,0,31,0,11,0,190,0,102,0,176,0,0,0,238,0,0,0,119,0,211,0,9,0,16,0,97,0,190,0,120,0,172,0,22,0,142,0,0,0,37,0,0,0,255,0,211,0,166,0,101,0,117,0,0,0,0,0,127,0,185,0,0,0,18,0,12,0,183,0,131,0,77,0,203,0,0,0,197,0,235,0,254,0,37,0,103,0,132,0,152,0,206,0,212,0,48,0,181,0,0,0,121,0,0,0,61,0,121,0,45,0,108,0,199,0,163,0,0,0,0,0,159,0,127,0,148,0,180,0,99,0,0,0,129,0,22,0,236,0,19,0,149,0,189,0,74,0,3,0,0,0,0,0,0,0,204,0,99,0,136,0,103,0,0,0,120,0,148,0,100,0,78,0,0,0,12,0,196,0,150,0,201,0,106,0,8,0,181,0,151,0,71,0,169,0,141,0,240,0,59,0,16,0,165,0,70,0,47,0,70,0,31,0,250,0,118,0,196,0,50,0,205,0,184,0,44,0,21,0,0,0,43,0,12,0,234,0,78,0,255,0,230,0,80,0,158,0,26,0,0,0,0,0,0,0,0,0,249,0,19,0,239,0,0,0,136,0,232,0,70,0,74,0,215,0,255,0,108,0,0,0,85,0,110,0,8,0,252,0,76,0,89,0,38,0,105,0,0,0,169,0,69,0,0,0,0,0,178,0,0,0,47,0,0,0,157,0,100,0,0,0,100,0,95,0,178,0,171,0,64,0,28,0,0,0,248,0,5,0,248,0,47,0,215,0,16,0,192,0,87,0,29,0,144,0,99,0,42,0,91,0,0,0,0,0,120,0,26,0,0,0,181,0,69,0,137,0,57,0,14,0,57,0,79,0,0,0,23,0,61,0,40,0,120,0,170,0,94,0,114,0,225,0,215,0,254,0,66,0,48,0,176,0,0,0,201,0,150,0,120,0,248,0,106,0,145,0,194,0,0,0,0,0,0,0,0,0,43,0,35,0,96,0,0,0,156,0,92,0,88,0,83,0,0,0,231,0,173,0,0,0,127,0,142,0,155,0,76,0,182,0,127,0,195,0,232,0,158,0,153,0,0,0,163,0,62,0,220,0,229,0,69,0,33,0,0,0,168,0,108,0,238,0,253,0,209,0,20,0,100,0,50,0,5,0,2,0,68,0,214,0,133,0,0,0,0,0,74,0,230,0,0,0,66,0,0,0,135,0,96,0,7,0,162,0,32,0,39,0,0,0,36,0,147,0,211,0,0,0,81,0,145,0,0,0,34,0,0,0,155,0,213,0,168,0,6,0,81,0,43,0,197,0,199,0,139,0,157,0,39,0,112,0,94,0,95,0,80,0,243,0,150,0,160,0,229,0,0,0,231,0,0,0,108,0,149,0,30,0,19,0,250,0,152,0,20,0,34,0,92,0,203,0,237,0,72,0,32,0,228,0,72,0,0,0,51,0,109,0,132,0,0,0,151,0,128,0,168,0,0,0,207,0,145,0,183,0,238,0,0,0,72,0,57,0,243,0,0,0,0,0,25,0,5,0,157,0,237,0,35,0,169,0,106,0,199,0,111,0,55,0,17,0,181,0,0,0,187,0,0,0,50,0,144,0,0,0,172,0,230,0,85,0,143,0,0,0,121,0,250,0,17,0,225,0,12,0,158,0,236,0,0,0,235,0,22,0,243,0,0,0,106,0,0,0,197,0,28,0,199,0,0,0,143,0,113,0,0,0,0,0,105,0,0,0,216,0,0,0,146,0,57,0,255,0,64,0,0,0,25,0,55,0,0,0,30,0,33,0,181,0,178,0,111,0,251,0,143,0,0,0,0,0,0,0);
signal scenario_full  : scenario_type := (11,31,30,31,84,31,8,31,4,31,18,31,75,31,18,31,75,31,80,31,167,31,74,31,74,30,122,31,220,31,46,31,203,31,82,31,172,31,196,31,145,31,142,31,92,31,59,31,130,31,247,31,5,31,108,31,34,31,157,31,99,31,99,30,158,31,158,30,158,29,207,31,53,31,53,30,53,29,53,28,53,27,200,31,175,31,142,31,158,31,158,30,158,29,78,31,243,31,191,31,5,31,121,31,216,31,46,31,46,30,35,31,35,30,155,31,230,31,230,30,209,31,10,31,208,31,117,31,64,31,155,31,155,30,220,31,234,31,234,30,11,31,220,31,144,31,83,31,235,31,18,31,53,31,37,31,249,31,195,31,143,31,143,30,179,31,179,30,6,31,147,31,231,31,150,31,224,31,212,31,212,30,111,31,56,31,200,31,200,30,124,31,223,31,230,31,230,30,248,31,248,30,147,31,130,31,188,31,113,31,171,31,171,30,157,31,216,31,216,30,236,31,164,31,164,30,168,31,168,30,119,31,96,31,33,31,133,31,133,30,133,29,133,28,113,31,154,31,59,31,59,30,204,31,15,31,251,31,109,31,38,31,15,31,92,31,92,30,241,31,123,31,217,31,177,31,177,30,177,29,176,31,27,31,220,31,136,31,2,31,2,30,113,31,229,31,155,31,252,31,229,31,156,31,48,31,113,31,99,31,77,31,231,31,123,31,20,31,78,31,25,31,25,30,241,31,241,30,241,29,198,31,198,30,140,31,47,31,12,31,24,31,24,30,86,31,56,31,56,30,13,31,146,31,77,31,192,31,129,31,26,31,202,31,217,31,26,31,80,31,149,31,2,31,2,30,26,31,41,31,141,31,148,31,196,31,132,31,198,31,77,31,199,31,199,30,178,31,214,31,143,31,143,30,122,31,122,30,37,31,37,30,117,31,210,31,210,30,245,31,240,31,161,31,242,31,251,31,14,31,56,31,141,31,141,30,35,31,13,31,79,31,15,31,92,31,243,31,100,31,192,31,225,31,8,31,6,31,121,31,38,31,38,30,38,29,38,28,202,31,29,31,213,31,213,30,255,31,255,30,255,29,213,31,213,30,60,31,213,31,184,31,48,31,48,30,48,29,48,28,48,27,48,26,242,31,90,31,90,30,90,29,164,31,12,31,12,30,120,31,107,31,107,30,109,31,60,31,60,30,60,29,3,31,241,31,35,31,35,30,35,29,70,31,70,31,230,31,19,31,19,30,104,31,247,31,176,31,25,31,25,30,128,31,139,31,132,31,132,30,239,31,76,31,200,31,200,30,210,31,139,31,51,31,51,30,242,31,60,31,103,31,142,31,114,31,105,31,17,31,226,31,87,31,114,31,141,31,141,30,38,31,174,31,167,31,93,31,90,31,130,31,53,31,35,31,135,31,133,31,133,30,3,31,168,31,164,31,43,31,208,31,120,31,231,31,79,31,230,31,16,31,16,30,211,31,230,31,64,31,111,31,8,31,8,30,204,31,138,31,78,31,78,30,200,31,28,31,144,31,89,31,89,30,70,31,193,31,77,31,196,31,38,31,38,30,109,31,217,31,76,31,76,30,33,31,197,31,70,31,36,31,80,31,194,31,50,31,244,31,244,30,39,31,39,30,20,31,40,31,83,31,114,31,130,31,130,30,194,31,39,31,203,31,203,30,203,29,4,31,4,30,4,29,147,31,223,31,223,30,223,29,10,31,49,31,49,30,247,31,93,31,11,31,117,31,239,31,197,31,241,31,219,31,219,30,185,31,185,30,165,31,165,30,72,31,72,30,213,31,61,31,61,30,123,31,83,31,103,31,96,31,33,31,33,30,33,29,94,31,14,31,239,31,159,31,159,30,31,31,11,31,190,31,102,31,176,31,176,30,238,31,238,30,119,31,211,31,9,31,16,31,97,31,190,31,120,31,172,31,22,31,142,31,142,30,37,31,37,30,255,31,211,31,166,31,101,31,117,31,117,30,117,29,127,31,185,31,185,30,18,31,12,31,183,31,131,31,77,31,203,31,203,30,197,31,235,31,254,31,37,31,103,31,132,31,152,31,206,31,212,31,48,31,181,31,181,30,121,31,121,30,61,31,121,31,45,31,108,31,199,31,163,31,163,30,163,29,159,31,127,31,148,31,180,31,99,31,99,30,129,31,22,31,236,31,19,31,149,31,189,31,74,31,3,31,3,30,3,29,3,28,204,31,99,31,136,31,103,31,103,30,120,31,148,31,100,31,78,31,78,30,12,31,196,31,150,31,201,31,106,31,8,31,181,31,151,31,71,31,169,31,141,31,240,31,59,31,16,31,165,31,70,31,47,31,70,31,31,31,250,31,118,31,196,31,50,31,205,31,184,31,44,31,21,31,21,30,43,31,12,31,234,31,78,31,255,31,230,31,80,31,158,31,26,31,26,30,26,29,26,28,26,27,249,31,19,31,239,31,239,30,136,31,232,31,70,31,74,31,215,31,255,31,108,31,108,30,85,31,110,31,8,31,252,31,76,31,89,31,38,31,105,31,105,30,169,31,69,31,69,30,69,29,178,31,178,30,47,31,47,30,157,31,100,31,100,30,100,31,95,31,178,31,171,31,64,31,28,31,28,30,248,31,5,31,248,31,47,31,215,31,16,31,192,31,87,31,29,31,144,31,99,31,42,31,91,31,91,30,91,29,120,31,26,31,26,30,181,31,69,31,137,31,57,31,14,31,57,31,79,31,79,30,23,31,61,31,40,31,120,31,170,31,94,31,114,31,225,31,215,31,254,31,66,31,48,31,176,31,176,30,201,31,150,31,120,31,248,31,106,31,145,31,194,31,194,30,194,29,194,28,194,27,43,31,35,31,96,31,96,30,156,31,92,31,88,31,83,31,83,30,231,31,173,31,173,30,127,31,142,31,155,31,76,31,182,31,127,31,195,31,232,31,158,31,153,31,153,30,163,31,62,31,220,31,229,31,69,31,33,31,33,30,168,31,108,31,238,31,253,31,209,31,20,31,100,31,50,31,5,31,2,31,68,31,214,31,133,31,133,30,133,29,74,31,230,31,230,30,66,31,66,30,135,31,96,31,7,31,162,31,32,31,39,31,39,30,36,31,147,31,211,31,211,30,81,31,145,31,145,30,34,31,34,30,155,31,213,31,168,31,6,31,81,31,43,31,197,31,199,31,139,31,157,31,39,31,112,31,94,31,95,31,80,31,243,31,150,31,160,31,229,31,229,30,231,31,231,30,108,31,149,31,30,31,19,31,250,31,152,31,20,31,34,31,92,31,203,31,237,31,72,31,32,31,228,31,72,31,72,30,51,31,109,31,132,31,132,30,151,31,128,31,168,31,168,30,207,31,145,31,183,31,238,31,238,30,72,31,57,31,243,31,243,30,243,29,25,31,5,31,157,31,237,31,35,31,169,31,106,31,199,31,111,31,55,31,17,31,181,31,181,30,187,31,187,30,50,31,144,31,144,30,172,31,230,31,85,31,143,31,143,30,121,31,250,31,17,31,225,31,12,31,158,31,236,31,236,30,235,31,22,31,243,31,243,30,106,31,106,30,197,31,28,31,199,31,199,30,143,31,113,31,113,30,113,29,105,31,105,30,216,31,216,30,146,31,57,31,255,31,64,31,64,30,25,31,55,31,55,30,30,31,33,31,181,31,178,31,111,31,251,31,143,31,143,30,143,29,143,28);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
