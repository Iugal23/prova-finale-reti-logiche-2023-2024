-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 441;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (115,0,0,0,120,0,57,0,185,0,0,0,120,0,209,0,123,0,215,0,0,0,49,0,0,0,95,0,83,0,0,0,49,0,52,0,154,0,0,0,205,0,224,0,0,0,0,0,207,0,194,0,252,0,205,0,51,0,218,0,0,0,0,0,12,0,222,0,85,0,196,0,0,0,0,0,243,0,111,0,51,0,254,0,0,0,72,0,27,0,212,0,0,0,65,0,0,0,14,0,0,0,59,0,57,0,82,0,0,0,0,0,51,0,0,0,66,0,234,0,23,0,107,0,17,0,254,0,33,0,1,0,131,0,0,0,0,0,37,0,90,0,90,0,111,0,245,0,160,0,41,0,3,0,0,0,81,0,107,0,56,0,0,0,46,0,250,0,214,0,8,0,0,0,0,0,200,0,189,0,92,0,121,0,251,0,0,0,0,0,0,0,0,0,67,0,119,0,219,0,41,0,81,0,40,0,30,0,71,0,15,0,119,0,98,0,0,0,51,0,198,0,41,0,158,0,183,0,97,0,0,0,201,0,84,0,231,0,0,0,46,0,77,0,100,0,0,0,180,0,55,0,81,0,251,0,207,0,0,0,92,0,117,0,153,0,138,0,152,0,28,0,95,0,47,0,126,0,249,0,49,0,88,0,22,0,6,0,85,0,45,0,165,0,66,0,0,0,68,0,234,0,214,0,0,0,0,0,124,0,0,0,185,0,126,0,182,0,137,0,196,0,122,0,24,0,0,0,182,0,217,0,0,0,0,0,222,0,42,0,137,0,4,0,135,0,98,0,241,0,191,0,168,0,0,0,37,0,39,0,100,0,0,0,197,0,217,0,187,0,0,0,207,0,203,0,149,0,0,0,125,0,0,0,127,0,193,0,172,0,240,0,0,0,0,0,71,0,218,0,0,0,0,0,108,0,176,0,138,0,159,0,6,0,94,0,126,0,76,0,8,0,52,0,15,0,0,0,0,0,0,0,45,0,130,0,130,0,196,0,79,0,0,0,218,0,0,0,160,0,195,0,0,0,103,0,0,0,49,0,191,0,152,0,101,0,148,0,215,0,180,0,223,0,236,0,0,0,160,0,144,0,0,0,182,0,0,0,130,0,0,0,235,0,135,0,209,0,13,0,11,0,0,0,0,0,43,0,0,0,0,0,105,0,126,0,33,0,134,0,92,0,73,0,211,0,253,0,97,0,0,0,253,0,168,0,122,0,137,0,138,0,0,0,0,0,222,0,133,0,83,0,86,0,80,0,65,0,226,0,28,0,181,0,240,0,233,0,0,0,79,0,0,0,98,0,0,0,107,0,0,0,100,0,197,0,102,0,210,0,0,0,119,0,0,0,174,0,21,0,184,0,108,0,197,0,197,0,185,0,151,0,58,0,169,0,88,0,103,0,162,0,123,0,78,0,129,0,192,0,25,0,213,0,137,0,71,0,54,0,146,0,252,0,0,0,44,0,228,0,83,0,246,0,53,0,0,0,187,0,4,0,165,0,0,0,218,0,139,0,198,0,123,0,44,0,19,0,63,0,150,0,51,0,144,0,154,0,175,0,0,0,7,0,222,0,155,0,21,0,240,0,28,0,0,0,51,0,113,0,112,0,0,0,77,0,12,0,25,0,203,0,155,0,87,0,23,0,166,0,52,0,227,0,63,0,184,0,47,0,0,0,241,0,82,0,0,0,150,0,0,0,97,0,58,0,230,0,29,0,223,0,0,0,38,0,0,0,7,0,3,0,119,0,42,0,165,0,0,0,176,0,59,0,0,0,0,0,239,0,43,0,58,0,120,0,139,0,185,0,38,0,168,0,127,0,0,0,103,0,157,0,0,0,88,0,115,0,76,0,101,0,182,0,0,0,196,0,235,0,0,0,9,0,0,0,0,0,0,0,177,0,12,0,146,0,81,0,0,0,211,0,77,0,203,0,163,0,42,0,30,0,253,0,11,0,118,0,203,0,0,0,180,0,232,0,0,0,80,0,0,0);
signal scenario_full  : scenario_type := (115,31,115,30,120,31,57,31,185,31,185,30,120,31,209,31,123,31,215,31,215,30,49,31,49,30,95,31,83,31,83,30,49,31,52,31,154,31,154,30,205,31,224,31,224,30,224,29,207,31,194,31,252,31,205,31,51,31,218,31,218,30,218,29,12,31,222,31,85,31,196,31,196,30,196,29,243,31,111,31,51,31,254,31,254,30,72,31,27,31,212,31,212,30,65,31,65,30,14,31,14,30,59,31,57,31,82,31,82,30,82,29,51,31,51,30,66,31,234,31,23,31,107,31,17,31,254,31,33,31,1,31,131,31,131,30,131,29,37,31,90,31,90,31,111,31,245,31,160,31,41,31,3,31,3,30,81,31,107,31,56,31,56,30,46,31,250,31,214,31,8,31,8,30,8,29,200,31,189,31,92,31,121,31,251,31,251,30,251,29,251,28,251,27,67,31,119,31,219,31,41,31,81,31,40,31,30,31,71,31,15,31,119,31,98,31,98,30,51,31,198,31,41,31,158,31,183,31,97,31,97,30,201,31,84,31,231,31,231,30,46,31,77,31,100,31,100,30,180,31,55,31,81,31,251,31,207,31,207,30,92,31,117,31,153,31,138,31,152,31,28,31,95,31,47,31,126,31,249,31,49,31,88,31,22,31,6,31,85,31,45,31,165,31,66,31,66,30,68,31,234,31,214,31,214,30,214,29,124,31,124,30,185,31,126,31,182,31,137,31,196,31,122,31,24,31,24,30,182,31,217,31,217,30,217,29,222,31,42,31,137,31,4,31,135,31,98,31,241,31,191,31,168,31,168,30,37,31,39,31,100,31,100,30,197,31,217,31,187,31,187,30,207,31,203,31,149,31,149,30,125,31,125,30,127,31,193,31,172,31,240,31,240,30,240,29,71,31,218,31,218,30,218,29,108,31,176,31,138,31,159,31,6,31,94,31,126,31,76,31,8,31,52,31,15,31,15,30,15,29,15,28,45,31,130,31,130,31,196,31,79,31,79,30,218,31,218,30,160,31,195,31,195,30,103,31,103,30,49,31,191,31,152,31,101,31,148,31,215,31,180,31,223,31,236,31,236,30,160,31,144,31,144,30,182,31,182,30,130,31,130,30,235,31,135,31,209,31,13,31,11,31,11,30,11,29,43,31,43,30,43,29,105,31,126,31,33,31,134,31,92,31,73,31,211,31,253,31,97,31,97,30,253,31,168,31,122,31,137,31,138,31,138,30,138,29,222,31,133,31,83,31,86,31,80,31,65,31,226,31,28,31,181,31,240,31,233,31,233,30,79,31,79,30,98,31,98,30,107,31,107,30,100,31,197,31,102,31,210,31,210,30,119,31,119,30,174,31,21,31,184,31,108,31,197,31,197,31,185,31,151,31,58,31,169,31,88,31,103,31,162,31,123,31,78,31,129,31,192,31,25,31,213,31,137,31,71,31,54,31,146,31,252,31,252,30,44,31,228,31,83,31,246,31,53,31,53,30,187,31,4,31,165,31,165,30,218,31,139,31,198,31,123,31,44,31,19,31,63,31,150,31,51,31,144,31,154,31,175,31,175,30,7,31,222,31,155,31,21,31,240,31,28,31,28,30,51,31,113,31,112,31,112,30,77,31,12,31,25,31,203,31,155,31,87,31,23,31,166,31,52,31,227,31,63,31,184,31,47,31,47,30,241,31,82,31,82,30,150,31,150,30,97,31,58,31,230,31,29,31,223,31,223,30,38,31,38,30,7,31,3,31,119,31,42,31,165,31,165,30,176,31,59,31,59,30,59,29,239,31,43,31,58,31,120,31,139,31,185,31,38,31,168,31,127,31,127,30,103,31,157,31,157,30,88,31,115,31,76,31,101,31,182,31,182,30,196,31,235,31,235,30,9,31,9,30,9,29,9,28,177,31,12,31,146,31,81,31,81,30,211,31,77,31,203,31,163,31,42,31,30,31,253,31,11,31,118,31,203,31,203,30,180,31,232,31,232,30,80,31,80,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
