-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_427 is
end project_tb_427;

architecture project_tb_arch_427 of project_tb_427 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 884;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,23,0,108,0,68,0,59,0,6,0,43,0,229,0,66,0,197,0,0,0,154,0,7,0,0,0,12,0,81,0,0,0,0,0,100,0,17,0,68,0,118,0,108,0,214,0,237,0,107,0,0,0,104,0,0,0,196,0,0,0,71,0,236,0,214,0,0,0,215,0,197,0,136,0,0,0,0,0,0,0,55,0,133,0,0,0,0,0,72,0,0,0,20,0,22,0,89,0,76,0,56,0,28,0,0,0,0,0,249,0,83,0,111,0,216,0,87,0,0,0,160,0,223,0,0,0,137,0,70,0,25,0,32,0,154,0,178,0,208,0,58,0,51,0,248,0,0,0,187,0,229,0,242,0,127,0,119,0,26,0,244,0,130,0,72,0,99,0,66,0,0,0,3,0,86,0,98,0,0,0,0,0,140,0,44,0,0,0,198,0,0,0,7,0,70,0,0,0,0,0,227,0,196,0,180,0,107,0,57,0,0,0,167,0,0,0,0,0,160,0,0,0,164,0,214,0,21,0,225,0,236,0,0,0,0,0,0,0,9,0,165,0,0,0,148,0,32,0,185,0,113,0,83,0,172,0,0,0,92,0,214,0,246,0,172,0,107,0,212,0,20,0,0,0,0,0,145,0,184,0,224,0,27,0,0,0,38,0,44,0,155,0,228,0,0,0,93,0,203,0,80,0,0,0,171,0,219,0,40,0,84,0,0,0,227,0,124,0,219,0,119,0,170,0,34,0,100,0,129,0,141,0,84,0,109,0,88,0,26,0,60,0,0,0,237,0,194,0,105,0,49,0,0,0,0,0,69,0,0,0,86,0,6,0,5,0,179,0,205,0,58,0,79,0,141,0,145,0,250,0,3,0,5,0,13,0,25,0,0,0,0,0,150,0,74,0,156,0,92,0,158,0,182,0,14,0,100,0,134,0,0,0,238,0,206,0,106,0,181,0,239,0,0,0,231,0,162,0,0,0,0,0,236,0,164,0,149,0,255,0,241,0,192,0,195,0,128,0,111,0,14,0,98,0,0,0,4,0,163,0,238,0,46,0,223,0,162,0,0,0,0,0,50,0,227,0,0,0,53,0,84,0,0,0,87,0,107,0,32,0,0,0,83,0,38,0,89,0,194,0,211,0,0,0,169,0,38,0,86,0,62,0,41,0,9,0,75,0,40,0,49,0,9,0,235,0,79,0,227,0,226,0,178,0,0,0,10,0,0,0,0,0,131,0,130,0,0,0,158,0,105,0,220,0,0,0,0,0,244,0,0,0,135,0,88,0,36,0,163,0,245,0,0,0,0,0,91,0,18,0,81,0,60,0,26,0,0,0,67,0,94,0,0,0,0,0,77,0,162,0,6,0,0,0,131,0,121,0,0,0,147,0,242,0,26,0,39,0,133,0,58,0,30,0,43,0,2,0,0,0,27,0,0,0,0,0,198,0,120,0,0,0,86,0,246,0,79,0,143,0,247,0,63,0,195,0,0,0,12,0,196,0,9,0,65,0,251,0,44,0,0,0,124,0,231,0,47,0,110,0,238,0,148,0,214,0,232,0,145,0,207,0,120,0,243,0,231,0,122,0,20,0,37,0,8,0,252,0,0,0,150,0,80,0,29,0,178,0,120,0,84,0,0,0,0,0,187,0,23,0,0,0,232,0,23,0,62,0,0,0,62,0,230,0,50,0,221,0,198,0,162,0,180,0,0,0,229,0,142,0,34,0,97,0,0,0,193,0,182,0,0,0,87,0,211,0,49,0,198,0,0,0,0,0,242,0,179,0,59,0,0,0,120,0,0,0,92,0,209,0,0,0,65,0,157,0,132,0,207,0,0,0,0,0,157,0,119,0,222,0,84,0,17,0,0,0,42,0,41,0,131,0,0,0,0,0,186,0,0,0,16,0,75,0,127,0,105,0,136,0,135,0,127,0,207,0,0,0,50,0,252,0,139,0,0,0,0,0,0,0,217,0,233,0,180,0,224,0,124,0,60,0,60,0,4,0,0,0,168,0,108,0,137,0,0,0,87,0,0,0,188,0,137,0,181,0,14,0,0,0,67,0,38,0,64,0,134,0,35,0,141,0,99,0,103,0,93,0,40,0,0,0,69,0,88,0,22,0,0,0,36,0,249,0,9,0,201,0,167,0,148,0,97,0,0,0,132,0,184,0,179,0,99,0,0,0,17,0,0,0,0,0,117,0,215,0,36,0,149,0,48,0,231,0,248,0,129,0,68,0,0,0,114,0,89,0,24,0,243,0,158,0,0,0,43,0,116,0,69,0,51,0,0,0,189,0,206,0,50,0,0,0,53,0,143,0,64,0,133,0,121,0,250,0,0,0,2,0,167,0,0,0,248,0,138,0,122,0,28,0,230,0,197,0,0,0,9,0,178,0,0,0,29,0,9,0,161,0,6,0,149,0,255,0,0,0,0,0,196,0,177,0,24,0,249,0,67,0,73,0,112,0,9,0,57,0,42,0,176,0,198,0,53,0,255,0,214,0,193,0,0,0,0,0,0,0,0,0,40,0,239,0,178,0,101,0,79,0,246,0,146,0,250,0,64,0,47,0,153,0,80,0,144,0,170,0,0,0,209,0,0,0,92,0,214,0,4,0,197,0,0,0,147,0,55,0,0,0,230,0,128,0,0,0,0,0,0,0,54,0,182,0,0,0,251,0,233,0,0,0,203,0,184,0,37,0,226,0,192,0,228,0,0,0,15,0,0,0,85,0,249,0,9,0,110,0,111,0,0,0,53,0,223,0,185,0,114,0,253,0,69,0,211,0,117,0,249,0,0,0,0,0,0,0,150,0,194,0,1,0,222,0,47,0,110,0,0,0,215,0,141,0,165,0,169,0,0,0,32,0,190,0,13,0,52,0,82,0,0,0,0,0,205,0,0,0,56,0,242,0,21,0,165,0,219,0,0,0,0,0,36,0,205,0,23,0,0,0,0,0,188,0,190,0,122,0,141,0,0,0,182,0,193,0,223,0,83,0,195,0,96,0,231,0,104,0,0,0,0,0,172,0,79,0,30,0,184,0,177,0,79,0,0,0,168,0,0,0,133,0,0,0,204,0,208,0,180,0,48,0,94,0,209,0,250,0,151,0,0,0,201,0,0,0,21,0,240,0,102,0,0,0,165,0,236,0,0,0,3,0,0,0,60,0,100,0,0,0,0,0,77,0,120,0,137,0,1,0,89,0,199,0,243,0,163,0,0,0,170,0,249,0,150,0,0,0,0,0,134,0,0,0,177,0,193,0,122,0,0,0,102,0,220,0,112,0,243,0,232,0,0,0,251,0,22,0,187,0,0,0,162,0,0,0,0,0,88,0,205,0,229,0,228,0,71,0,88,0,249,0,46,0,73,0,0,0,115,0,232,0,13,0,231,0,118,0,48,0,219,0,73,0,37,0,0,0,254,0,227,0,61,0,91,0,225,0,171,0,239,0,178,0,239,0,70,0,0,0,0,0,205,0,60,0,169,0,9,0,13,0,0,0,242,0,84,0,99,0,69,0,76,0,246,0,33,0,0,0,0,0,61,0,0,0,220,0,96,0,221,0,123,0,42,0,12,0,253,0,165,0,99,0,43,0,218,0,0,0,0,0,184,0,75,0,0,0,0,0,237,0,162,0,147,0,72,0,124,0,0,0,44,0,0,0,129,0,0,0,101,0,27,0,215,0,0,0,18,0,216,0,39,0,80,0,0,0,126,0,51,0,120,0,10,0,57,0,180,0,27,0,165,0,27,0,0,0,115,0,72,0,171,0,159,0,254,0,61,0,0,0,89,0,253,0,85,0,214,0,93,0,226,0,83,0,128,0,40,0,35,0,0,0,0,0,211,0,2,0,0,0,0,0,227,0,193,0,41,0,214,0,86,0,188,0,2,0,230,0,25,0,240,0,98,0,0,0,239,0,144,0,115,0,33,0,0,0,0,0,0,0,146,0,121,0,0,0,65,0,205,0,89,0,0,0,64,0);
signal scenario_full  : scenario_type := (0,0,23,31,108,31,68,31,59,31,6,31,43,31,229,31,66,31,197,31,197,30,154,31,7,31,7,30,12,31,81,31,81,30,81,29,100,31,17,31,68,31,118,31,108,31,214,31,237,31,107,31,107,30,104,31,104,30,196,31,196,30,71,31,236,31,214,31,214,30,215,31,197,31,136,31,136,30,136,29,136,28,55,31,133,31,133,30,133,29,72,31,72,30,20,31,22,31,89,31,76,31,56,31,28,31,28,30,28,29,249,31,83,31,111,31,216,31,87,31,87,30,160,31,223,31,223,30,137,31,70,31,25,31,32,31,154,31,178,31,208,31,58,31,51,31,248,31,248,30,187,31,229,31,242,31,127,31,119,31,26,31,244,31,130,31,72,31,99,31,66,31,66,30,3,31,86,31,98,31,98,30,98,29,140,31,44,31,44,30,198,31,198,30,7,31,70,31,70,30,70,29,227,31,196,31,180,31,107,31,57,31,57,30,167,31,167,30,167,29,160,31,160,30,164,31,214,31,21,31,225,31,236,31,236,30,236,29,236,28,9,31,165,31,165,30,148,31,32,31,185,31,113,31,83,31,172,31,172,30,92,31,214,31,246,31,172,31,107,31,212,31,20,31,20,30,20,29,145,31,184,31,224,31,27,31,27,30,38,31,44,31,155,31,228,31,228,30,93,31,203,31,80,31,80,30,171,31,219,31,40,31,84,31,84,30,227,31,124,31,219,31,119,31,170,31,34,31,100,31,129,31,141,31,84,31,109,31,88,31,26,31,60,31,60,30,237,31,194,31,105,31,49,31,49,30,49,29,69,31,69,30,86,31,6,31,5,31,179,31,205,31,58,31,79,31,141,31,145,31,250,31,3,31,5,31,13,31,25,31,25,30,25,29,150,31,74,31,156,31,92,31,158,31,182,31,14,31,100,31,134,31,134,30,238,31,206,31,106,31,181,31,239,31,239,30,231,31,162,31,162,30,162,29,236,31,164,31,149,31,255,31,241,31,192,31,195,31,128,31,111,31,14,31,98,31,98,30,4,31,163,31,238,31,46,31,223,31,162,31,162,30,162,29,50,31,227,31,227,30,53,31,84,31,84,30,87,31,107,31,32,31,32,30,83,31,38,31,89,31,194,31,211,31,211,30,169,31,38,31,86,31,62,31,41,31,9,31,75,31,40,31,49,31,9,31,235,31,79,31,227,31,226,31,178,31,178,30,10,31,10,30,10,29,131,31,130,31,130,30,158,31,105,31,220,31,220,30,220,29,244,31,244,30,135,31,88,31,36,31,163,31,245,31,245,30,245,29,91,31,18,31,81,31,60,31,26,31,26,30,67,31,94,31,94,30,94,29,77,31,162,31,6,31,6,30,131,31,121,31,121,30,147,31,242,31,26,31,39,31,133,31,58,31,30,31,43,31,2,31,2,30,27,31,27,30,27,29,198,31,120,31,120,30,86,31,246,31,79,31,143,31,247,31,63,31,195,31,195,30,12,31,196,31,9,31,65,31,251,31,44,31,44,30,124,31,231,31,47,31,110,31,238,31,148,31,214,31,232,31,145,31,207,31,120,31,243,31,231,31,122,31,20,31,37,31,8,31,252,31,252,30,150,31,80,31,29,31,178,31,120,31,84,31,84,30,84,29,187,31,23,31,23,30,232,31,23,31,62,31,62,30,62,31,230,31,50,31,221,31,198,31,162,31,180,31,180,30,229,31,142,31,34,31,97,31,97,30,193,31,182,31,182,30,87,31,211,31,49,31,198,31,198,30,198,29,242,31,179,31,59,31,59,30,120,31,120,30,92,31,209,31,209,30,65,31,157,31,132,31,207,31,207,30,207,29,157,31,119,31,222,31,84,31,17,31,17,30,42,31,41,31,131,31,131,30,131,29,186,31,186,30,16,31,75,31,127,31,105,31,136,31,135,31,127,31,207,31,207,30,50,31,252,31,139,31,139,30,139,29,139,28,217,31,233,31,180,31,224,31,124,31,60,31,60,31,4,31,4,30,168,31,108,31,137,31,137,30,87,31,87,30,188,31,137,31,181,31,14,31,14,30,67,31,38,31,64,31,134,31,35,31,141,31,99,31,103,31,93,31,40,31,40,30,69,31,88,31,22,31,22,30,36,31,249,31,9,31,201,31,167,31,148,31,97,31,97,30,132,31,184,31,179,31,99,31,99,30,17,31,17,30,17,29,117,31,215,31,36,31,149,31,48,31,231,31,248,31,129,31,68,31,68,30,114,31,89,31,24,31,243,31,158,31,158,30,43,31,116,31,69,31,51,31,51,30,189,31,206,31,50,31,50,30,53,31,143,31,64,31,133,31,121,31,250,31,250,30,2,31,167,31,167,30,248,31,138,31,122,31,28,31,230,31,197,31,197,30,9,31,178,31,178,30,29,31,9,31,161,31,6,31,149,31,255,31,255,30,255,29,196,31,177,31,24,31,249,31,67,31,73,31,112,31,9,31,57,31,42,31,176,31,198,31,53,31,255,31,214,31,193,31,193,30,193,29,193,28,193,27,40,31,239,31,178,31,101,31,79,31,246,31,146,31,250,31,64,31,47,31,153,31,80,31,144,31,170,31,170,30,209,31,209,30,92,31,214,31,4,31,197,31,197,30,147,31,55,31,55,30,230,31,128,31,128,30,128,29,128,28,54,31,182,31,182,30,251,31,233,31,233,30,203,31,184,31,37,31,226,31,192,31,228,31,228,30,15,31,15,30,85,31,249,31,9,31,110,31,111,31,111,30,53,31,223,31,185,31,114,31,253,31,69,31,211,31,117,31,249,31,249,30,249,29,249,28,150,31,194,31,1,31,222,31,47,31,110,31,110,30,215,31,141,31,165,31,169,31,169,30,32,31,190,31,13,31,52,31,82,31,82,30,82,29,205,31,205,30,56,31,242,31,21,31,165,31,219,31,219,30,219,29,36,31,205,31,23,31,23,30,23,29,188,31,190,31,122,31,141,31,141,30,182,31,193,31,223,31,83,31,195,31,96,31,231,31,104,31,104,30,104,29,172,31,79,31,30,31,184,31,177,31,79,31,79,30,168,31,168,30,133,31,133,30,204,31,208,31,180,31,48,31,94,31,209,31,250,31,151,31,151,30,201,31,201,30,21,31,240,31,102,31,102,30,165,31,236,31,236,30,3,31,3,30,60,31,100,31,100,30,100,29,77,31,120,31,137,31,1,31,89,31,199,31,243,31,163,31,163,30,170,31,249,31,150,31,150,30,150,29,134,31,134,30,177,31,193,31,122,31,122,30,102,31,220,31,112,31,243,31,232,31,232,30,251,31,22,31,187,31,187,30,162,31,162,30,162,29,88,31,205,31,229,31,228,31,71,31,88,31,249,31,46,31,73,31,73,30,115,31,232,31,13,31,231,31,118,31,48,31,219,31,73,31,37,31,37,30,254,31,227,31,61,31,91,31,225,31,171,31,239,31,178,31,239,31,70,31,70,30,70,29,205,31,60,31,169,31,9,31,13,31,13,30,242,31,84,31,99,31,69,31,76,31,246,31,33,31,33,30,33,29,61,31,61,30,220,31,96,31,221,31,123,31,42,31,12,31,253,31,165,31,99,31,43,31,218,31,218,30,218,29,184,31,75,31,75,30,75,29,237,31,162,31,147,31,72,31,124,31,124,30,44,31,44,30,129,31,129,30,101,31,27,31,215,31,215,30,18,31,216,31,39,31,80,31,80,30,126,31,51,31,120,31,10,31,57,31,180,31,27,31,165,31,27,31,27,30,115,31,72,31,171,31,159,31,254,31,61,31,61,30,89,31,253,31,85,31,214,31,93,31,226,31,83,31,128,31,40,31,35,31,35,30,35,29,211,31,2,31,2,30,2,29,227,31,193,31,41,31,214,31,86,31,188,31,2,31,230,31,25,31,240,31,98,31,98,30,239,31,144,31,115,31,33,31,33,30,33,29,33,28,146,31,121,31,121,30,65,31,205,31,89,31,89,30,64,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
