-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_78 is
end project_tb_78;

architecture project_tb_arch_78 of project_tb_78 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 770;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (159,0,0,0,22,0,151,0,161,0,229,0,254,0,96,0,51,0,94,0,120,0,179,0,70,0,13,0,0,0,1,0,54,0,0,0,64,0,0,0,170,0,41,0,216,0,39,0,249,0,7,0,212,0,67,0,252,0,197,0,0,0,121,0,0,0,201,0,177,0,33,0,207,0,142,0,0,0,216,0,97,0,183,0,115,0,120,0,90,0,20,0,249,0,0,0,28,0,92,0,55,0,238,0,0,0,239,0,33,0,97,0,0,0,253,0,220,0,99,0,117,0,216,0,54,0,191,0,98,0,0,0,155,0,61,0,217,0,246,0,44,0,83,0,223,0,242,0,11,0,168,0,0,0,50,0,141,0,143,0,76,0,0,0,75,0,0,0,14,0,19,0,93,0,211,0,162,0,147,0,213,0,69,0,160,0,0,0,86,0,239,0,41,0,0,0,175,0,73,0,0,0,238,0,29,0,8,0,248,0,73,0,0,0,57,0,200,0,214,0,84,0,162,0,5,0,246,0,136,0,151,0,171,0,229,0,116,0,135,0,211,0,49,0,177,0,221,0,100,0,70,0,107,0,105,0,0,0,116,0,13,0,0,0,94,0,109,0,183,0,43,0,35,0,159,0,22,0,0,0,0,0,10,0,37,0,56,0,0,0,0,0,85,0,82,0,42,0,245,0,137,0,61,0,145,0,4,0,145,0,133,0,97,0,123,0,88,0,0,0,109,0,77,0,101,0,159,0,134,0,151,0,74,0,119,0,152,0,199,0,141,0,0,0,14,0,245,0,231,0,0,0,151,0,232,0,0,0,57,0,73,0,67,0,142,0,207,0,53,0,59,0,21,0,225,0,17,0,245,0,107,0,0,0,0,0,12,0,42,0,0,0,112,0,118,0,0,0,85,0,157,0,115,0,87,0,76,0,0,0,102,0,82,0,136,0,70,0,136,0,75,0,1,0,220,0,0,0,95,0,143,0,240,0,191,0,134,0,6,0,167,0,133,0,202,0,241,0,94,0,119,0,3,0,196,0,181,0,0,0,19,0,224,0,157,0,222,0,113,0,84,0,73,0,210,0,216,0,0,0,0,0,255,0,57,0,197,0,176,0,144,0,20,0,12,0,66,0,37,0,187,0,170,0,143,0,0,0,236,0,225,0,140,0,179,0,210,0,0,0,164,0,0,0,222,0,0,0,242,0,236,0,0,0,0,0,155,0,28,0,205,0,169,0,213,0,101,0,0,0,119,0,182,0,238,0,0,0,117,0,0,0,153,0,78,0,135,0,0,0,64,0,0,0,250,0,165,0,76,0,241,0,227,0,187,0,150,0,196,0,0,0,0,0,0,0,160,0,0,0,135,0,72,0,0,0,0,0,171,0,223,0,8,0,119,0,11,0,123,0,221,0,57,0,214,0,11,0,117,0,131,0,51,0,0,0,228,0,94,0,203,0,171,0,4,0,19,0,0,0,0,0,113,0,58,0,0,0,218,0,60,0,215,0,221,0,35,0,217,0,75,0,157,0,223,0,242,0,116,0,207,0,111,0,5,0,12,0,0,0,137,0,24,0,56,0,0,0,203,0,27,0,231,0,170,0,1,0,65,0,67,0,130,0,0,0,40,0,0,0,0,0,172,0,237,0,148,0,0,0,168,0,188,0,15,0,0,0,0,0,194,0,0,0,0,0,242,0,19,0,38,0,127,0,211,0,244,0,151,0,0,0,129,0,216,0,0,0,232,0,117,0,96,0,254,0,0,0,74,0,163,0,0,0,216,0,0,0,208,0,111,0,0,0,216,0,188,0,0,0,121,0,170,0,42,0,0,0,249,0,225,0,27,0,11,0,183,0,118,0,172,0,0,0,179,0,129,0,0,0,0,0,197,0,0,0,0,0,57,0,18,0,212,0,206,0,198,0,15,0,28,0,175,0,162,0,27,0,201,0,17,0,179,0,0,0,184,0,0,0,0,0,48,0,55,0,175,0,51,0,144,0,147,0,250,0,240,0,253,0,106,0,243,0,34,0,42,0,100,0,112,0,244,0,241,0,64,0,50,0,0,0,21,0,42,0,125,0,237,0,0,0,155,0,0,0,41,0,52,0,0,0,234,0,91,0,0,0,202,0,152,0,10,0,53,0,198,0,144,0,81,0,210,0,108,0,5,0,32,0,196,0,89,0,172,0,254,0,1,0,0,0,63,0,77,0,8,0,101,0,0,0,147,0,68,0,0,0,0,0,146,0,121,0,12,0,0,0,217,0,233,0,176,0,132,0,145,0,0,0,0,0,146,0,10,0,160,0,250,0,0,0,230,0,0,0,125,0,167,0,221,0,18,0,230,0,100,0,18,0,157,0,128,0,36,0,0,0,28,0,208,0,0,0,8,0,176,0,41,0,0,0,184,0,0,0,128,0,150,0,36,0,78,0,250,0,108,0,45,0,118,0,25,0,126,0,125,0,0,0,2,0,105,0,212,0,104,0,82,0,78,0,0,0,5,0,226,0,53,0,142,0,0,0,11,0,87,0,4,0,136,0,218,0,228,0,95,0,0,0,211,0,70,0,0,0,116,0,37,0,160,0,156,0,131,0,122,0,36,0,248,0,183,0,241,0,0,0,94,0,158,0,5,0,0,0,0,0,0,0,10,0,116,0,122,0,89,0,0,0,138,0,159,0,60,0,240,0,82,0,0,0,21,0,238,0,26,0,31,0,29,0,140,0,220,0,70,0,74,0,78,0,0,0,227,0,84,0,153,0,114,0,22,0,121,0,89,0,250,0,103,0,94,0,176,0,0,0,250,0,204,0,182,0,103,0,83,0,0,0,0,0,41,0,0,0,231,0,204,0,125,0,58,0,46,0,169,0,72,0,0,0,0,0,37,0,119,0,122,0,187,0,9,0,124,0,88,0,0,0,86,0,195,0,245,0,69,0,105,0,116,0,30,0,188,0,195,0,97,0,0,0,168,0,0,0,0,0,215,0,101,0,155,0,0,0,0,0,31,0,223,0,90,0,0,0,111,0,120,0,109,0,141,0,207,0,18,0,76,0,84,0,173,0,20,0,0,0,36,0,56,0,36,0,72,0,165,0,233,0,89,0,0,0,220,0,128,0,11,0,38,0,181,0,113,0,171,0,0,0,0,0,112,0,18,0,148,0,134,0,194,0,0,0,15,0,222,0,72,0,0,0,136,0,210,0,145,0,229,0,254,0,162,0,0,0,163,0,217,0,255,0,247,0,187,0,0,0,10,0,182,0,49,0,110,0,0,0,222,0,0,0,189,0,114,0,0,0,3,0,80,0,114,0,85,0,73,0,4,0,78,0,114,0,21,0,94,0,75,0,107,0,0,0,61,0,216,0,124,0,12,0,255,0,89,0,0,0,140,0,204,0,39,0,121,0,30,0,0,0,227,0,96,0,30,0,45,0,0,0,166,0,50,0,0,0,4,0,93,0,0,0,110,0,192,0,146,0,178,0);
signal scenario_full  : scenario_type := (159,31,159,30,22,31,151,31,161,31,229,31,254,31,96,31,51,31,94,31,120,31,179,31,70,31,13,31,13,30,1,31,54,31,54,30,64,31,64,30,170,31,41,31,216,31,39,31,249,31,7,31,212,31,67,31,252,31,197,31,197,30,121,31,121,30,201,31,177,31,33,31,207,31,142,31,142,30,216,31,97,31,183,31,115,31,120,31,90,31,20,31,249,31,249,30,28,31,92,31,55,31,238,31,238,30,239,31,33,31,97,31,97,30,253,31,220,31,99,31,117,31,216,31,54,31,191,31,98,31,98,30,155,31,61,31,217,31,246,31,44,31,83,31,223,31,242,31,11,31,168,31,168,30,50,31,141,31,143,31,76,31,76,30,75,31,75,30,14,31,19,31,93,31,211,31,162,31,147,31,213,31,69,31,160,31,160,30,86,31,239,31,41,31,41,30,175,31,73,31,73,30,238,31,29,31,8,31,248,31,73,31,73,30,57,31,200,31,214,31,84,31,162,31,5,31,246,31,136,31,151,31,171,31,229,31,116,31,135,31,211,31,49,31,177,31,221,31,100,31,70,31,107,31,105,31,105,30,116,31,13,31,13,30,94,31,109,31,183,31,43,31,35,31,159,31,22,31,22,30,22,29,10,31,37,31,56,31,56,30,56,29,85,31,82,31,42,31,245,31,137,31,61,31,145,31,4,31,145,31,133,31,97,31,123,31,88,31,88,30,109,31,77,31,101,31,159,31,134,31,151,31,74,31,119,31,152,31,199,31,141,31,141,30,14,31,245,31,231,31,231,30,151,31,232,31,232,30,57,31,73,31,67,31,142,31,207,31,53,31,59,31,21,31,225,31,17,31,245,31,107,31,107,30,107,29,12,31,42,31,42,30,112,31,118,31,118,30,85,31,157,31,115,31,87,31,76,31,76,30,102,31,82,31,136,31,70,31,136,31,75,31,1,31,220,31,220,30,95,31,143,31,240,31,191,31,134,31,6,31,167,31,133,31,202,31,241,31,94,31,119,31,3,31,196,31,181,31,181,30,19,31,224,31,157,31,222,31,113,31,84,31,73,31,210,31,216,31,216,30,216,29,255,31,57,31,197,31,176,31,144,31,20,31,12,31,66,31,37,31,187,31,170,31,143,31,143,30,236,31,225,31,140,31,179,31,210,31,210,30,164,31,164,30,222,31,222,30,242,31,236,31,236,30,236,29,155,31,28,31,205,31,169,31,213,31,101,31,101,30,119,31,182,31,238,31,238,30,117,31,117,30,153,31,78,31,135,31,135,30,64,31,64,30,250,31,165,31,76,31,241,31,227,31,187,31,150,31,196,31,196,30,196,29,196,28,160,31,160,30,135,31,72,31,72,30,72,29,171,31,223,31,8,31,119,31,11,31,123,31,221,31,57,31,214,31,11,31,117,31,131,31,51,31,51,30,228,31,94,31,203,31,171,31,4,31,19,31,19,30,19,29,113,31,58,31,58,30,218,31,60,31,215,31,221,31,35,31,217,31,75,31,157,31,223,31,242,31,116,31,207,31,111,31,5,31,12,31,12,30,137,31,24,31,56,31,56,30,203,31,27,31,231,31,170,31,1,31,65,31,67,31,130,31,130,30,40,31,40,30,40,29,172,31,237,31,148,31,148,30,168,31,188,31,15,31,15,30,15,29,194,31,194,30,194,29,242,31,19,31,38,31,127,31,211,31,244,31,151,31,151,30,129,31,216,31,216,30,232,31,117,31,96,31,254,31,254,30,74,31,163,31,163,30,216,31,216,30,208,31,111,31,111,30,216,31,188,31,188,30,121,31,170,31,42,31,42,30,249,31,225,31,27,31,11,31,183,31,118,31,172,31,172,30,179,31,129,31,129,30,129,29,197,31,197,30,197,29,57,31,18,31,212,31,206,31,198,31,15,31,28,31,175,31,162,31,27,31,201,31,17,31,179,31,179,30,184,31,184,30,184,29,48,31,55,31,175,31,51,31,144,31,147,31,250,31,240,31,253,31,106,31,243,31,34,31,42,31,100,31,112,31,244,31,241,31,64,31,50,31,50,30,21,31,42,31,125,31,237,31,237,30,155,31,155,30,41,31,52,31,52,30,234,31,91,31,91,30,202,31,152,31,10,31,53,31,198,31,144,31,81,31,210,31,108,31,5,31,32,31,196,31,89,31,172,31,254,31,1,31,1,30,63,31,77,31,8,31,101,31,101,30,147,31,68,31,68,30,68,29,146,31,121,31,12,31,12,30,217,31,233,31,176,31,132,31,145,31,145,30,145,29,146,31,10,31,160,31,250,31,250,30,230,31,230,30,125,31,167,31,221,31,18,31,230,31,100,31,18,31,157,31,128,31,36,31,36,30,28,31,208,31,208,30,8,31,176,31,41,31,41,30,184,31,184,30,128,31,150,31,36,31,78,31,250,31,108,31,45,31,118,31,25,31,126,31,125,31,125,30,2,31,105,31,212,31,104,31,82,31,78,31,78,30,5,31,226,31,53,31,142,31,142,30,11,31,87,31,4,31,136,31,218,31,228,31,95,31,95,30,211,31,70,31,70,30,116,31,37,31,160,31,156,31,131,31,122,31,36,31,248,31,183,31,241,31,241,30,94,31,158,31,5,31,5,30,5,29,5,28,10,31,116,31,122,31,89,31,89,30,138,31,159,31,60,31,240,31,82,31,82,30,21,31,238,31,26,31,31,31,29,31,140,31,220,31,70,31,74,31,78,31,78,30,227,31,84,31,153,31,114,31,22,31,121,31,89,31,250,31,103,31,94,31,176,31,176,30,250,31,204,31,182,31,103,31,83,31,83,30,83,29,41,31,41,30,231,31,204,31,125,31,58,31,46,31,169,31,72,31,72,30,72,29,37,31,119,31,122,31,187,31,9,31,124,31,88,31,88,30,86,31,195,31,245,31,69,31,105,31,116,31,30,31,188,31,195,31,97,31,97,30,168,31,168,30,168,29,215,31,101,31,155,31,155,30,155,29,31,31,223,31,90,31,90,30,111,31,120,31,109,31,141,31,207,31,18,31,76,31,84,31,173,31,20,31,20,30,36,31,56,31,36,31,72,31,165,31,233,31,89,31,89,30,220,31,128,31,11,31,38,31,181,31,113,31,171,31,171,30,171,29,112,31,18,31,148,31,134,31,194,31,194,30,15,31,222,31,72,31,72,30,136,31,210,31,145,31,229,31,254,31,162,31,162,30,163,31,217,31,255,31,247,31,187,31,187,30,10,31,182,31,49,31,110,31,110,30,222,31,222,30,189,31,114,31,114,30,3,31,80,31,114,31,85,31,73,31,4,31,78,31,114,31,21,31,94,31,75,31,107,31,107,30,61,31,216,31,124,31,12,31,255,31,89,31,89,30,140,31,204,31,39,31,121,31,30,31,30,30,227,31,96,31,30,31,45,31,45,30,166,31,50,31,50,30,4,31,93,31,93,30,110,31,192,31,146,31,178,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
