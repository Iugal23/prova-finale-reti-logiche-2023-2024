-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 172;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (87,0,209,0,0,0,39,0,55,0,107,0,148,0,193,0,0,0,102,0,211,0,213,0,18,0,159,0,35,0,80,0,7,0,183,0,153,0,69,0,236,0,170,0,0,0,209,0,54,0,0,0,109,0,35,0,86,0,0,0,67,0,81,0,149,0,0,0,138,0,1,0,0,0,26,0,186,0,217,0,0,0,140,0,67,0,28,0,175,0,0,0,3,0,0,0,0,0,242,0,238,0,131,0,240,0,160,0,177,0,1,0,0,0,204,0,75,0,97,0,0,0,216,0,248,0,36,0,214,0,77,0,114,0,0,0,83,0,231,0,141,0,106,0,16,0,253,0,62,0,0,0,226,0,0,0,182,0,232,0,190,0,146,0,71,0,75,0,35,0,160,0,16,0,53,0,85,0,0,0,181,0,94,0,157,0,64,0,209,0,13,0,0,0,0,0,120,0,54,0,0,0,254,0,41,0,150,0,0,0,78,0,0,0,234,0,0,0,0,0,43,0,38,0,169,0,241,0,42,0,214,0,0,0,14,0,9,0,223,0,58,0,0,0,57,0,72,0,161,0,197,0,0,0,98,0,54,0,108,0,153,0,125,0,95,0,116,0,152,0,246,0,226,0,0,0,166,0,41,0,254,0,0,0,191,0,199,0,231,0,234,0,46,0,133,0,0,0,124,0,0,0,162,0,236,0,215,0,38,0,143,0,207,0,245,0,241,0,210,0,69,0,166,0,24,0,142,0,181,0,15,0,148,0,12,0,0,0,179,0,0,0,20,0);
signal scenario_full  : scenario_type := (87,31,209,31,209,30,39,31,55,31,107,31,148,31,193,31,193,30,102,31,211,31,213,31,18,31,159,31,35,31,80,31,7,31,183,31,153,31,69,31,236,31,170,31,170,30,209,31,54,31,54,30,109,31,35,31,86,31,86,30,67,31,81,31,149,31,149,30,138,31,1,31,1,30,26,31,186,31,217,31,217,30,140,31,67,31,28,31,175,31,175,30,3,31,3,30,3,29,242,31,238,31,131,31,240,31,160,31,177,31,1,31,1,30,204,31,75,31,97,31,97,30,216,31,248,31,36,31,214,31,77,31,114,31,114,30,83,31,231,31,141,31,106,31,16,31,253,31,62,31,62,30,226,31,226,30,182,31,232,31,190,31,146,31,71,31,75,31,35,31,160,31,16,31,53,31,85,31,85,30,181,31,94,31,157,31,64,31,209,31,13,31,13,30,13,29,120,31,54,31,54,30,254,31,41,31,150,31,150,30,78,31,78,30,234,31,234,30,234,29,43,31,38,31,169,31,241,31,42,31,214,31,214,30,14,31,9,31,223,31,58,31,58,30,57,31,72,31,161,31,197,31,197,30,98,31,54,31,108,31,153,31,125,31,95,31,116,31,152,31,246,31,226,31,226,30,166,31,41,31,254,31,254,30,191,31,199,31,231,31,234,31,46,31,133,31,133,30,124,31,124,30,162,31,236,31,215,31,38,31,143,31,207,31,245,31,241,31,210,31,69,31,166,31,24,31,142,31,181,31,15,31,148,31,12,31,12,30,179,31,179,30,20,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
