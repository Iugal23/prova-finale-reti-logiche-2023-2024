-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_155 is
end project_tb_155;

architecture project_tb_arch_155 of project_tb_155 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 674;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (233,0,248,0,83,0,0,0,105,0,0,0,23,0,156,0,255,0,9,0,95,0,99,0,43,0,221,0,120,0,135,0,26,0,56,0,144,0,148,0,75,0,98,0,191,0,129,0,242,0,214,0,73,0,0,0,174,0,233,0,25,0,217,0,0,0,0,0,235,0,134,0,28,0,136,0,80,0,132,0,182,0,121,0,56,0,194,0,238,0,0,0,0,0,226,0,148,0,47,0,251,0,190,0,193,0,198,0,99,0,220,0,163,0,0,0,58,0,0,0,73,0,0,0,60,0,0,0,241,0,95,0,237,0,12,0,0,0,233,0,25,0,73,0,64,0,108,0,52,0,17,0,172,0,221,0,0,0,0,0,181,0,10,0,7,0,0,0,57,0,0,0,21,0,146,0,13,0,214,0,0,0,130,0,0,0,166,0,0,0,186,0,161,0,101,0,153,0,200,0,0,0,171,0,95,0,145,0,97,0,233,0,54,0,123,0,0,0,0,0,11,0,219,0,107,0,99,0,163,0,0,0,230,0,64,0,245,0,0,0,101,0,0,0,201,0,78,0,90,0,0,0,43,0,32,0,0,0,100,0,232,0,228,0,124,0,227,0,148,0,0,0,226,0,0,0,243,0,223,0,47,0,228,0,29,0,127,0,0,0,5,0,71,0,0,0,212,0,128,0,49,0,208,0,109,0,113,0,0,0,40,0,183,0,215,0,136,0,121,0,216,0,173,0,9,0,140,0,150,0,135,0,207,0,0,0,59,0,59,0,0,0,249,0,78,0,198,0,23,0,0,0,233,0,0,0,151,0,169,0,196,0,14,0,27,0,0,0,2,0,47,0,10,0,129,0,236,0,49,0,93,0,238,0,177,0,0,0,40,0,0,0,22,0,92,0,82,0,0,0,158,0,185,0,0,0,0,0,0,0,206,0,150,0,33,0,171,0,214,0,124,0,0,0,0,0,128,0,183,0,0,0,219,0,200,0,74,0,0,0,35,0,51,0,201,0,0,0,91,0,0,0,159,0,119,0,75,0,37,0,232,0,28,0,182,0,179,0,153,0,239,0,201,0,0,0,0,0,23,0,95,0,0,0,233,0,1,0,0,0,253,0,31,0,131,0,0,0,168,0,204,0,135,0,90,0,68,0,0,0,84,0,236,0,0,0,95,0,100,0,168,0,0,0,53,0,53,0,0,0,59,0,202,0,0,0,48,0,199,0,170,0,215,0,0,0,40,0,15,0,83,0,149,0,159,0,75,0,166,0,184,0,251,0,175,0,90,0,214,0,136,0,220,0,0,0,117,0,16,0,151,0,91,0,180,0,232,0,248,0,26,0,73,0,223,0,242,0,5,0,233,0,0,0,32,0,247,0,118,0,54,0,0,0,0,0,29,0,0,0,171,0,0,0,174,0,153,0,177,0,0,0,220,0,65,0,74,0,95,0,63,0,84,0,193,0,97,0,154,0,175,0,49,0,96,0,250,0,126,0,132,0,16,0,54,0,208,0,217,0,228,0,230,0,0,0,244,0,229,0,0,0,203,0,28,0,111,0,0,0,26,0,136,0,0,0,154,0,0,0,143,0,128,0,0,0,240,0,71,0,0,0,206,0,27,0,0,0,0,0,211,0,183,0,160,0,90,0,254,0,162,0,52,0,131,0,206,0,163,0,0,0,0,0,0,0,235,0,155,0,237,0,211,0,197,0,124,0,0,0,0,0,154,0,64,0,24,0,12,0,0,0,235,0,103,0,0,0,160,0,206,0,200,0,251,0,152,0,79,0,96,0,165,0,46,0,5,0,171,0,131,0,90,0,1,0,255,0,141,0,114,0,252,0,0,0,0,0,20,0,11,0,141,0,0,0,194,0,69,0,48,0,234,0,197,0,218,0,54,0,0,0,114,0,48,0,0,0,26,0,159,0,0,0,252,0,175,0,169,0,100,0,0,0,0,0,0,0,128,0,243,0,0,0,223,0,195,0,40,0,92,0,138,0,234,0,0,0,183,0,97,0,87,0,0,0,127,0,80,0,109,0,0,0,0,0,94,0,221,0,138,0,219,0,15,0,33,0,190,0,195,0,0,0,219,0,234,0,22,0,20,0,231,0,146,0,114,0,181,0,3,0,132,0,8,0,75,0,132,0,154,0,246,0,143,0,0,0,115,0,146,0,188,0,120,0,193,0,203,0,85,0,49,0,43,0,83,0,109,0,197,0,28,0,132,0,168,0,224,0,203,0,0,0,91,0,45,0,198,0,45,0,242,0,0,0,184,0,0,0,91,0,0,0,0,0,200,0,58,0,43,0,0,0,0,0,11,0,205,0,128,0,18,0,33,0,191,0,52,0,88,0,68,0,67,0,116,0,226,0,243,0,206,0,144,0,0,0,86,0,204,0,115,0,0,0,72,0,78,0,0,0,77,0,191,0,227,0,129,0,132,0,48,0,182,0,194,0,19,0,25,0,37,0,123,0,208,0,225,0,250,0,0,0,185,0,97,0,214,0,88,0,73,0,0,0,0,0,39,0,181,0,131,0,192,0,0,0,46,0,0,0,198,0,88,0,125,0,8,0,0,0,0,0,228,0,76,0,213,0,0,0,157,0,85,0,67,0,97,0,89,0,58,0,243,0,182,0,69,0,167,0,199,0,58,0,155,0,96,0,191,0,22,0,179,0,67,0,108,0,188,0,101,0,34,0,169,0,230,0,0,0,40,0,0,0,133,0,43,0,9,0,237,0,0,0,19,0,69,0,119,0,194,0,0,0,164,0,112,0,206,0,56,0,233,0,246,0,145,0,84,0,255,0,212,0,111,0,176,0,177,0,59,0,46,0,0,0,45,0,202,0,56,0,70,0,197,0,172,0,103,0,165,0,231,0,16,0,246,0,94,0,165,0,116,0,95,0,46,0,248,0,203,0,58,0,77,0,6,0,108,0,244,0,96,0,55,0,104,0,0,0,147,0,157,0,99,0,171,0,141,0,17,0,58,0,76,0,229,0,50,0,187,0,252,0,248,0,0,0,217,0,142,0,204,0,0,0);
signal scenario_full  : scenario_type := (233,31,248,31,83,31,83,30,105,31,105,30,23,31,156,31,255,31,9,31,95,31,99,31,43,31,221,31,120,31,135,31,26,31,56,31,144,31,148,31,75,31,98,31,191,31,129,31,242,31,214,31,73,31,73,30,174,31,233,31,25,31,217,31,217,30,217,29,235,31,134,31,28,31,136,31,80,31,132,31,182,31,121,31,56,31,194,31,238,31,238,30,238,29,226,31,148,31,47,31,251,31,190,31,193,31,198,31,99,31,220,31,163,31,163,30,58,31,58,30,73,31,73,30,60,31,60,30,241,31,95,31,237,31,12,31,12,30,233,31,25,31,73,31,64,31,108,31,52,31,17,31,172,31,221,31,221,30,221,29,181,31,10,31,7,31,7,30,57,31,57,30,21,31,146,31,13,31,214,31,214,30,130,31,130,30,166,31,166,30,186,31,161,31,101,31,153,31,200,31,200,30,171,31,95,31,145,31,97,31,233,31,54,31,123,31,123,30,123,29,11,31,219,31,107,31,99,31,163,31,163,30,230,31,64,31,245,31,245,30,101,31,101,30,201,31,78,31,90,31,90,30,43,31,32,31,32,30,100,31,232,31,228,31,124,31,227,31,148,31,148,30,226,31,226,30,243,31,223,31,47,31,228,31,29,31,127,31,127,30,5,31,71,31,71,30,212,31,128,31,49,31,208,31,109,31,113,31,113,30,40,31,183,31,215,31,136,31,121,31,216,31,173,31,9,31,140,31,150,31,135,31,207,31,207,30,59,31,59,31,59,30,249,31,78,31,198,31,23,31,23,30,233,31,233,30,151,31,169,31,196,31,14,31,27,31,27,30,2,31,47,31,10,31,129,31,236,31,49,31,93,31,238,31,177,31,177,30,40,31,40,30,22,31,92,31,82,31,82,30,158,31,185,31,185,30,185,29,185,28,206,31,150,31,33,31,171,31,214,31,124,31,124,30,124,29,128,31,183,31,183,30,219,31,200,31,74,31,74,30,35,31,51,31,201,31,201,30,91,31,91,30,159,31,119,31,75,31,37,31,232,31,28,31,182,31,179,31,153,31,239,31,201,31,201,30,201,29,23,31,95,31,95,30,233,31,1,31,1,30,253,31,31,31,131,31,131,30,168,31,204,31,135,31,90,31,68,31,68,30,84,31,236,31,236,30,95,31,100,31,168,31,168,30,53,31,53,31,53,30,59,31,202,31,202,30,48,31,199,31,170,31,215,31,215,30,40,31,15,31,83,31,149,31,159,31,75,31,166,31,184,31,251,31,175,31,90,31,214,31,136,31,220,31,220,30,117,31,16,31,151,31,91,31,180,31,232,31,248,31,26,31,73,31,223,31,242,31,5,31,233,31,233,30,32,31,247,31,118,31,54,31,54,30,54,29,29,31,29,30,171,31,171,30,174,31,153,31,177,31,177,30,220,31,65,31,74,31,95,31,63,31,84,31,193,31,97,31,154,31,175,31,49,31,96,31,250,31,126,31,132,31,16,31,54,31,208,31,217,31,228,31,230,31,230,30,244,31,229,31,229,30,203,31,28,31,111,31,111,30,26,31,136,31,136,30,154,31,154,30,143,31,128,31,128,30,240,31,71,31,71,30,206,31,27,31,27,30,27,29,211,31,183,31,160,31,90,31,254,31,162,31,52,31,131,31,206,31,163,31,163,30,163,29,163,28,235,31,155,31,237,31,211,31,197,31,124,31,124,30,124,29,154,31,64,31,24,31,12,31,12,30,235,31,103,31,103,30,160,31,206,31,200,31,251,31,152,31,79,31,96,31,165,31,46,31,5,31,171,31,131,31,90,31,1,31,255,31,141,31,114,31,252,31,252,30,252,29,20,31,11,31,141,31,141,30,194,31,69,31,48,31,234,31,197,31,218,31,54,31,54,30,114,31,48,31,48,30,26,31,159,31,159,30,252,31,175,31,169,31,100,31,100,30,100,29,100,28,128,31,243,31,243,30,223,31,195,31,40,31,92,31,138,31,234,31,234,30,183,31,97,31,87,31,87,30,127,31,80,31,109,31,109,30,109,29,94,31,221,31,138,31,219,31,15,31,33,31,190,31,195,31,195,30,219,31,234,31,22,31,20,31,231,31,146,31,114,31,181,31,3,31,132,31,8,31,75,31,132,31,154,31,246,31,143,31,143,30,115,31,146,31,188,31,120,31,193,31,203,31,85,31,49,31,43,31,83,31,109,31,197,31,28,31,132,31,168,31,224,31,203,31,203,30,91,31,45,31,198,31,45,31,242,31,242,30,184,31,184,30,91,31,91,30,91,29,200,31,58,31,43,31,43,30,43,29,11,31,205,31,128,31,18,31,33,31,191,31,52,31,88,31,68,31,67,31,116,31,226,31,243,31,206,31,144,31,144,30,86,31,204,31,115,31,115,30,72,31,78,31,78,30,77,31,191,31,227,31,129,31,132,31,48,31,182,31,194,31,19,31,25,31,37,31,123,31,208,31,225,31,250,31,250,30,185,31,97,31,214,31,88,31,73,31,73,30,73,29,39,31,181,31,131,31,192,31,192,30,46,31,46,30,198,31,88,31,125,31,8,31,8,30,8,29,228,31,76,31,213,31,213,30,157,31,85,31,67,31,97,31,89,31,58,31,243,31,182,31,69,31,167,31,199,31,58,31,155,31,96,31,191,31,22,31,179,31,67,31,108,31,188,31,101,31,34,31,169,31,230,31,230,30,40,31,40,30,133,31,43,31,9,31,237,31,237,30,19,31,69,31,119,31,194,31,194,30,164,31,112,31,206,31,56,31,233,31,246,31,145,31,84,31,255,31,212,31,111,31,176,31,177,31,59,31,46,31,46,30,45,31,202,31,56,31,70,31,197,31,172,31,103,31,165,31,231,31,16,31,246,31,94,31,165,31,116,31,95,31,46,31,248,31,203,31,58,31,77,31,6,31,108,31,244,31,96,31,55,31,104,31,104,30,147,31,157,31,99,31,171,31,141,31,17,31,58,31,76,31,229,31,50,31,187,31,252,31,248,31,248,30,217,31,142,31,204,31,204,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
