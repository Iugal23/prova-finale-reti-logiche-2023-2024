-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_913 is
end project_tb_913;

architecture project_tb_arch_913 of project_tb_913 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 749;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (30,0,95,0,34,0,0,0,0,0,44,0,42,0,0,0,0,0,147,0,81,0,0,0,142,0,51,0,54,0,174,0,29,0,0,0,193,0,0,0,0,0,98,0,0,0,31,0,0,0,1,0,102,0,105,0,16,0,105,0,0,0,18,0,182,0,176,0,123,0,50,0,160,0,65,0,156,0,62,0,130,0,186,0,0,0,125,0,107,0,238,0,91,0,103,0,234,0,219,0,0,0,59,0,241,0,154,0,221,0,0,0,174,0,196,0,50,0,47,0,5,0,214,0,44,0,143,0,180,0,42,0,112,0,0,0,219,0,153,0,194,0,125,0,46,0,0,0,71,0,128,0,0,0,193,0,127,0,187,0,0,0,238,0,0,0,114,0,180,0,108,0,241,0,110,0,0,0,225,0,37,0,207,0,230,0,126,0,15,0,46,0,62,0,138,0,0,0,7,0,130,0,0,0,98,0,121,0,44,0,91,0,118,0,0,0,129,0,227,0,0,0,0,0,20,0,248,0,0,0,191,0,0,0,0,0,0,0,0,0,169,0,225,0,0,0,206,0,0,0,172,0,0,0,115,0,138,0,106,0,197,0,0,0,128,0,207,0,38,0,0,0,0,0,200,0,77,0,76,0,90,0,29,0,215,0,0,0,15,0,15,0,128,0,62,0,33,0,238,0,12,0,221,0,254,0,215,0,138,0,255,0,206,0,85,0,40,0,245,0,132,0,0,0,58,0,0,0,52,0,0,0,125,0,211,0,50,0,173,0,31,0,0,0,133,0,217,0,94,0,122,0,221,0,233,0,24,0,121,0,220,0,0,0,127,0,208,0,51,0,159,0,221,0,0,0,174,0,108,0,46,0,155,0,139,0,48,0,244,0,109,0,212,0,132,0,253,0,178,0,39,0,233,0,37,0,41,0,0,0,166,0,245,0,181,0,165,0,101,0,0,0,254,0,139,0,174,0,14,0,93,0,188,0,223,0,52,0,0,0,0,0,40,0,9,0,95,0,166,0,219,0,171,0,104,0,29,0,160,0,185,0,176,0,0,0,15,0,0,0,140,0,0,0,199,0,10,0,254,0,0,0,103,0,209,0,180,0,224,0,0,0,0,0,236,0,149,0,191,0,201,0,0,0,223,0,29,0,197,0,22,0,205,0,168,0,83,0,0,0,100,0,50,0,179,0,12,0,121,0,0,0,0,0,196,0,4,0,0,0,71,0,142,0,0,0,60,0,220,0,27,0,0,0,90,0,0,0,163,0,135,0,1,0,186,0,234,0,111,0,0,0,36,0,135,0,183,0,206,0,185,0,179,0,212,0,226,0,0,0,7,0,48,0,100,0,215,0,75,0,102,0,0,0,172,0,59,0,204,0,0,0,99,0,127,0,110,0,4,0,131,0,54,0,160,0,160,0,216,0,55,0,0,0,150,0,98,0,8,0,254,0,0,0,114,0,33,0,0,0,64,0,217,0,231,0,130,0,138,0,171,0,252,0,27,0,0,0,122,0,0,0,200,0,22,0,134,0,0,0,166,0,6,0,65,0,156,0,178,0,104,0,113,0,0,0,0,0,206,0,145,0,92,0,0,0,0,0,0,0,214,0,137,0,54,0,39,0,161,0,65,0,118,0,0,0,226,0,39,0,0,0,162,0,145,0,169,0,166,0,0,0,0,0,116,0,95,0,32,0,230,0,0,0,243,0,75,0,83,0,216,0,119,0,207,0,192,0,197,0,54,0,30,0,167,0,249,0,3,0,0,0,0,0,42,0,247,0,103,0,176,0,0,0,154,0,0,0,0,0,75,0,89,0,0,0,0,0,0,0,172,0,53,0,44,0,210,0,0,0,129,0,0,0,45,0,77,0,32,0,205,0,233,0,104,0,180,0,89,0,4,0,228,0,231,0,0,0,230,0,220,0,193,0,0,0,254,0,45,0,17,0,160,0,22,0,29,0,139,0,84,0,59,0,44,0,0,0,175,0,106,0,91,0,42,0,0,0,59,0,178,0,101,0,177,0,113,0,213,0,246,0,120,0,0,0,110,0,29,0,50,0,163,0,187,0,195,0,67,0,107,0,1,0,46,0,115,0,175,0,232,0,218,0,176,0,0,0,91,0,0,0,219,0,0,0,13,0,127,0,129,0,14,0,0,0,7,0,99,0,97,0,89,0,195,0,134,0,0,0,107,0,66,0,0,0,69,0,0,0,228,0,232,0,54,0,212,0,99,0,1,0,116,0,180,0,186,0,145,0,0,0,243,0,175,0,165,0,75,0,175,0,0,0,24,0,224,0,96,0,203,0,43,0,245,0,0,0,84,0,240,0,28,0,0,0,11,0,0,0,119,0,191,0,0,0,31,0,170,0,151,0,104,0,49,0,2,0,0,0,144,0,80,0,68,0,129,0,92,0,77,0,90,0,172,0,253,0,174,0,85,0,0,0,189,0,0,0,190,0,145,0,180,0,47,0,34,0,6,0,157,0,0,0,224,0,10,0,120,0,73,0,0,0,0,0,147,0,0,0,0,0,202,0,68,0,242,0,38,0,0,0,0,0,0,0,141,0,116,0,186,0,238,0,83,0,0,0,104,0,0,0,82,0,233,0,198,0,145,0,39,0,42,0,88,0,0,0,147,0,0,0,75,0,171,0,105,0,201,0,105,0,0,0,52,0,77,0,181,0,85,0,167,0,70,0,214,0,254,0,0,0,16,0,253,0,123,0,166,0,155,0,2,0,5,0,0,0,0,0,59,0,233,0,76,0,183,0,0,0,131,0,209,0,150,0,254,0,91,0,0,0,245,0,49,0,99,0,14,0,207,0,147,0,152,0,28,0,211,0,213,0,0,0,34,0,12,0,205,0,18,0,0,0,0,0,0,0,167,0,189,0,170,0,232,0,156,0,99,0,127,0,214,0,202,0,0,0,219,0,160,0,0,0,60,0,108,0,0,0,114,0,245,0,227,0,150,0,89,0,242,0,144,0,0,0,0,0,83,0,0,0,190,0,82,0,223,0,0,0,199,0,104,0,0,0,98,0,0,0,90,0,198,0,73,0,0,0,0,0,0,0,221,0,207,0,49,0,209,0,0,0,70,0,228,0,67,0,57,0,200,0,91,0,155,0,227,0,87,0,191,0,76,0,0,0,94,0,64,0,37,0,70,0,43,0,0,0,239,0,0,0,50,0,115,0,242,0,111,0,129,0,36,0,146,0,47,0,37,0,233,0,0,0,0,0,0,0,173,0,242,0,0,0,193,0,136,0,0,0,115,0,83,0,0,0,108,0,186,0,147,0,81,0,219,0,154,0,0,0,0,0,0,0,76,0,49,0,236,0,0,0,0,0,0,0,237,0,197,0,156,0,0,0,39,0,214,0);
signal scenario_full  : scenario_type := (30,31,95,31,34,31,34,30,34,29,44,31,42,31,42,30,42,29,147,31,81,31,81,30,142,31,51,31,54,31,174,31,29,31,29,30,193,31,193,30,193,29,98,31,98,30,31,31,31,30,1,31,102,31,105,31,16,31,105,31,105,30,18,31,182,31,176,31,123,31,50,31,160,31,65,31,156,31,62,31,130,31,186,31,186,30,125,31,107,31,238,31,91,31,103,31,234,31,219,31,219,30,59,31,241,31,154,31,221,31,221,30,174,31,196,31,50,31,47,31,5,31,214,31,44,31,143,31,180,31,42,31,112,31,112,30,219,31,153,31,194,31,125,31,46,31,46,30,71,31,128,31,128,30,193,31,127,31,187,31,187,30,238,31,238,30,114,31,180,31,108,31,241,31,110,31,110,30,225,31,37,31,207,31,230,31,126,31,15,31,46,31,62,31,138,31,138,30,7,31,130,31,130,30,98,31,121,31,44,31,91,31,118,31,118,30,129,31,227,31,227,30,227,29,20,31,248,31,248,30,191,31,191,30,191,29,191,28,191,27,169,31,225,31,225,30,206,31,206,30,172,31,172,30,115,31,138,31,106,31,197,31,197,30,128,31,207,31,38,31,38,30,38,29,200,31,77,31,76,31,90,31,29,31,215,31,215,30,15,31,15,31,128,31,62,31,33,31,238,31,12,31,221,31,254,31,215,31,138,31,255,31,206,31,85,31,40,31,245,31,132,31,132,30,58,31,58,30,52,31,52,30,125,31,211,31,50,31,173,31,31,31,31,30,133,31,217,31,94,31,122,31,221,31,233,31,24,31,121,31,220,31,220,30,127,31,208,31,51,31,159,31,221,31,221,30,174,31,108,31,46,31,155,31,139,31,48,31,244,31,109,31,212,31,132,31,253,31,178,31,39,31,233,31,37,31,41,31,41,30,166,31,245,31,181,31,165,31,101,31,101,30,254,31,139,31,174,31,14,31,93,31,188,31,223,31,52,31,52,30,52,29,40,31,9,31,95,31,166,31,219,31,171,31,104,31,29,31,160,31,185,31,176,31,176,30,15,31,15,30,140,31,140,30,199,31,10,31,254,31,254,30,103,31,209,31,180,31,224,31,224,30,224,29,236,31,149,31,191,31,201,31,201,30,223,31,29,31,197,31,22,31,205,31,168,31,83,31,83,30,100,31,50,31,179,31,12,31,121,31,121,30,121,29,196,31,4,31,4,30,71,31,142,31,142,30,60,31,220,31,27,31,27,30,90,31,90,30,163,31,135,31,1,31,186,31,234,31,111,31,111,30,36,31,135,31,183,31,206,31,185,31,179,31,212,31,226,31,226,30,7,31,48,31,100,31,215,31,75,31,102,31,102,30,172,31,59,31,204,31,204,30,99,31,127,31,110,31,4,31,131,31,54,31,160,31,160,31,216,31,55,31,55,30,150,31,98,31,8,31,254,31,254,30,114,31,33,31,33,30,64,31,217,31,231,31,130,31,138,31,171,31,252,31,27,31,27,30,122,31,122,30,200,31,22,31,134,31,134,30,166,31,6,31,65,31,156,31,178,31,104,31,113,31,113,30,113,29,206,31,145,31,92,31,92,30,92,29,92,28,214,31,137,31,54,31,39,31,161,31,65,31,118,31,118,30,226,31,39,31,39,30,162,31,145,31,169,31,166,31,166,30,166,29,116,31,95,31,32,31,230,31,230,30,243,31,75,31,83,31,216,31,119,31,207,31,192,31,197,31,54,31,30,31,167,31,249,31,3,31,3,30,3,29,42,31,247,31,103,31,176,31,176,30,154,31,154,30,154,29,75,31,89,31,89,30,89,29,89,28,172,31,53,31,44,31,210,31,210,30,129,31,129,30,45,31,77,31,32,31,205,31,233,31,104,31,180,31,89,31,4,31,228,31,231,31,231,30,230,31,220,31,193,31,193,30,254,31,45,31,17,31,160,31,22,31,29,31,139,31,84,31,59,31,44,31,44,30,175,31,106,31,91,31,42,31,42,30,59,31,178,31,101,31,177,31,113,31,213,31,246,31,120,31,120,30,110,31,29,31,50,31,163,31,187,31,195,31,67,31,107,31,1,31,46,31,115,31,175,31,232,31,218,31,176,31,176,30,91,31,91,30,219,31,219,30,13,31,127,31,129,31,14,31,14,30,7,31,99,31,97,31,89,31,195,31,134,31,134,30,107,31,66,31,66,30,69,31,69,30,228,31,232,31,54,31,212,31,99,31,1,31,116,31,180,31,186,31,145,31,145,30,243,31,175,31,165,31,75,31,175,31,175,30,24,31,224,31,96,31,203,31,43,31,245,31,245,30,84,31,240,31,28,31,28,30,11,31,11,30,119,31,191,31,191,30,31,31,170,31,151,31,104,31,49,31,2,31,2,30,144,31,80,31,68,31,129,31,92,31,77,31,90,31,172,31,253,31,174,31,85,31,85,30,189,31,189,30,190,31,145,31,180,31,47,31,34,31,6,31,157,31,157,30,224,31,10,31,120,31,73,31,73,30,73,29,147,31,147,30,147,29,202,31,68,31,242,31,38,31,38,30,38,29,38,28,141,31,116,31,186,31,238,31,83,31,83,30,104,31,104,30,82,31,233,31,198,31,145,31,39,31,42,31,88,31,88,30,147,31,147,30,75,31,171,31,105,31,201,31,105,31,105,30,52,31,77,31,181,31,85,31,167,31,70,31,214,31,254,31,254,30,16,31,253,31,123,31,166,31,155,31,2,31,5,31,5,30,5,29,59,31,233,31,76,31,183,31,183,30,131,31,209,31,150,31,254,31,91,31,91,30,245,31,49,31,99,31,14,31,207,31,147,31,152,31,28,31,211,31,213,31,213,30,34,31,12,31,205,31,18,31,18,30,18,29,18,28,167,31,189,31,170,31,232,31,156,31,99,31,127,31,214,31,202,31,202,30,219,31,160,31,160,30,60,31,108,31,108,30,114,31,245,31,227,31,150,31,89,31,242,31,144,31,144,30,144,29,83,31,83,30,190,31,82,31,223,31,223,30,199,31,104,31,104,30,98,31,98,30,90,31,198,31,73,31,73,30,73,29,73,28,221,31,207,31,49,31,209,31,209,30,70,31,228,31,67,31,57,31,200,31,91,31,155,31,227,31,87,31,191,31,76,31,76,30,94,31,64,31,37,31,70,31,43,31,43,30,239,31,239,30,50,31,115,31,242,31,111,31,129,31,36,31,146,31,47,31,37,31,233,31,233,30,233,29,233,28,173,31,242,31,242,30,193,31,136,31,136,30,115,31,83,31,83,30,108,31,186,31,147,31,81,31,219,31,154,31,154,30,154,29,154,28,76,31,49,31,236,31,236,30,236,29,236,28,237,31,197,31,156,31,156,30,39,31,214,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
