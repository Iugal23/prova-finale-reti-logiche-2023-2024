-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_13 is
end project_tb_13;

architecture project_tb_arch_13 of project_tb_13 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 217;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (45,0,213,0,210,0,250,0,184,0,1,0,21,0,214,0,199,0,95,0,88,0,58,0,211,0,0,0,20,0,14,0,75,0,222,0,0,0,162,0,65,0,176,0,88,0,0,0,46,0,145,0,162,0,164,0,54,0,79,0,54,0,25,0,0,0,142,0,43,0,25,0,5,0,190,0,24,0,0,0,0,0,100,0,122,0,101,0,202,0,74,0,0,0,156,0,73,0,48,0,101,0,103,0,169,0,99,0,74,0,80,0,0,0,0,0,41,0,213,0,56,0,34,0,89,0,115,0,219,0,112,0,80,0,229,0,24,0,0,0,2,0,154,0,0,0,0,0,143,0,141,0,148,0,0,0,193,0,65,0,0,0,202,0,0,0,61,0,188,0,162,0,184,0,124,0,0,0,0,0,0,0,211,0,97,0,229,0,117,0,90,0,130,0,9,0,0,0,158,0,46,0,18,0,151,0,199,0,24,0,182,0,52,0,199,0,20,0,0,0,16,0,0,0,24,0,86,0,103,0,140,0,0,0,204,0,0,0,0,0,255,0,163,0,205,0,158,0,0,0,195,0,3,0,225,0,0,0,240,0,134,0,218,0,0,0,100,0,195,0,100,0,199,0,158,0,206,0,191,0,163,0,151,0,190,0,31,0,180,0,180,0,222,0,27,0,58,0,170,0,96,0,80,0,226,0,212,0,174,0,0,0,0,0,111,0,116,0,170,0,1,0,136,0,20,0,0,0,24,0,73,0,79,0,31,0,0,0,100,0,0,0,135,0,159,0,19,0,38,0,129,0,86,0,198,0,184,0,86,0,168,0,7,0,124,0,247,0,191,0,23,0,0,0,101,0,0,0,0,0,244,0,145,0,23,0,38,0,3,0,234,0,0,0,104,0,0,0,69,0,155,0,220,0,192,0,233,0,102,0,128,0,29,0,105,0,36,0,0,0,0,0,160,0,0,0,0,0,160,0,173,0,20,0);
signal scenario_full  : scenario_type := (45,31,213,31,210,31,250,31,184,31,1,31,21,31,214,31,199,31,95,31,88,31,58,31,211,31,211,30,20,31,14,31,75,31,222,31,222,30,162,31,65,31,176,31,88,31,88,30,46,31,145,31,162,31,164,31,54,31,79,31,54,31,25,31,25,30,142,31,43,31,25,31,5,31,190,31,24,31,24,30,24,29,100,31,122,31,101,31,202,31,74,31,74,30,156,31,73,31,48,31,101,31,103,31,169,31,99,31,74,31,80,31,80,30,80,29,41,31,213,31,56,31,34,31,89,31,115,31,219,31,112,31,80,31,229,31,24,31,24,30,2,31,154,31,154,30,154,29,143,31,141,31,148,31,148,30,193,31,65,31,65,30,202,31,202,30,61,31,188,31,162,31,184,31,124,31,124,30,124,29,124,28,211,31,97,31,229,31,117,31,90,31,130,31,9,31,9,30,158,31,46,31,18,31,151,31,199,31,24,31,182,31,52,31,199,31,20,31,20,30,16,31,16,30,24,31,86,31,103,31,140,31,140,30,204,31,204,30,204,29,255,31,163,31,205,31,158,31,158,30,195,31,3,31,225,31,225,30,240,31,134,31,218,31,218,30,100,31,195,31,100,31,199,31,158,31,206,31,191,31,163,31,151,31,190,31,31,31,180,31,180,31,222,31,27,31,58,31,170,31,96,31,80,31,226,31,212,31,174,31,174,30,174,29,111,31,116,31,170,31,1,31,136,31,20,31,20,30,24,31,73,31,79,31,31,31,31,30,100,31,100,30,135,31,159,31,19,31,38,31,129,31,86,31,198,31,184,31,86,31,168,31,7,31,124,31,247,31,191,31,23,31,23,30,101,31,101,30,101,29,244,31,145,31,23,31,38,31,3,31,234,31,234,30,104,31,104,30,69,31,155,31,220,31,192,31,233,31,102,31,128,31,29,31,105,31,36,31,36,30,36,29,160,31,160,30,160,29,160,31,173,31,20,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
