-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_226 is
end project_tb_226;

architecture project_tb_arch_226 of project_tb_226 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 900;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (52,0,62,0,28,0,5,0,188,0,201,0,15,0,177,0,58,0,57,0,128,0,186,0,48,0,94,0,171,0,0,0,0,0,250,0,0,0,80,0,229,0,27,0,120,0,18,0,238,0,36,0,89,0,255,0,212,0,199,0,0,0,0,0,167,0,141,0,255,0,193,0,101,0,182,0,0,0,204,0,8,0,60,0,132,0,138,0,254,0,131,0,168,0,0,0,27,0,166,0,246,0,0,0,117,0,0,0,126,0,3,0,248,0,97,0,0,0,194,0,44,0,166,0,171,0,19,0,237,0,0,0,125,0,183,0,240,0,74,0,82,0,0,0,105,0,0,0,246,0,96,0,234,0,13,0,98,0,170,0,85,0,173,0,241,0,0,0,214,0,0,0,99,0,216,0,6,0,83,0,246,0,2,0,186,0,0,0,165,0,1,0,183,0,0,0,198,0,215,0,212,0,106,0,0,0,240,0,240,0,50,0,16,0,118,0,16,0,146,0,0,0,210,0,213,0,247,0,25,0,50,0,144,0,0,0,184,0,173,0,204,0,77,0,50,0,0,0,201,0,44,0,11,0,40,0,125,0,79,0,24,0,178,0,0,0,208,0,217,0,239,0,0,0,47,0,58,0,26,0,26,0,0,0,107,0,183,0,151,0,49,0,122,0,20,0,93,0,152,0,0,0,0,0,215,0,40,0,55,0,76,0,89,0,50,0,83,0,75,0,17,0,187,0,28,0,203,0,0,0,0,0,163,0,190,0,0,0,124,0,195,0,0,0,96,0,68,0,202,0,118,0,185,0,48,0,176,0,225,0,216,0,229,0,71,0,62,0,236,0,217,0,214,0,145,0,156,0,3,0,158,0,81,0,236,0,108,0,87,0,187,0,29,0,188,0,0,0,169,0,0,0,0,0,229,0,151,0,0,0,0,0,0,0,127,0,65,0,164,0,162,0,0,0,47,0,200,0,92,0,21,0,0,0,0,0,0,0,87,0,165,0,153,0,168,0,25,0,61,0,19,0,236,0,158,0,171,0,195,0,81,0,24,0,187,0,238,0,0,0,17,0,250,0,0,0,45,0,11,0,44,0,185,0,0,0,0,0,0,0,63,0,58,0,94,0,204,0,134,0,158,0,85,0,163,0,136,0,119,0,112,0,223,0,127,0,0,0,198,0,35,0,0,0,164,0,0,0,174,0,70,0,228,0,0,0,128,0,91,0,33,0,115,0,14,0,237,0,188,0,0,0,0,0,52,0,233,0,0,0,253,0,191,0,145,0,7,0,196,0,0,0,33,0,0,0,158,0,43,0,0,0,0,0,0,0,17,0,164,0,44,0,101,0,213,0,120,0,0,0,0,0,51,0,191,0,66,0,76,0,121,0,0,0,24,0,3,0,155,0,147,0,46,0,115,0,0,0,0,0,5,0,78,0,108,0,238,0,0,0,200,0,169,0,0,0,147,0,195,0,92,0,36,0,42,0,0,0,0,0,151,0,236,0,0,0,139,0,49,0,185,0,117,0,171,0,141,0,124,0,193,0,0,0,115,0,174,0,224,0,0,0,164,0,132,0,238,0,74,0,17,0,6,0,0,0,182,0,176,0,172,0,2,0,246,0,64,0,0,0,109,0,23,0,210,0,24,0,131,0,176,0,100,0,154,0,20,0,97,0,239,0,0,0,150,0,137,0,94,0,147,0,30,0,58,0,140,0,240,0,57,0,35,0,0,0,246,0,249,0,156,0,0,0,202,0,26,0,5,0,31,0,0,0,221,0,42,0,0,0,229,0,40,0,107,0,97,0,62,0,0,0,141,0,117,0,109,0,68,0,178,0,111,0,243,0,0,0,43,0,4,0,112,0,43,0,124,0,15,0,0,0,249,0,150,0,75,0,0,0,176,0,0,0,27,0,224,0,0,0,107,0,243,0,142,0,0,0,5,0,147,0,219,0,0,0,25,0,133,0,70,0,96,0,182,0,47,0,221,0,0,0,0,0,120,0,169,0,0,0,0,0,221,0,209,0,122,0,127,0,83,0,0,0,116,0,0,0,116,0,230,0,148,0,255,0,199,0,43,0,80,0,109,0,14,0,45,0,0,0,233,0,21,0,46,0,60,0,144,0,122,0,37,0,0,0,178,0,0,0,148,0,0,0,1,0,58,0,109,0,32,0,78,0,73,0,254,0,126,0,116,0,73,0,211,0,0,0,118,0,123,0,166,0,0,0,0,0,184,0,104,0,243,0,69,0,0,0,25,0,242,0,239,0,0,0,99,0,0,0,37,0,192,0,99,0,154,0,232,0,137,0,0,0,248,0,0,0,17,0,26,0,0,0,0,0,6,0,15,0,107,0,124,0,225,0,202,0,145,0,13,0,0,0,132,0,150,0,0,0,4,0,219,0,225,0,213,0,0,0,40,0,21,0,0,0,3,0,233,0,0,0,23,0,70,0,96,0,160,0,64,0,78,0,156,0,7,0,52,0,70,0,210,0,26,0,151,0,0,0,244,0,138,0,150,0,100,0,183,0,0,0,0,0,0,0,0,0,0,0,221,0,79,0,35,0,155,0,39,0,184,0,151,0,247,0,96,0,33,0,109,0,193,0,49,0,67,0,0,0,61,0,120,0,0,0,77,0,95,0,207,0,91,0,139,0,44,0,98,0,0,0,173,0,0,0,54,0,183,0,154,0,189,0,0,0,205,0,243,0,249,0,58,0,104,0,0,0,89,0,0,0,88,0,83,0,201,0,243,0,150,0,0,0,205,0,15,0,168,0,0,0,29,0,243,0,112,0,117,0,0,0,194,0,10,0,198,0,147,0,208,0,0,0,32,0,200,0,33,0,79,0,170,0,143,0,148,0,193,0,12,0,251,0,65,0,80,0,0,0,189,0,7,0,75,0,130,0,36,0,0,0,218,0,105,0,16,0,56,0,220,0,171,0,89,0,41,0,54,0,95,0,214,0,24,0,0,0,10,0,0,0,61,0,34,0,54,0,163,0,9,0,1,0,56,0,25,0,146,0,0,0,77,0,1,0,42,0,238,0,0,0,0,0,237,0,0,0,64,0,2,0,110,0,102,0,240,0,4,0,0,0,121,0,0,0,206,0,52,0,231,0,236,0,72,0,37,0,155,0,0,0,167,0,233,0,191,0,71,0,239,0,246,0,0,0,57,0,205,0,176,0,247,0,29,0,0,0,115,0,44,0,79,0,25,0,202,0,40,0,82,0,9,0,11,0,27,0,97,0,15,0,0,0,252,0,224,0,171,0,222,0,0,0,0,0,66,0,117,0,60,0,41,0,6,0,143,0,128,0,0,0,91,0,101,0,250,0,216,0,68,0,111,0,0,0,0,0,0,0,201,0,105,0,0,0,124,0,0,0,94,0,16,0,239,0,0,0,31,0,23,0,21,0,32,0,220,0,0,0,195,0,177,0,0,0,6,0,0,0,106,0,0,0,166,0,0,0,124,0,112,0,53,0,138,0,46,0,104,0,167,0,162,0,0,0,0,0,236,0,0,0,0,0,0,0,183,0,213,0,217,0,0,0,41,0,0,0,218,0,13,0,72,0,43,0,194,0,16,0,169,0,0,0,0,0,139,0,154,0,173,0,0,0,36,0,26,0,206,0,12,0,26,0,188,0,61,0,0,0,0,0,50,0,236,0,118,0,90,0,91,0,167,0,0,0,79,0,204,0,74,0,163,0,194,0,243,0,131,0,0,0,25,0,0,0,0,0,120,0,243,0,251,0,175,0,39,0,246,0,105,0,117,0,118,0,116,0,0,0,237,0,213,0,214,0,135,0,0,0,32,0,63,0,139,0,90,0,144,0,238,0,242,0,151,0,67,0,202,0,200,0,10,0,0,0,0,0,200,0,157,0,33,0,83,0,12,0,3,0,65,0,174,0,190,0,13,0,0,0,190,0,188,0,0,0,180,0,67,0,116,0,79,0,8,0,224,0,201,0,145,0,59,0,27,0,232,0,214,0,148,0,0,0,0,0,140,0,26,0,157,0,230,0,0,0,93,0,3,0,32,0,48,0,52,0,26,0,186,0);
signal scenario_full  : scenario_type := (52,31,62,31,28,31,5,31,188,31,201,31,15,31,177,31,58,31,57,31,128,31,186,31,48,31,94,31,171,31,171,30,171,29,250,31,250,30,80,31,229,31,27,31,120,31,18,31,238,31,36,31,89,31,255,31,212,31,199,31,199,30,199,29,167,31,141,31,255,31,193,31,101,31,182,31,182,30,204,31,8,31,60,31,132,31,138,31,254,31,131,31,168,31,168,30,27,31,166,31,246,31,246,30,117,31,117,30,126,31,3,31,248,31,97,31,97,30,194,31,44,31,166,31,171,31,19,31,237,31,237,30,125,31,183,31,240,31,74,31,82,31,82,30,105,31,105,30,246,31,96,31,234,31,13,31,98,31,170,31,85,31,173,31,241,31,241,30,214,31,214,30,99,31,216,31,6,31,83,31,246,31,2,31,186,31,186,30,165,31,1,31,183,31,183,30,198,31,215,31,212,31,106,31,106,30,240,31,240,31,50,31,16,31,118,31,16,31,146,31,146,30,210,31,213,31,247,31,25,31,50,31,144,31,144,30,184,31,173,31,204,31,77,31,50,31,50,30,201,31,44,31,11,31,40,31,125,31,79,31,24,31,178,31,178,30,208,31,217,31,239,31,239,30,47,31,58,31,26,31,26,31,26,30,107,31,183,31,151,31,49,31,122,31,20,31,93,31,152,31,152,30,152,29,215,31,40,31,55,31,76,31,89,31,50,31,83,31,75,31,17,31,187,31,28,31,203,31,203,30,203,29,163,31,190,31,190,30,124,31,195,31,195,30,96,31,68,31,202,31,118,31,185,31,48,31,176,31,225,31,216,31,229,31,71,31,62,31,236,31,217,31,214,31,145,31,156,31,3,31,158,31,81,31,236,31,108,31,87,31,187,31,29,31,188,31,188,30,169,31,169,30,169,29,229,31,151,31,151,30,151,29,151,28,127,31,65,31,164,31,162,31,162,30,47,31,200,31,92,31,21,31,21,30,21,29,21,28,87,31,165,31,153,31,168,31,25,31,61,31,19,31,236,31,158,31,171,31,195,31,81,31,24,31,187,31,238,31,238,30,17,31,250,31,250,30,45,31,11,31,44,31,185,31,185,30,185,29,185,28,63,31,58,31,94,31,204,31,134,31,158,31,85,31,163,31,136,31,119,31,112,31,223,31,127,31,127,30,198,31,35,31,35,30,164,31,164,30,174,31,70,31,228,31,228,30,128,31,91,31,33,31,115,31,14,31,237,31,188,31,188,30,188,29,52,31,233,31,233,30,253,31,191,31,145,31,7,31,196,31,196,30,33,31,33,30,158,31,43,31,43,30,43,29,43,28,17,31,164,31,44,31,101,31,213,31,120,31,120,30,120,29,51,31,191,31,66,31,76,31,121,31,121,30,24,31,3,31,155,31,147,31,46,31,115,31,115,30,115,29,5,31,78,31,108,31,238,31,238,30,200,31,169,31,169,30,147,31,195,31,92,31,36,31,42,31,42,30,42,29,151,31,236,31,236,30,139,31,49,31,185,31,117,31,171,31,141,31,124,31,193,31,193,30,115,31,174,31,224,31,224,30,164,31,132,31,238,31,74,31,17,31,6,31,6,30,182,31,176,31,172,31,2,31,246,31,64,31,64,30,109,31,23,31,210,31,24,31,131,31,176,31,100,31,154,31,20,31,97,31,239,31,239,30,150,31,137,31,94,31,147,31,30,31,58,31,140,31,240,31,57,31,35,31,35,30,246,31,249,31,156,31,156,30,202,31,26,31,5,31,31,31,31,30,221,31,42,31,42,30,229,31,40,31,107,31,97,31,62,31,62,30,141,31,117,31,109,31,68,31,178,31,111,31,243,31,243,30,43,31,4,31,112,31,43,31,124,31,15,31,15,30,249,31,150,31,75,31,75,30,176,31,176,30,27,31,224,31,224,30,107,31,243,31,142,31,142,30,5,31,147,31,219,31,219,30,25,31,133,31,70,31,96,31,182,31,47,31,221,31,221,30,221,29,120,31,169,31,169,30,169,29,221,31,209,31,122,31,127,31,83,31,83,30,116,31,116,30,116,31,230,31,148,31,255,31,199,31,43,31,80,31,109,31,14,31,45,31,45,30,233,31,21,31,46,31,60,31,144,31,122,31,37,31,37,30,178,31,178,30,148,31,148,30,1,31,58,31,109,31,32,31,78,31,73,31,254,31,126,31,116,31,73,31,211,31,211,30,118,31,123,31,166,31,166,30,166,29,184,31,104,31,243,31,69,31,69,30,25,31,242,31,239,31,239,30,99,31,99,30,37,31,192,31,99,31,154,31,232,31,137,31,137,30,248,31,248,30,17,31,26,31,26,30,26,29,6,31,15,31,107,31,124,31,225,31,202,31,145,31,13,31,13,30,132,31,150,31,150,30,4,31,219,31,225,31,213,31,213,30,40,31,21,31,21,30,3,31,233,31,233,30,23,31,70,31,96,31,160,31,64,31,78,31,156,31,7,31,52,31,70,31,210,31,26,31,151,31,151,30,244,31,138,31,150,31,100,31,183,31,183,30,183,29,183,28,183,27,183,26,221,31,79,31,35,31,155,31,39,31,184,31,151,31,247,31,96,31,33,31,109,31,193,31,49,31,67,31,67,30,61,31,120,31,120,30,77,31,95,31,207,31,91,31,139,31,44,31,98,31,98,30,173,31,173,30,54,31,183,31,154,31,189,31,189,30,205,31,243,31,249,31,58,31,104,31,104,30,89,31,89,30,88,31,83,31,201,31,243,31,150,31,150,30,205,31,15,31,168,31,168,30,29,31,243,31,112,31,117,31,117,30,194,31,10,31,198,31,147,31,208,31,208,30,32,31,200,31,33,31,79,31,170,31,143,31,148,31,193,31,12,31,251,31,65,31,80,31,80,30,189,31,7,31,75,31,130,31,36,31,36,30,218,31,105,31,16,31,56,31,220,31,171,31,89,31,41,31,54,31,95,31,214,31,24,31,24,30,10,31,10,30,61,31,34,31,54,31,163,31,9,31,1,31,56,31,25,31,146,31,146,30,77,31,1,31,42,31,238,31,238,30,238,29,237,31,237,30,64,31,2,31,110,31,102,31,240,31,4,31,4,30,121,31,121,30,206,31,52,31,231,31,236,31,72,31,37,31,155,31,155,30,167,31,233,31,191,31,71,31,239,31,246,31,246,30,57,31,205,31,176,31,247,31,29,31,29,30,115,31,44,31,79,31,25,31,202,31,40,31,82,31,9,31,11,31,27,31,97,31,15,31,15,30,252,31,224,31,171,31,222,31,222,30,222,29,66,31,117,31,60,31,41,31,6,31,143,31,128,31,128,30,91,31,101,31,250,31,216,31,68,31,111,31,111,30,111,29,111,28,201,31,105,31,105,30,124,31,124,30,94,31,16,31,239,31,239,30,31,31,23,31,21,31,32,31,220,31,220,30,195,31,177,31,177,30,6,31,6,30,106,31,106,30,166,31,166,30,124,31,112,31,53,31,138,31,46,31,104,31,167,31,162,31,162,30,162,29,236,31,236,30,236,29,236,28,183,31,213,31,217,31,217,30,41,31,41,30,218,31,13,31,72,31,43,31,194,31,16,31,169,31,169,30,169,29,139,31,154,31,173,31,173,30,36,31,26,31,206,31,12,31,26,31,188,31,61,31,61,30,61,29,50,31,236,31,118,31,90,31,91,31,167,31,167,30,79,31,204,31,74,31,163,31,194,31,243,31,131,31,131,30,25,31,25,30,25,29,120,31,243,31,251,31,175,31,39,31,246,31,105,31,117,31,118,31,116,31,116,30,237,31,213,31,214,31,135,31,135,30,32,31,63,31,139,31,90,31,144,31,238,31,242,31,151,31,67,31,202,31,200,31,10,31,10,30,10,29,200,31,157,31,33,31,83,31,12,31,3,31,65,31,174,31,190,31,13,31,13,30,190,31,188,31,188,30,180,31,67,31,116,31,79,31,8,31,224,31,201,31,145,31,59,31,27,31,232,31,214,31,148,31,148,30,148,29,140,31,26,31,157,31,230,31,230,30,93,31,3,31,32,31,48,31,52,31,26,31,186,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
