-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 906;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (159,0,161,0,123,0,158,0,163,0,132,0,118,0,33,0,87,0,78,0,240,0,0,0,45,0,221,0,180,0,32,0,0,0,0,0,62,0,200,0,181,0,143,0,199,0,195,0,107,0,163,0,0,0,242,0,36,0,0,0,4,0,255,0,135,0,107,0,63,0,55,0,150,0,39,0,243,0,237,0,236,0,88,0,0,0,0,0,90,0,39,0,152,0,97,0,46,0,215,0,117,0,0,0,204,0,160,0,0,0,0,0,0,0,246,0,176,0,0,0,43,0,121,0,20,0,170,0,49,0,0,0,254,0,181,0,93,0,70,0,22,0,174,0,0,0,0,0,223,0,80,0,75,0,88,0,0,0,5,0,78,0,138,0,103,0,228,0,5,0,56,0,0,0,0,0,38,0,105,0,220,0,245,0,2,0,34,0,134,0,65,0,0,0,0,0,159,0,0,0,123,0,151,0,0,0,0,0,133,0,0,0,0,0,0,0,87,0,206,0,113,0,129,0,184,0,210,0,73,0,1,0,42,0,153,0,92,0,116,0,0,0,73,0,0,0,41,0,171,0,126,0,130,0,117,0,39,0,232,0,238,0,206,0,26,0,190,0,180,0,35,0,229,0,0,0,56,0,11,0,225,0,249,0,112,0,207,0,0,0,0,0,6,0,85,0,17,0,193,0,49,0,88,0,104,0,244,0,38,0,134,0,238,0,168,0,33,0,175,0,70,0,0,0,254,0,0,0,118,0,0,0,188,0,60,0,147,0,43,0,109,0,0,0,47,0,49,0,0,0,0,0,203,0,40,0,59,0,0,0,2,0,39,0,78,0,0,0,63,0,0,0,246,0,52,0,244,0,14,0,0,0,37,0,120,0,199,0,0,0,190,0,112,0,211,0,0,0,0,0,5,0,102,0,128,0,212,0,30,0,87,0,87,0,0,0,26,0,1,0,44,0,184,0,11,0,189,0,0,0,0,0,27,0,52,0,72,0,88,0,51,0,0,0,96,0,193,0,159,0,210,0,81,0,0,0,222,0,167,0,38,0,214,0,214,0,19,0,164,0,135,0,12,0,31,0,22,0,20,0,0,0,59,0,8,0,68,0,0,0,49,0,228,0,137,0,156,0,0,0,45,0,24,0,225,0,146,0,10,0,180,0,180,0,19,0,28,0,113,0,102,0,0,0,0,0,214,0,118,0,142,0,107,0,30,0,0,0,210,0,47,0,75,0,0,0,0,0,0,0,59,0,165,0,32,0,229,0,188,0,29,0,190,0,23,0,48,0,98,0,185,0,119,0,251,0,75,0,28,0,152,0,15,0,164,0,93,0,98,0,134,0,207,0,186,0,62,0,14,0,81,0,87,0,120,0,214,0,11,0,0,0,0,0,134,0,83,0,140,0,94,0,34,0,0,0,13,0,36,0,0,0,13,0,12,0,69,0,45,0,205,0,178,0,68,0,235,0,58,0,0,0,0,0,176,0,236,0,62,0,117,0,61,0,0,0,179,0,35,0,0,0,195,0,137,0,45,0,24,0,215,0,0,0,91,0,128,0,113,0,42,0,0,0,49,0,195,0,154,0,156,0,176,0,1,0,0,0,167,0,11,0,82,0,77,0,193,0,236,0,169,0,42,0,206,0,155,0,27,0,146,0,68,0,254,0,128,0,10,0,68,0,0,0,221,0,92,0,104,0,209,0,28,0,35,0,12,0,247,0,0,0,129,0,84,0,90,0,0,0,151,0,84,0,0,0,225,0,0,0,110,0,78,0,47,0,0,0,68,0,211,0,0,0,29,0,246,0,253,0,54,0,43,0,226,0,42,0,102,0,0,0,0,0,41,0,64,0,250,0,0,0,0,0,0,0,127,0,0,0,0,0,15,0,52,0,28,0,23,0,53,0,166,0,245,0,94,0,0,0,91,0,182,0,0,0,154,0,0,0,114,0,175,0,0,0,0,0,30,0,199,0,37,0,86,0,249,0,64,0,227,0,111,0,0,0,235,0,240,0,155,0,46,0,141,0,247,0,198,0,214,0,152,0,87,0,153,0,42,0,182,0,175,0,31,0,181,0,88,0,100,0,118,0,0,0,206,0,152,0,192,0,0,0,12,0,168,0,139,0,184,0,106,0,98,0,0,0,0,0,0,0,249,0,234,0,0,0,0,0,0,0,232,0,0,0,57,0,68,0,117,0,43,0,108,0,0,0,46,0,0,0,17,0,0,0,37,0,4,0,170,0,176,0,25,0,169,0,0,0,219,0,26,0,223,0,98,0,113,0,94,0,0,0,0,0,209,0,211,0,132,0,0,0,121,0,108,0,23,0,0,0,190,0,201,0,79,0,196,0,0,0,89,0,101,0,0,0,0,0,4,0,168,0,18,0,131,0,209,0,243,0,4,0,185,0,49,0,0,0,168,0,150,0,197,0,104,0,164,0,149,0,222,0,198,0,120,0,237,0,8,0,76,0,216,0,28,0,119,0,96,0,238,0,0,0,239,0,117,0,236,0,0,0,172,0,34,0,54,0,166,0,86,0,212,0,83,0,242,0,0,0,243,0,0,0,0,0,228,0,5,0,0,0,0,0,52,0,0,0,135,0,100,0,180,0,92,0,254,0,35,0,64,0,0,0,48,0,105,0,0,0,74,0,182,0,0,0,239,0,130,0,103,0,176,0,225,0,253,0,76,0,44,0,6,0,0,0,191,0,37,0,73,0,214,0,236,0,180,0,230,0,34,0,109,0,132,0,179,0,0,0,21,0,0,0,198,0,94,0,75,0,50,0,0,0,96,0,185,0,240,0,118,0,0,0,47,0,200,0,145,0,203,0,143,0,207,0,0,0,19,0,0,0,171,0,53,0,173,0,147,0,103,0,172,0,167,0,20,0,124,0,54,0,0,0,109,0,239,0,9,0,206,0,15,0,207,0,103,0,0,0,186,0,0,0,180,0,48,0,107,0,16,0,60,0,34,0,103,0,144,0,0,0,71,0,51,0,0,0,46,0,29,0,200,0,0,0,205,0,205,0,126,0,0,0,244,0,54,0,169,0,100,0,151,0,0,0,240,0,148,0,119,0,65,0,0,0,0,0,188,0,196,0,36,0,227,0,156,0,0,0,0,0,220,0,0,0,0,0,243,0,103,0,0,0,0,0,161,0,62,0,0,0,10,0,68,0,162,0,106,0,167,0,0,0,179,0,124,0,134,0,164,0,12,0,227,0,0,0,130,0,120,0,164,0,164,0,0,0,212,0,41,0,108,0,0,0,48,0,0,0,217,0,106,0,0,0,175,0,236,0,0,0,172,0,171,0,0,0,0,0,208,0,0,0,180,0,68,0,127,0,213,0,203,0,32,0,0,0,4,0,26,0,205,0,148,0,143,0,0,0,156,0,239,0,94,0,56,0,203,0,215,0,0,0,75,0,93,0,159,0,73,0,173,0,142,0,13,0,167,0,81,0,231,0,145,0,31,0,27,0,0,0,30,0,175,0,222,0,43,0,110,0,39,0,0,0,132,0,0,0,115,0,116,0,113,0,42,0,82,0,0,0,141,0,45,0,230,0,202,0,27,0,116,0,0,0,223,0,79,0,212,0,0,0,164,0,99,0,0,0,102,0,55,0,76,0,70,0,187,0,56,0,0,0,193,0,49,0,211,0,115,0,62,0,60,0,49,0,14,0,93,0,62,0,230,0,39,0,0,0,160,0,140,0,0,0,25,0,15,0,100,0,96,0,0,0,172,0,253,0,76,0,174,0,194,0,0,0,0,0,0,0,192,0,238,0,157,0,69,0,24,0,150,0,0,0,233,0,36,0,167,0,110,0,31,0,0,0,51,0,44,0,0,0,83,0,0,0,17,0,7,0,0,0,131,0,179,0,33,0,0,0,231,0,183,0,83,0,65,0,0,0,251,0,105,0,35,0,20,0,225,0,242,0,200,0,82,0,36,0,0,0,227,0,211,0,243,0,12,0,144,0,0,0,40,0,4,0,237,0,0,0,0,0,53,0,0,0,177,0,0,0,5,0,0,0,193,0,91,0,0,0,0,0,81,0,0,0,74,0,84,0,145,0,106,0,201,0,149,0);
signal scenario_full  : scenario_type := (159,31,161,31,123,31,158,31,163,31,132,31,118,31,33,31,87,31,78,31,240,31,240,30,45,31,221,31,180,31,32,31,32,30,32,29,62,31,200,31,181,31,143,31,199,31,195,31,107,31,163,31,163,30,242,31,36,31,36,30,4,31,255,31,135,31,107,31,63,31,55,31,150,31,39,31,243,31,237,31,236,31,88,31,88,30,88,29,90,31,39,31,152,31,97,31,46,31,215,31,117,31,117,30,204,31,160,31,160,30,160,29,160,28,246,31,176,31,176,30,43,31,121,31,20,31,170,31,49,31,49,30,254,31,181,31,93,31,70,31,22,31,174,31,174,30,174,29,223,31,80,31,75,31,88,31,88,30,5,31,78,31,138,31,103,31,228,31,5,31,56,31,56,30,56,29,38,31,105,31,220,31,245,31,2,31,34,31,134,31,65,31,65,30,65,29,159,31,159,30,123,31,151,31,151,30,151,29,133,31,133,30,133,29,133,28,87,31,206,31,113,31,129,31,184,31,210,31,73,31,1,31,42,31,153,31,92,31,116,31,116,30,73,31,73,30,41,31,171,31,126,31,130,31,117,31,39,31,232,31,238,31,206,31,26,31,190,31,180,31,35,31,229,31,229,30,56,31,11,31,225,31,249,31,112,31,207,31,207,30,207,29,6,31,85,31,17,31,193,31,49,31,88,31,104,31,244,31,38,31,134,31,238,31,168,31,33,31,175,31,70,31,70,30,254,31,254,30,118,31,118,30,188,31,60,31,147,31,43,31,109,31,109,30,47,31,49,31,49,30,49,29,203,31,40,31,59,31,59,30,2,31,39,31,78,31,78,30,63,31,63,30,246,31,52,31,244,31,14,31,14,30,37,31,120,31,199,31,199,30,190,31,112,31,211,31,211,30,211,29,5,31,102,31,128,31,212,31,30,31,87,31,87,31,87,30,26,31,1,31,44,31,184,31,11,31,189,31,189,30,189,29,27,31,52,31,72,31,88,31,51,31,51,30,96,31,193,31,159,31,210,31,81,31,81,30,222,31,167,31,38,31,214,31,214,31,19,31,164,31,135,31,12,31,31,31,22,31,20,31,20,30,59,31,8,31,68,31,68,30,49,31,228,31,137,31,156,31,156,30,45,31,24,31,225,31,146,31,10,31,180,31,180,31,19,31,28,31,113,31,102,31,102,30,102,29,214,31,118,31,142,31,107,31,30,31,30,30,210,31,47,31,75,31,75,30,75,29,75,28,59,31,165,31,32,31,229,31,188,31,29,31,190,31,23,31,48,31,98,31,185,31,119,31,251,31,75,31,28,31,152,31,15,31,164,31,93,31,98,31,134,31,207,31,186,31,62,31,14,31,81,31,87,31,120,31,214,31,11,31,11,30,11,29,134,31,83,31,140,31,94,31,34,31,34,30,13,31,36,31,36,30,13,31,12,31,69,31,45,31,205,31,178,31,68,31,235,31,58,31,58,30,58,29,176,31,236,31,62,31,117,31,61,31,61,30,179,31,35,31,35,30,195,31,137,31,45,31,24,31,215,31,215,30,91,31,128,31,113,31,42,31,42,30,49,31,195,31,154,31,156,31,176,31,1,31,1,30,167,31,11,31,82,31,77,31,193,31,236,31,169,31,42,31,206,31,155,31,27,31,146,31,68,31,254,31,128,31,10,31,68,31,68,30,221,31,92,31,104,31,209,31,28,31,35,31,12,31,247,31,247,30,129,31,84,31,90,31,90,30,151,31,84,31,84,30,225,31,225,30,110,31,78,31,47,31,47,30,68,31,211,31,211,30,29,31,246,31,253,31,54,31,43,31,226,31,42,31,102,31,102,30,102,29,41,31,64,31,250,31,250,30,250,29,250,28,127,31,127,30,127,29,15,31,52,31,28,31,23,31,53,31,166,31,245,31,94,31,94,30,91,31,182,31,182,30,154,31,154,30,114,31,175,31,175,30,175,29,30,31,199,31,37,31,86,31,249,31,64,31,227,31,111,31,111,30,235,31,240,31,155,31,46,31,141,31,247,31,198,31,214,31,152,31,87,31,153,31,42,31,182,31,175,31,31,31,181,31,88,31,100,31,118,31,118,30,206,31,152,31,192,31,192,30,12,31,168,31,139,31,184,31,106,31,98,31,98,30,98,29,98,28,249,31,234,31,234,30,234,29,234,28,232,31,232,30,57,31,68,31,117,31,43,31,108,31,108,30,46,31,46,30,17,31,17,30,37,31,4,31,170,31,176,31,25,31,169,31,169,30,219,31,26,31,223,31,98,31,113,31,94,31,94,30,94,29,209,31,211,31,132,31,132,30,121,31,108,31,23,31,23,30,190,31,201,31,79,31,196,31,196,30,89,31,101,31,101,30,101,29,4,31,168,31,18,31,131,31,209,31,243,31,4,31,185,31,49,31,49,30,168,31,150,31,197,31,104,31,164,31,149,31,222,31,198,31,120,31,237,31,8,31,76,31,216,31,28,31,119,31,96,31,238,31,238,30,239,31,117,31,236,31,236,30,172,31,34,31,54,31,166,31,86,31,212,31,83,31,242,31,242,30,243,31,243,30,243,29,228,31,5,31,5,30,5,29,52,31,52,30,135,31,100,31,180,31,92,31,254,31,35,31,64,31,64,30,48,31,105,31,105,30,74,31,182,31,182,30,239,31,130,31,103,31,176,31,225,31,253,31,76,31,44,31,6,31,6,30,191,31,37,31,73,31,214,31,236,31,180,31,230,31,34,31,109,31,132,31,179,31,179,30,21,31,21,30,198,31,94,31,75,31,50,31,50,30,96,31,185,31,240,31,118,31,118,30,47,31,200,31,145,31,203,31,143,31,207,31,207,30,19,31,19,30,171,31,53,31,173,31,147,31,103,31,172,31,167,31,20,31,124,31,54,31,54,30,109,31,239,31,9,31,206,31,15,31,207,31,103,31,103,30,186,31,186,30,180,31,48,31,107,31,16,31,60,31,34,31,103,31,144,31,144,30,71,31,51,31,51,30,46,31,29,31,200,31,200,30,205,31,205,31,126,31,126,30,244,31,54,31,169,31,100,31,151,31,151,30,240,31,148,31,119,31,65,31,65,30,65,29,188,31,196,31,36,31,227,31,156,31,156,30,156,29,220,31,220,30,220,29,243,31,103,31,103,30,103,29,161,31,62,31,62,30,10,31,68,31,162,31,106,31,167,31,167,30,179,31,124,31,134,31,164,31,12,31,227,31,227,30,130,31,120,31,164,31,164,31,164,30,212,31,41,31,108,31,108,30,48,31,48,30,217,31,106,31,106,30,175,31,236,31,236,30,172,31,171,31,171,30,171,29,208,31,208,30,180,31,68,31,127,31,213,31,203,31,32,31,32,30,4,31,26,31,205,31,148,31,143,31,143,30,156,31,239,31,94,31,56,31,203,31,215,31,215,30,75,31,93,31,159,31,73,31,173,31,142,31,13,31,167,31,81,31,231,31,145,31,31,31,27,31,27,30,30,31,175,31,222,31,43,31,110,31,39,31,39,30,132,31,132,30,115,31,116,31,113,31,42,31,82,31,82,30,141,31,45,31,230,31,202,31,27,31,116,31,116,30,223,31,79,31,212,31,212,30,164,31,99,31,99,30,102,31,55,31,76,31,70,31,187,31,56,31,56,30,193,31,49,31,211,31,115,31,62,31,60,31,49,31,14,31,93,31,62,31,230,31,39,31,39,30,160,31,140,31,140,30,25,31,15,31,100,31,96,31,96,30,172,31,253,31,76,31,174,31,194,31,194,30,194,29,194,28,192,31,238,31,157,31,69,31,24,31,150,31,150,30,233,31,36,31,167,31,110,31,31,31,31,30,51,31,44,31,44,30,83,31,83,30,17,31,7,31,7,30,131,31,179,31,33,31,33,30,231,31,183,31,83,31,65,31,65,30,251,31,105,31,35,31,20,31,225,31,242,31,200,31,82,31,36,31,36,30,227,31,211,31,243,31,12,31,144,31,144,30,40,31,4,31,237,31,237,30,237,29,53,31,53,30,177,31,177,30,5,31,5,30,193,31,91,31,91,30,91,29,81,31,81,30,74,31,84,31,145,31,106,31,201,31,149,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
