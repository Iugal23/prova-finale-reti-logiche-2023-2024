-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 399;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,18,0,0,0,94,0,154,0,91,0,180,0,46,0,4,0,24,0,242,0,87,0,156,0,130,0,244,0,126,0,126,0,251,0,0,0,175,0,68,0,16,0,220,0,0,0,0,0,141,0,255,0,190,0,202,0,120,0,21,0,167,0,143,0,201,0,178,0,108,0,91,0,45,0,0,0,0,0,155,0,147,0,75,0,240,0,232,0,0,0,196,0,242,0,0,0,216,0,142,0,130,0,201,0,247,0,0,0,102,0,0,0,3,0,91,0,99,0,52,0,97,0,14,0,202,0,83,0,0,0,229,0,60,0,0,0,0,0,0,0,208,0,131,0,34,0,73,0,245,0,95,0,52,0,77,0,225,0,0,0,0,0,191,0,160,0,65,0,0,0,252,0,75,0,109,0,2,0,113,0,0,0,194,0,143,0,14,0,127,0,25,0,233,0,29,0,230,0,201,0,52,0,125,0,0,0,77,0,0,0,112,0,166,0,159,0,143,0,14,0,242,0,56,0,184,0,223,0,0,0,0,0,159,0,0,0,158,0,224,0,0,0,44,0,60,0,254,0,190,0,166,0,162,0,0,0,56,0,198,0,241,0,153,0,0,0,0,0,240,0,0,0,26,0,0,0,70,0,205,0,218,0,135,0,84,0,158,0,0,0,0,0,159,0,179,0,250,0,0,0,0,0,227,0,190,0,107,0,33,0,0,0,92,0,106,0,112,0,231,0,134,0,47,0,154,0,11,0,192,0,45,0,83,0,32,0,203,0,85,0,236,0,191,0,195,0,224,0,0,0,134,0,129,0,244,0,48,0,120,0,82,0,0,0,28,0,58,0,99,0,211,0,189,0,57,0,0,0,96,0,218,0,116,0,160,0,0,0,0,0,82,0,0,0,134,0,0,0,0,0,0,0,129,0,41,0,43,0,183,0,209,0,157,0,191,0,122,0,53,0,3,0,153,0,0,0,0,0,100,0,8,0,134,0,168,0,67,0,116,0,155,0,76,0,44,0,0,0,210,0,217,0,150,0,0,0,117,0,215,0,109,0,114,0,101,0,47,0,140,0,122,0,64,0,211,0,68,0,127,0,0,0,214,0,148,0,10,0,0,0,161,0,0,0,6,0,184,0,40,0,145,0,95,0,108,0,168,0,74,0,246,0,3,0,4,0,90,0,1,0,10,0,252,0,159,0,221,0,118,0,106,0,54,0,232,0,0,0,215,0,195,0,190,0,196,0,109,0,169,0,223,0,177,0,90,0,28,0,43,0,48,0,195,0,238,0,41,0,51,0,48,0,240,0,161,0,116,0,91,0,94,0,0,0,75,0,0,0,0,0,245,0,163,0,17,0,108,0,0,0,5,0,219,0,0,0,0,0,133,0,142,0,0,0,162,0,199,0,204,0,169,0,20,0,1,0,209,0,27,0,208,0,81,0,203,0,220,0,8,0,70,0,172,0,53,0,129,0,64,0,59,0,22,0,59,0,161,0,0,0,0,0,89,0,124,0,186,0,0,0,37,0,229,0,0,0,22,0,146,0,99,0,66,0,38,0,126,0,165,0,77,0,0,0,83,0,78,0,43,0,98,0,81,0,148,0,100,0,0,0,6,0,241,0,0,0,227,0,175,0,66,0,109,0,148,0,221,0,47,0,71,0,0,0,1,0,87,0,143,0,141,0,0,0,14,0,0,0,104,0,11,0,165,0,70,0,242,0,125,0,207,0,185,0,0,0,0,0,52,0,109,0,111,0,251,0,0,0,219,0,0,0,181,0,83,0,106,0,0,0,26,0,183,0,0,0);
signal scenario_full  : scenario_type := (0,0,18,31,18,30,94,31,154,31,91,31,180,31,46,31,4,31,24,31,242,31,87,31,156,31,130,31,244,31,126,31,126,31,251,31,251,30,175,31,68,31,16,31,220,31,220,30,220,29,141,31,255,31,190,31,202,31,120,31,21,31,167,31,143,31,201,31,178,31,108,31,91,31,45,31,45,30,45,29,155,31,147,31,75,31,240,31,232,31,232,30,196,31,242,31,242,30,216,31,142,31,130,31,201,31,247,31,247,30,102,31,102,30,3,31,91,31,99,31,52,31,97,31,14,31,202,31,83,31,83,30,229,31,60,31,60,30,60,29,60,28,208,31,131,31,34,31,73,31,245,31,95,31,52,31,77,31,225,31,225,30,225,29,191,31,160,31,65,31,65,30,252,31,75,31,109,31,2,31,113,31,113,30,194,31,143,31,14,31,127,31,25,31,233,31,29,31,230,31,201,31,52,31,125,31,125,30,77,31,77,30,112,31,166,31,159,31,143,31,14,31,242,31,56,31,184,31,223,31,223,30,223,29,159,31,159,30,158,31,224,31,224,30,44,31,60,31,254,31,190,31,166,31,162,31,162,30,56,31,198,31,241,31,153,31,153,30,153,29,240,31,240,30,26,31,26,30,70,31,205,31,218,31,135,31,84,31,158,31,158,30,158,29,159,31,179,31,250,31,250,30,250,29,227,31,190,31,107,31,33,31,33,30,92,31,106,31,112,31,231,31,134,31,47,31,154,31,11,31,192,31,45,31,83,31,32,31,203,31,85,31,236,31,191,31,195,31,224,31,224,30,134,31,129,31,244,31,48,31,120,31,82,31,82,30,28,31,58,31,99,31,211,31,189,31,57,31,57,30,96,31,218,31,116,31,160,31,160,30,160,29,82,31,82,30,134,31,134,30,134,29,134,28,129,31,41,31,43,31,183,31,209,31,157,31,191,31,122,31,53,31,3,31,153,31,153,30,153,29,100,31,8,31,134,31,168,31,67,31,116,31,155,31,76,31,44,31,44,30,210,31,217,31,150,31,150,30,117,31,215,31,109,31,114,31,101,31,47,31,140,31,122,31,64,31,211,31,68,31,127,31,127,30,214,31,148,31,10,31,10,30,161,31,161,30,6,31,184,31,40,31,145,31,95,31,108,31,168,31,74,31,246,31,3,31,4,31,90,31,1,31,10,31,252,31,159,31,221,31,118,31,106,31,54,31,232,31,232,30,215,31,195,31,190,31,196,31,109,31,169,31,223,31,177,31,90,31,28,31,43,31,48,31,195,31,238,31,41,31,51,31,48,31,240,31,161,31,116,31,91,31,94,31,94,30,75,31,75,30,75,29,245,31,163,31,17,31,108,31,108,30,5,31,219,31,219,30,219,29,133,31,142,31,142,30,162,31,199,31,204,31,169,31,20,31,1,31,209,31,27,31,208,31,81,31,203,31,220,31,8,31,70,31,172,31,53,31,129,31,64,31,59,31,22,31,59,31,161,31,161,30,161,29,89,31,124,31,186,31,186,30,37,31,229,31,229,30,22,31,146,31,99,31,66,31,38,31,126,31,165,31,77,31,77,30,83,31,78,31,43,31,98,31,81,31,148,31,100,31,100,30,6,31,241,31,241,30,227,31,175,31,66,31,109,31,148,31,221,31,47,31,71,31,71,30,1,31,87,31,143,31,141,31,141,30,14,31,14,30,104,31,11,31,165,31,70,31,242,31,125,31,207,31,185,31,185,30,185,29,52,31,109,31,111,31,251,31,251,30,219,31,219,30,181,31,83,31,106,31,106,30,26,31,183,31,183,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
