-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 807;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (241,0,0,0,109,0,45,0,87,0,14,0,249,0,180,0,10,0,145,0,0,0,0,0,17,0,164,0,255,0,0,0,0,0,0,0,135,0,49,0,224,0,251,0,216,0,160,0,121,0,185,0,214,0,128,0,63,0,236,0,254,0,253,0,88,0,255,0,0,0,0,0,57,0,167,0,197,0,96,0,86,0,108,0,7,0,194,0,4,0,235,0,42,0,179,0,87,0,125,0,116,0,0,0,4,0,0,0,10,0,11,0,47,0,129,0,68,0,61,0,71,0,137,0,5,0,159,0,224,0,0,0,0,0,25,0,0,0,16,0,0,0,225,0,191,0,223,0,68,0,0,0,138,0,133,0,157,0,196,0,155,0,217,0,217,0,253,0,102,0,166,0,68,0,44,0,167,0,224,0,52,0,0,0,54,0,52,0,183,0,206,0,9,0,219,0,252,0,17,0,0,0,0,0,105,0,191,0,45,0,60,0,183,0,134,0,172,0,144,0,152,0,148,0,69,0,0,0,117,0,98,0,26,0,209,0,40,0,134,0,141,0,16,0,114,0,236,0,222,0,191,0,129,0,84,0,82,0,42,0,87,0,237,0,148,0,224,0,74,0,203,0,133,0,130,0,129,0,21,0,255,0,0,0,217,0,0,0,14,0,114,0,101,0,202,0,0,0,79,0,0,0,158,0,67,0,7,0,0,0,1,0,0,0,0,0,18,0,0,0,0,0,99,0,232,0,5,0,0,0,214,0,59,0,14,0,66,0,80,0,176,0,0,0,76,0,79,0,198,0,131,0,217,0,157,0,73,0,232,0,132,0,163,0,0,0,1,0,123,0,223,0,142,0,226,0,251,0,34,0,174,0,45,0,216,0,0,0,0,0,103,0,160,0,0,0,128,0,0,0,0,0,119,0,59,0,104,0,8,0,123,0,35,0,53,0,41,0,193,0,215,0,135,0,91,0,26,0,195,0,48,0,206,0,62,0,192,0,192,0,159,0,52,0,0,0,36,0,208,0,135,0,75,0,215,0,249,0,193,0,177,0,182,0,132,0,48,0,175,0,88,0,173,0,0,0,116,0,0,0,245,0,210,0,49,0,38,0,146,0,103,0,0,0,150,0,195,0,127,0,48,0,16,0,155,0,0,0,175,0,0,0,71,0,0,0,191,0,0,0,80,0,103,0,76,0,215,0,73,0,45,0,178,0,64,0,152,0,138,0,105,0,231,0,0,0,0,0,110,0,134,0,161,0,197,0,175,0,158,0,214,0,0,0,142,0,230,0,215,0,76,0,224,0,100,0,233,0,74,0,127,0,157,0,0,0,111,0,0,0,180,0,0,0,92,0,0,0,101,0,65,0,160,0,151,0,0,0,181,0,203,0,219,0,116,0,133,0,0,0,71,0,149,0,0,0,66,0,0,0,0,0,251,0,191,0,14,0,115,0,169,0,204,0,148,0,208,0,0,0,64,0,182,0,159,0,77,0,47,0,0,0,199,0,65,0,0,0,69,0,142,0,119,0,223,0,147,0,72,0,227,0,88,0,165,0,213,0,107,0,0,0,0,0,115,0,75,0,118,0,0,0,30,0,94,0,99,0,74,0,0,0,58,0,100,0,199,0,249,0,0,0,205,0,42,0,23,0,132,0,37,0,59,0,150,0,214,0,163,0,33,0,139,0,57,0,12,0,0,0,49,0,44,0,229,0,250,0,84,0,53,0,32,0,80,0,192,0,86,0,24,0,222,0,42,0,202,0,28,0,22,0,91,0,70,0,0,0,84,0,150,0,211,0,186,0,94,0,5,0,21,0,228,0,30,0,159,0,0,0,230,0,21,0,178,0,35,0,126,0,97,0,0,0,25,0,107,0,208,0,93,0,125,0,24,0,70,0,100,0,148,0,0,0,105,0,0,0,203,0,22,0,95,0,139,0,115,0,89,0,0,0,78,0,98,0,97,0,122,0,226,0,226,0,32,0,192,0,244,0,0,0,218,0,169,0,52,0,26,0,13,0,69,0,206,0,141,0,57,0,22,0,1,0,160,0,0,0,96,0,147,0,40,0,236,0,244,0,159,0,180,0,199,0,3,0,65,0,0,0,0,0,0,0,95,0,181,0,206,0,36,0,246,0,56,0,166,0,0,0,10,0,139,0,245,0,161,0,82,0,90,0,15,0,89,0,248,0,210,0,47,0,133,0,0,0,0,0,111,0,252,0,241,0,0,0,0,0,173,0,190,0,56,0,178,0,0,0,237,0,168,0,190,0,22,0,202,0,92,0,0,0,91,0,0,0,35,0,255,0,125,0,189,0,189,0,211,0,227,0,250,0,98,0,187,0,129,0,248,0,86,0,71,0,132,0,153,0,17,0,160,0,30,0,179,0,95,0,248,0,245,0,40,0,164,0,126,0,234,0,174,0,0,0,78,0,139,0,23,0,159,0,109,0,46,0,0,0,147,0,147,0,143,0,30,0,105,0,227,0,220,0,8,0,110,0,122,0,0,0,246,0,145,0,18,0,0,0,207,0,194,0,125,0,173,0,208,0,0,0,0,0,240,0,66,0,175,0,0,0,0,0,106,0,196,0,112,0,214,0,202,0,0,0,0,0,225,0,179,0,113,0,0,0,8,0,135,0,14,0,71,0,0,0,194,0,7,0,255,0,119,0,39,0,61,0,55,0,0,0,50,0,32,0,0,0,244,0,164,0,94,0,114,0,0,0,79,0,70,0,25,0,84,0,14,0,157,0,134,0,123,0,167,0,190,0,43,0,72,0,197,0,0,0,123,0,71,0,137,0,27,0,40,0,6,0,254,0,0,0,55,0,160,0,27,0,192,0,251,0,0,0,0,0,91,0,137,0,239,0,0,0,246,0,136,0,11,0,0,0,50,0,0,0,87,0,65,0,36,0,125,0,70,0,0,0,234,0,194,0,45,0,89,0,72,0,221,0,84,0,244,0,116,0,236,0,0,0,5,0,106,0,251,0,174,0,40,0,209,0,243,0,249,0,0,0,181,0,34,0,69,0,84,0,13,0,222,0,40,0,229,0,212,0,130,0,211,0,0,0,79,0,0,0,26,0,191,0,0,0,0,0,5,0,252,0,111,0,253,0,78,0,254,0,8,0,84,0,0,0,0,0,249,0,0,0,130,0,0,0,72,0,195,0,107,0,110,0,12,0,236,0,0,0,218,0,163,0,84,0,46,0,126,0,221,0,15,0,75,0,246,0,175,0,46,0,60,0,47,0,199,0,0,0,146,0,42,0,201,0,235,0,0,0,142,0,0,0,98,0,137,0,162,0,108,0,209,0,8,0,231,0,51,0,0,0,139,0,104,0,10,0,141,0,102,0,235,0,96,0,122,0,0,0,132,0,126,0,135,0,133,0,214,0,145,0,167,0,109,0,39,0,58,0,180,0,180,0,191,0,122,0,246,0,15,0,151,0,94,0,248,0,0,0,123,0,0,0,127,0,236,0,125,0,0,0,234,0,0,0,143,0,0,0,188,0,0,0,162,0,0,0,23,0,0,0,56,0,250,0,92,0,55,0,121,0,82,0,25,0,55,0,0,0,232,0,0,0,67,0,20,0,107,0,67,0,131,0,185,0,1,0,50,0,178,0,151,0,0,0,2,0,64,0);
signal scenario_full  : scenario_type := (241,31,241,30,109,31,45,31,87,31,14,31,249,31,180,31,10,31,145,31,145,30,145,29,17,31,164,31,255,31,255,30,255,29,255,28,135,31,49,31,224,31,251,31,216,31,160,31,121,31,185,31,214,31,128,31,63,31,236,31,254,31,253,31,88,31,255,31,255,30,255,29,57,31,167,31,197,31,96,31,86,31,108,31,7,31,194,31,4,31,235,31,42,31,179,31,87,31,125,31,116,31,116,30,4,31,4,30,10,31,11,31,47,31,129,31,68,31,61,31,71,31,137,31,5,31,159,31,224,31,224,30,224,29,25,31,25,30,16,31,16,30,225,31,191,31,223,31,68,31,68,30,138,31,133,31,157,31,196,31,155,31,217,31,217,31,253,31,102,31,166,31,68,31,44,31,167,31,224,31,52,31,52,30,54,31,52,31,183,31,206,31,9,31,219,31,252,31,17,31,17,30,17,29,105,31,191,31,45,31,60,31,183,31,134,31,172,31,144,31,152,31,148,31,69,31,69,30,117,31,98,31,26,31,209,31,40,31,134,31,141,31,16,31,114,31,236,31,222,31,191,31,129,31,84,31,82,31,42,31,87,31,237,31,148,31,224,31,74,31,203,31,133,31,130,31,129,31,21,31,255,31,255,30,217,31,217,30,14,31,114,31,101,31,202,31,202,30,79,31,79,30,158,31,67,31,7,31,7,30,1,31,1,30,1,29,18,31,18,30,18,29,99,31,232,31,5,31,5,30,214,31,59,31,14,31,66,31,80,31,176,31,176,30,76,31,79,31,198,31,131,31,217,31,157,31,73,31,232,31,132,31,163,31,163,30,1,31,123,31,223,31,142,31,226,31,251,31,34,31,174,31,45,31,216,31,216,30,216,29,103,31,160,31,160,30,128,31,128,30,128,29,119,31,59,31,104,31,8,31,123,31,35,31,53,31,41,31,193,31,215,31,135,31,91,31,26,31,195,31,48,31,206,31,62,31,192,31,192,31,159,31,52,31,52,30,36,31,208,31,135,31,75,31,215,31,249,31,193,31,177,31,182,31,132,31,48,31,175,31,88,31,173,31,173,30,116,31,116,30,245,31,210,31,49,31,38,31,146,31,103,31,103,30,150,31,195,31,127,31,48,31,16,31,155,31,155,30,175,31,175,30,71,31,71,30,191,31,191,30,80,31,103,31,76,31,215,31,73,31,45,31,178,31,64,31,152,31,138,31,105,31,231,31,231,30,231,29,110,31,134,31,161,31,197,31,175,31,158,31,214,31,214,30,142,31,230,31,215,31,76,31,224,31,100,31,233,31,74,31,127,31,157,31,157,30,111,31,111,30,180,31,180,30,92,31,92,30,101,31,65,31,160,31,151,31,151,30,181,31,203,31,219,31,116,31,133,31,133,30,71,31,149,31,149,30,66,31,66,30,66,29,251,31,191,31,14,31,115,31,169,31,204,31,148,31,208,31,208,30,64,31,182,31,159,31,77,31,47,31,47,30,199,31,65,31,65,30,69,31,142,31,119,31,223,31,147,31,72,31,227,31,88,31,165,31,213,31,107,31,107,30,107,29,115,31,75,31,118,31,118,30,30,31,94,31,99,31,74,31,74,30,58,31,100,31,199,31,249,31,249,30,205,31,42,31,23,31,132,31,37,31,59,31,150,31,214,31,163,31,33,31,139,31,57,31,12,31,12,30,49,31,44,31,229,31,250,31,84,31,53,31,32,31,80,31,192,31,86,31,24,31,222,31,42,31,202,31,28,31,22,31,91,31,70,31,70,30,84,31,150,31,211,31,186,31,94,31,5,31,21,31,228,31,30,31,159,31,159,30,230,31,21,31,178,31,35,31,126,31,97,31,97,30,25,31,107,31,208,31,93,31,125,31,24,31,70,31,100,31,148,31,148,30,105,31,105,30,203,31,22,31,95,31,139,31,115,31,89,31,89,30,78,31,98,31,97,31,122,31,226,31,226,31,32,31,192,31,244,31,244,30,218,31,169,31,52,31,26,31,13,31,69,31,206,31,141,31,57,31,22,31,1,31,160,31,160,30,96,31,147,31,40,31,236,31,244,31,159,31,180,31,199,31,3,31,65,31,65,30,65,29,65,28,95,31,181,31,206,31,36,31,246,31,56,31,166,31,166,30,10,31,139,31,245,31,161,31,82,31,90,31,15,31,89,31,248,31,210,31,47,31,133,31,133,30,133,29,111,31,252,31,241,31,241,30,241,29,173,31,190,31,56,31,178,31,178,30,237,31,168,31,190,31,22,31,202,31,92,31,92,30,91,31,91,30,35,31,255,31,125,31,189,31,189,31,211,31,227,31,250,31,98,31,187,31,129,31,248,31,86,31,71,31,132,31,153,31,17,31,160,31,30,31,179,31,95,31,248,31,245,31,40,31,164,31,126,31,234,31,174,31,174,30,78,31,139,31,23,31,159,31,109,31,46,31,46,30,147,31,147,31,143,31,30,31,105,31,227,31,220,31,8,31,110,31,122,31,122,30,246,31,145,31,18,31,18,30,207,31,194,31,125,31,173,31,208,31,208,30,208,29,240,31,66,31,175,31,175,30,175,29,106,31,196,31,112,31,214,31,202,31,202,30,202,29,225,31,179,31,113,31,113,30,8,31,135,31,14,31,71,31,71,30,194,31,7,31,255,31,119,31,39,31,61,31,55,31,55,30,50,31,32,31,32,30,244,31,164,31,94,31,114,31,114,30,79,31,70,31,25,31,84,31,14,31,157,31,134,31,123,31,167,31,190,31,43,31,72,31,197,31,197,30,123,31,71,31,137,31,27,31,40,31,6,31,254,31,254,30,55,31,160,31,27,31,192,31,251,31,251,30,251,29,91,31,137,31,239,31,239,30,246,31,136,31,11,31,11,30,50,31,50,30,87,31,65,31,36,31,125,31,70,31,70,30,234,31,194,31,45,31,89,31,72,31,221,31,84,31,244,31,116,31,236,31,236,30,5,31,106,31,251,31,174,31,40,31,209,31,243,31,249,31,249,30,181,31,34,31,69,31,84,31,13,31,222,31,40,31,229,31,212,31,130,31,211,31,211,30,79,31,79,30,26,31,191,31,191,30,191,29,5,31,252,31,111,31,253,31,78,31,254,31,8,31,84,31,84,30,84,29,249,31,249,30,130,31,130,30,72,31,195,31,107,31,110,31,12,31,236,31,236,30,218,31,163,31,84,31,46,31,126,31,221,31,15,31,75,31,246,31,175,31,46,31,60,31,47,31,199,31,199,30,146,31,42,31,201,31,235,31,235,30,142,31,142,30,98,31,137,31,162,31,108,31,209,31,8,31,231,31,51,31,51,30,139,31,104,31,10,31,141,31,102,31,235,31,96,31,122,31,122,30,132,31,126,31,135,31,133,31,214,31,145,31,167,31,109,31,39,31,58,31,180,31,180,31,191,31,122,31,246,31,15,31,151,31,94,31,248,31,248,30,123,31,123,30,127,31,236,31,125,31,125,30,234,31,234,30,143,31,143,30,188,31,188,30,162,31,162,30,23,31,23,30,56,31,250,31,92,31,55,31,121,31,82,31,25,31,55,31,55,30,232,31,232,30,67,31,20,31,107,31,67,31,131,31,185,31,1,31,50,31,178,31,151,31,151,30,2,31,64,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
