-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 975;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (168,0,0,0,0,0,16,0,248,0,56,0,195,0,221,0,74,0,74,0,156,0,41,0,145,0,0,0,103,0,0,0,137,0,4,0,5,0,47,0,175,0,158,0,135,0,0,0,0,0,24,0,64,0,161,0,183,0,229,0,181,0,229,0,0,0,177,0,90,0,0,0,0,0,55,0,53,0,0,0,182,0,254,0,0,0,122,0,107,0,162,0,216,0,113,0,229,0,124,0,101,0,85,0,175,0,34,0,15,0,23,0,82,0,157,0,149,0,0,0,121,0,0,0,159,0,181,0,0,0,0,0,172,0,0,0,113,0,88,0,54,0,52,0,44,0,0,0,93,0,189,0,236,0,96,0,140,0,181,0,137,0,0,0,184,0,113,0,30,0,108,0,42,0,226,0,128,0,77,0,175,0,156,0,0,0,226,0,244,0,251,0,252,0,193,0,192,0,239,0,27,0,230,0,238,0,170,0,0,0,8,0,55,0,138,0,0,0,56,0,61,0,231,0,135,0,41,0,87,0,103,0,238,0,170,0,230,0,42,0,51,0,0,0,0,0,211,0,157,0,121,0,248,0,104,0,131,0,136,0,44,0,108,0,47,0,19,0,0,0,51,0,0,0,132,0,18,0,54,0,0,0,170,0,23,0,23,0,0,0,2,0,62,0,212,0,158,0,132,0,118,0,54,0,207,0,0,0,200,0,65,0,0,0,253,0,217,0,93,0,199,0,147,0,149,0,191,0,213,0,192,0,19,0,93,0,227,0,142,0,0,0,45,0,0,0,133,0,143,0,234,0,249,0,0,0,0,0,0,0,10,0,214,0,249,0,87,0,0,0,52,0,52,0,234,0,183,0,100,0,104,0,91,0,207,0,99,0,19,0,123,0,156,0,164,0,159,0,237,0,76,0,110,0,224,0,242,0,185,0,236,0,65,0,168,0,214,0,189,0,253,0,143,0,15,0,25,0,231,0,205,0,94,0,115,0,174,0,14,0,0,0,211,0,0,0,250,0,52,0,218,0,49,0,217,0,242,0,48,0,37,0,0,0,16,0,147,0,107,0,66,0,8,0,122,0,91,0,233,0,0,0,69,0,28,0,168,0,136,0,151,0,134,0,156,0,185,0,170,0,168,0,255,0,212,0,232,0,208,0,73,0,62,0,157,0,38,0,148,0,0,0,238,0,44,0,209,0,156,0,0,0,230,0,89,0,0,0,24,0,0,0,0,0,61,0,63,0,60,0,209,0,243,0,14,0,43,0,68,0,11,0,58,0,193,0,160,0,11,0,24,0,132,0,175,0,125,0,199,0,101,0,0,0,0,0,136,0,125,0,138,0,80,0,37,0,216,0,28,0,14,0,208,0,61,0,0,0,36,0,239,0,0,0,184,0,0,0,80,0,0,0,22,0,194,0,178,0,217,0,79,0,30,0,154,0,158,0,57,0,241,0,137,0,210,0,91,0,158,0,2,0,94,0,29,0,181,0,224,0,0,0,67,0,114,0,166,0,65,0,75,0,74,0,253,0,77,0,88,0,114,0,181,0,23,0,0,0,0,0,28,0,0,0,197,0,191,0,244,0,72,0,0,0,69,0,25,0,0,0,255,0,179,0,73,0,121,0,146,0,250,0,198,0,121,0,100,0,223,0,0,0,0,0,119,0,0,0,235,0,148,0,63,0,0,0,175,0,180,0,102,0,0,0,87,0,189,0,24,0,239,0,58,0,217,0,0,0,183,0,131,0,57,0,29,0,31,0,82,0,138,0,42,0,0,0,4,0,0,0,150,0,178,0,20,0,192,0,30,0,0,0,215,0,85,0,111,0,220,0,231,0,101,0,241,0,159,0,199,0,189,0,54,0,187,0,85,0,0,0,100,0,46,0,56,0,159,0,125,0,0,0,27,0,0,0,123,0,126,0,0,0,102,0,74,0,0,0,0,0,120,0,176,0,125,0,130,0,253,0,226,0,106,0,187,0,0,0,208,0,49,0,15,0,0,0,110,0,93,0,174,0,87,0,152,0,203,0,83,0,0,0,0,0,149,0,0,0,0,0,13,0,0,0,182,0,113,0,168,0,119,0,0,0,149,0,115,0,67,0,126,0,103,0,0,0,0,0,0,0,227,0,0,0,54,0,153,0,39,0,173,0,49,0,19,0,0,0,101,0,176,0,44,0,136,0,91,0,0,0,198,0,14,0,150,0,0,0,136,0,0,0,0,0,87,0,231,0,133,0,65,0,132,0,24,0,83,0,175,0,87,0,59,0,0,0,128,0,93,0,0,0,150,0,168,0,0,0,0,0,62,0,60,0,22,0,91,0,0,0,222,0,0,0,82,0,193,0,239,0,0,0,217,0,161,0,55,0,235,0,106,0,157,0,46,0,201,0,209,0,154,0,154,0,182,0,66,0,87,0,0,0,0,0,100,0,0,0,0,0,217,0,74,0,1,0,156,0,46,0,0,0,199,0,90,0,145,0,186,0,106,0,75,0,48,0,0,0,13,0,21,0,0,0,162,0,0,0,0,0,0,0,68,0,205,0,89,0,220,0,122,0,26,0,179,0,229,0,237,0,218,0,223,0,0,0,35,0,91,0,67,0,84,0,175,0,245,0,61,0,0,0,130,0,241,0,155,0,0,0,65,0,220,0,243,0,51,0,0,0,27,0,0,0,203,0,3,0,215,0,204,0,222,0,105,0,224,0,216,0,248,0,237,0,25,0,72,0,9,0,99,0,201,0,0,0,116,0,9,0,157,0,204,0,111,0,174,0,212,0,0,0,0,0,0,0,65,0,116,0,0,0,67,0,213,0,172,0,149,0,144,0,51,0,45,0,233,0,204,0,198,0,11,0,106,0,19,0,100,0,0,0,0,0,0,0,148,0,217,0,165,0,27,0,206,0,208,0,164,0,0,0,55,0,204,0,157,0,0,0,164,0,171,0,189,0,234,0,231,0,237,0,121,0,0,0,0,0,114,0,214,0,0,0,130,0,0,0,0,0,179,0,92,0,32,0,143,0,81,0,0,0,56,0,116,0,155,0,0,0,60,0,176,0,6,0,165,0,209,0,46,0,202,0,229,0,79,0,16,0,147,0,10,0,31,0,244,0,0,0,103,0,211,0,0,0,111,0,7,0,116,0,239,0,44,0,165,0,202,0,199,0,28,0,203,0,34,0,0,0,155,0,26,0,227,0,0,0,31,0,146,0,175,0,197,0,186,0,113,0,0,0,175,0,0,0,234,0,108,0,113,0,0,0,130,0,227,0,57,0,72,0,174,0,217,0,0,0,175,0,65,0,19,0,168,0,126,0,191,0,93,0,8,0,243,0,104,0,87,0,38,0,130,0,147,0,136,0,236,0,196,0,138,0,143,0,218,0,13,0,84,0,58,0,116,0,187,0,150,0,130,0,60,0,247,0,0,0,44,0,164,0,109,0,252,0,238,0,123,0,71,0,188,0,189,0,207,0,227,0,4,0,232,0,102,0,0,0,234,0,92,0,214,0,220,0,59,0,19,0,113,0,207,0,0,0,128,0,225,0,85,0,0,0,25,0,0,0,67,0,202,0,21,0,37,0,0,0,56,0,55,0,251,0,89,0,0,0,0,0,98,0,0,0,88,0,87,0,25,0,201,0,235,0,131,0,179,0,184,0,4,0,191,0,61,0,238,0,0,0,0,0,222,0,99,0,84,0,0,0,82,0,142,0,118,0,0,0,83,0,224,0,100,0,0,0,217,0,242,0,36,0,204,0,0,0,22,0,145,0,0,0,0,0,135,0,61,0,20,0,241,0,66,0,112,0,92,0,11,0,196,0,254,0,244,0,176,0,167,0,169,0,0,0,219,0,21,0,51,0,171,0,169,0,0,0,144,0,50,0,88,0,181,0,133,0,33,0,20,0,81,0,218,0,0,0,130,0,94,0,0,0,164,0,0,0,159,0,0,0,186,0,0,0,0,0,0,0,104,0,241,0,231,0,156,0,105,0,183,0,165,0,184,0,34,0,0,0,12,0,184,0,200,0,0,0,131,0,109,0,76,0,123,0,0,0,112,0,0,0,0,0,107,0,22,0,0,0,114,0,46,0,178,0,202,0,136,0,105,0,0,0,160,0,0,0,7,0,216,0,144,0,0,0,15,0,65,0,85,0,235,0,183,0,188,0,58,0,72,0,94,0,0,0,107,0,0,0,233,0,91,0,221,0,0,0,0,0,91,0,62,0,174,0,54,0,0,0,60,0,24,0,0,0,254,0,63,0,0,0,0,0,96,0,253,0,199,0,233,0,37,0,78,0,208,0,98,0,142,0,240,0,91,0,104,0,148,0,169,0,39,0,94,0,0,0,74,0,0,0,15,0,185,0,239,0,172,0,139,0,0,0,90,0,72,0,3,0,53,0);
signal scenario_full  : scenario_type := (168,31,168,30,168,29,16,31,248,31,56,31,195,31,221,31,74,31,74,31,156,31,41,31,145,31,145,30,103,31,103,30,137,31,4,31,5,31,47,31,175,31,158,31,135,31,135,30,135,29,24,31,64,31,161,31,183,31,229,31,181,31,229,31,229,30,177,31,90,31,90,30,90,29,55,31,53,31,53,30,182,31,254,31,254,30,122,31,107,31,162,31,216,31,113,31,229,31,124,31,101,31,85,31,175,31,34,31,15,31,23,31,82,31,157,31,149,31,149,30,121,31,121,30,159,31,181,31,181,30,181,29,172,31,172,30,113,31,88,31,54,31,52,31,44,31,44,30,93,31,189,31,236,31,96,31,140,31,181,31,137,31,137,30,184,31,113,31,30,31,108,31,42,31,226,31,128,31,77,31,175,31,156,31,156,30,226,31,244,31,251,31,252,31,193,31,192,31,239,31,27,31,230,31,238,31,170,31,170,30,8,31,55,31,138,31,138,30,56,31,61,31,231,31,135,31,41,31,87,31,103,31,238,31,170,31,230,31,42,31,51,31,51,30,51,29,211,31,157,31,121,31,248,31,104,31,131,31,136,31,44,31,108,31,47,31,19,31,19,30,51,31,51,30,132,31,18,31,54,31,54,30,170,31,23,31,23,31,23,30,2,31,62,31,212,31,158,31,132,31,118,31,54,31,207,31,207,30,200,31,65,31,65,30,253,31,217,31,93,31,199,31,147,31,149,31,191,31,213,31,192,31,19,31,93,31,227,31,142,31,142,30,45,31,45,30,133,31,143,31,234,31,249,31,249,30,249,29,249,28,10,31,214,31,249,31,87,31,87,30,52,31,52,31,234,31,183,31,100,31,104,31,91,31,207,31,99,31,19,31,123,31,156,31,164,31,159,31,237,31,76,31,110,31,224,31,242,31,185,31,236,31,65,31,168,31,214,31,189,31,253,31,143,31,15,31,25,31,231,31,205,31,94,31,115,31,174,31,14,31,14,30,211,31,211,30,250,31,52,31,218,31,49,31,217,31,242,31,48,31,37,31,37,30,16,31,147,31,107,31,66,31,8,31,122,31,91,31,233,31,233,30,69,31,28,31,168,31,136,31,151,31,134,31,156,31,185,31,170,31,168,31,255,31,212,31,232,31,208,31,73,31,62,31,157,31,38,31,148,31,148,30,238,31,44,31,209,31,156,31,156,30,230,31,89,31,89,30,24,31,24,30,24,29,61,31,63,31,60,31,209,31,243,31,14,31,43,31,68,31,11,31,58,31,193,31,160,31,11,31,24,31,132,31,175,31,125,31,199,31,101,31,101,30,101,29,136,31,125,31,138,31,80,31,37,31,216,31,28,31,14,31,208,31,61,31,61,30,36,31,239,31,239,30,184,31,184,30,80,31,80,30,22,31,194,31,178,31,217,31,79,31,30,31,154,31,158,31,57,31,241,31,137,31,210,31,91,31,158,31,2,31,94,31,29,31,181,31,224,31,224,30,67,31,114,31,166,31,65,31,75,31,74,31,253,31,77,31,88,31,114,31,181,31,23,31,23,30,23,29,28,31,28,30,197,31,191,31,244,31,72,31,72,30,69,31,25,31,25,30,255,31,179,31,73,31,121,31,146,31,250,31,198,31,121,31,100,31,223,31,223,30,223,29,119,31,119,30,235,31,148,31,63,31,63,30,175,31,180,31,102,31,102,30,87,31,189,31,24,31,239,31,58,31,217,31,217,30,183,31,131,31,57,31,29,31,31,31,82,31,138,31,42,31,42,30,4,31,4,30,150,31,178,31,20,31,192,31,30,31,30,30,215,31,85,31,111,31,220,31,231,31,101,31,241,31,159,31,199,31,189,31,54,31,187,31,85,31,85,30,100,31,46,31,56,31,159,31,125,31,125,30,27,31,27,30,123,31,126,31,126,30,102,31,74,31,74,30,74,29,120,31,176,31,125,31,130,31,253,31,226,31,106,31,187,31,187,30,208,31,49,31,15,31,15,30,110,31,93,31,174,31,87,31,152,31,203,31,83,31,83,30,83,29,149,31,149,30,149,29,13,31,13,30,182,31,113,31,168,31,119,31,119,30,149,31,115,31,67,31,126,31,103,31,103,30,103,29,103,28,227,31,227,30,54,31,153,31,39,31,173,31,49,31,19,31,19,30,101,31,176,31,44,31,136,31,91,31,91,30,198,31,14,31,150,31,150,30,136,31,136,30,136,29,87,31,231,31,133,31,65,31,132,31,24,31,83,31,175,31,87,31,59,31,59,30,128,31,93,31,93,30,150,31,168,31,168,30,168,29,62,31,60,31,22,31,91,31,91,30,222,31,222,30,82,31,193,31,239,31,239,30,217,31,161,31,55,31,235,31,106,31,157,31,46,31,201,31,209,31,154,31,154,31,182,31,66,31,87,31,87,30,87,29,100,31,100,30,100,29,217,31,74,31,1,31,156,31,46,31,46,30,199,31,90,31,145,31,186,31,106,31,75,31,48,31,48,30,13,31,21,31,21,30,162,31,162,30,162,29,162,28,68,31,205,31,89,31,220,31,122,31,26,31,179,31,229,31,237,31,218,31,223,31,223,30,35,31,91,31,67,31,84,31,175,31,245,31,61,31,61,30,130,31,241,31,155,31,155,30,65,31,220,31,243,31,51,31,51,30,27,31,27,30,203,31,3,31,215,31,204,31,222,31,105,31,224,31,216,31,248,31,237,31,25,31,72,31,9,31,99,31,201,31,201,30,116,31,9,31,157,31,204,31,111,31,174,31,212,31,212,30,212,29,212,28,65,31,116,31,116,30,67,31,213,31,172,31,149,31,144,31,51,31,45,31,233,31,204,31,198,31,11,31,106,31,19,31,100,31,100,30,100,29,100,28,148,31,217,31,165,31,27,31,206,31,208,31,164,31,164,30,55,31,204,31,157,31,157,30,164,31,171,31,189,31,234,31,231,31,237,31,121,31,121,30,121,29,114,31,214,31,214,30,130,31,130,30,130,29,179,31,92,31,32,31,143,31,81,31,81,30,56,31,116,31,155,31,155,30,60,31,176,31,6,31,165,31,209,31,46,31,202,31,229,31,79,31,16,31,147,31,10,31,31,31,244,31,244,30,103,31,211,31,211,30,111,31,7,31,116,31,239,31,44,31,165,31,202,31,199,31,28,31,203,31,34,31,34,30,155,31,26,31,227,31,227,30,31,31,146,31,175,31,197,31,186,31,113,31,113,30,175,31,175,30,234,31,108,31,113,31,113,30,130,31,227,31,57,31,72,31,174,31,217,31,217,30,175,31,65,31,19,31,168,31,126,31,191,31,93,31,8,31,243,31,104,31,87,31,38,31,130,31,147,31,136,31,236,31,196,31,138,31,143,31,218,31,13,31,84,31,58,31,116,31,187,31,150,31,130,31,60,31,247,31,247,30,44,31,164,31,109,31,252,31,238,31,123,31,71,31,188,31,189,31,207,31,227,31,4,31,232,31,102,31,102,30,234,31,92,31,214,31,220,31,59,31,19,31,113,31,207,31,207,30,128,31,225,31,85,31,85,30,25,31,25,30,67,31,202,31,21,31,37,31,37,30,56,31,55,31,251,31,89,31,89,30,89,29,98,31,98,30,88,31,87,31,25,31,201,31,235,31,131,31,179,31,184,31,4,31,191,31,61,31,238,31,238,30,238,29,222,31,99,31,84,31,84,30,82,31,142,31,118,31,118,30,83,31,224,31,100,31,100,30,217,31,242,31,36,31,204,31,204,30,22,31,145,31,145,30,145,29,135,31,61,31,20,31,241,31,66,31,112,31,92,31,11,31,196,31,254,31,244,31,176,31,167,31,169,31,169,30,219,31,21,31,51,31,171,31,169,31,169,30,144,31,50,31,88,31,181,31,133,31,33,31,20,31,81,31,218,31,218,30,130,31,94,31,94,30,164,31,164,30,159,31,159,30,186,31,186,30,186,29,186,28,104,31,241,31,231,31,156,31,105,31,183,31,165,31,184,31,34,31,34,30,12,31,184,31,200,31,200,30,131,31,109,31,76,31,123,31,123,30,112,31,112,30,112,29,107,31,22,31,22,30,114,31,46,31,178,31,202,31,136,31,105,31,105,30,160,31,160,30,7,31,216,31,144,31,144,30,15,31,65,31,85,31,235,31,183,31,188,31,58,31,72,31,94,31,94,30,107,31,107,30,233,31,91,31,221,31,221,30,221,29,91,31,62,31,174,31,54,31,54,30,60,31,24,31,24,30,254,31,63,31,63,30,63,29,96,31,253,31,199,31,233,31,37,31,78,31,208,31,98,31,142,31,240,31,91,31,104,31,148,31,169,31,39,31,94,31,94,30,74,31,74,30,15,31,185,31,239,31,172,31,139,31,139,30,90,31,72,31,3,31,53,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
