-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 647;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (125,0,0,0,142,0,0,0,0,0,15,0,211,0,125,0,93,0,244,0,237,0,181,0,13,0,0,0,156,0,0,0,28,0,186,0,140,0,138,0,115,0,78,0,235,0,67,0,0,0,0,0,25,0,0,0,130,0,140,0,168,0,39,0,62,0,185,0,200,0,35,0,68,0,169,0,9,0,13,0,190,0,47,0,126,0,144,0,152,0,146,0,0,0,223,0,165,0,0,0,157,0,0,0,224,0,14,0,142,0,0,0,0,0,12,0,213,0,79,0,0,0,225,0,140,0,186,0,56,0,0,0,90,0,222,0,88,0,161,0,149,0,116,0,0,0,235,0,210,0,117,0,0,0,187,0,130,0,240,0,48,0,0,0,119,0,181,0,0,0,5,0,19,0,181,0,0,0,9,0,0,0,108,0,41,0,49,0,0,0,80,0,127,0,7,0,0,0,219,0,158,0,0,0,53,0,192,0,240,0,0,0,244,0,174,0,81,0,0,0,127,0,4,0,122,0,32,0,224,0,88,0,0,0,103,0,174,0,78,0,99,0,31,0,72,0,255,0,24,0,197,0,53,0,63,0,0,0,99,0,118,0,0,0,96,0,0,0,253,0,32,0,228,0,195,0,29,0,191,0,197,0,10,0,243,0,228,0,143,0,0,0,206,0,0,0,0,0,248,0,0,0,188,0,0,0,123,0,36,0,0,0,71,0,2,0,0,0,126,0,0,0,18,0,255,0,2,0,0,0,88,0,74,0,0,0,0,0,5,0,192,0,55,0,0,0,197,0,226,0,0,0,177,0,129,0,12,0,239,0,53,0,51,0,200,0,161,0,198,0,84,0,213,0,18,0,95,0,226,0,0,0,41,0,189,0,0,0,117,0,51,0,0,0,7,0,0,0,143,0,56,0,52,0,0,0,211,0,36,0,146,0,216,0,189,0,0,0,243,0,0,0,0,0,116,0,0,0,156,0,196,0,167,0,0,0,0,0,251,0,6,0,233,0,198,0,117,0,240,0,199,0,143,0,244,0,178,0,124,0,186,0,140,0,206,0,49,0,102,0,200,0,154,0,0,0,174,0,225,0,240,0,154,0,0,0,214,0,0,0,101,0,0,0,149,0,72,0,0,0,134,0,45,0,236,0,41,0,118,0,193,0,0,0,90,0,151,0,245,0,186,0,91,0,79,0,20,0,96,0,0,0,0,0,0,0,151,0,0,0,83,0,99,0,0,0,255,0,0,0,186,0,154,0,0,0,38,0,248,0,0,0,0,0,225,0,196,0,184,0,71,0,234,0,27,0,36,0,78,0,68,0,39,0,0,0,92,0,28,0,137,0,61,0,197,0,8,0,0,0,113,0,0,0,180,0,61,0,86,0,55,0,57,0,163,0,196,0,0,0,140,0,87,0,94,0,212,0,242,0,169,0,0,0,207,0,21,0,0,0,38,0,209,0,0,0,0,0,125,0,86,0,195,0,127,0,0,0,251,0,0,0,0,0,234,0,0,0,78,0,0,0,171,0,117,0,205,0,0,0,70,0,0,0,178,0,100,0,0,0,90,0,0,0,143,0,150,0,180,0,80,0,80,0,0,0,0,0,181,0,68,0,238,0,58,0,58,0,203,0,153,0,0,0,216,0,220,0,143,0,0,0,125,0,188,0,100,0,0,0,0,0,35,0,30,0,74,0,0,0,127,0,89,0,242,0,204,0,113,0,152,0,238,0,236,0,136,0,231,0,60,0,111,0,158,0,9,0,0,0,137,0,0,0,0,0,197,0,0,0,0,0,135,0,180,0,12,0,0,0,177,0,63,0,192,0,0,0,235,0,0,0,36,0,250,0,165,0,11,0,0,0,0,0,227,0,144,0,96,0,171,0,189,0,51,0,0,0,245,0,182,0,70,0,181,0,109,0,101,0,32,0,153,0,190,0,128,0,77,0,0,0,224,0,39,0,230,0,197,0,253,0,251,0,0,0,254,0,54,0,11,0,102,0,26,0,115,0,254,0,33,0,232,0,50,0,58,0,0,0,0,0,0,0,3,0,46,0,122,0,0,0,128,0,4,0,139,0,74,0,208,0,125,0,0,0,131,0,70,0,160,0,192,0,0,0,197,0,229,0,244,0,68,0,42,0,229,0,148,0,0,0,5,0,33,0,71,0,0,0,0,0,170,0,59,0,0,0,215,0,14,0,229,0,69,0,8,0,127,0,0,0,160,0,108,0,211,0,184,0,6,0,193,0,207,0,1,0,19,0,0,0,121,0,82,0,124,0,205,0,210,0,45,0,132,0,83,0,157,0,184,0,54,0,147,0,43,0,251,0,0,0,47,0,35,0,181,0,155,0,86,0,0,0,60,0,5,0,136,0,0,0,191,0,96,0,125,0,149,0,101,0,21,0,81,0,160,0,169,0,0,0,173,0,95,0,52,0,189,0,23,0,106,0,10,0,96,0,84,0,0,0,213,0,76,0,186,0,39,0,30,0,85,0,39,0,78,0,208,0,0,0,251,0,51,0,13,0,56,0,140,0,234,0,115,0,70,0,209,0,0,0,206,0,16,0,166,0,164,0,0,0,25,0,178,0,226,0,41,0,197,0,107,0,204,0,0,0,136,0,214,0,71,0,167,0,17,0,0,0,164,0,21,0,0,0,0,0,246,0,69,0,0,0,0,0,67,0,50,0,116,0,86,0,156,0,0,0,0,0,0,0,241,0,91,0,35,0,70,0,0,0,71,0,74,0,46,0,215,0,58,0,23,0,159,0,118,0,130,0,0,0,140,0,131,0,0,0,156,0,119,0,8,0,86,0,161,0,252,0,24,0,0,0,160,0,97,0,250,0,46,0,78,0,121,0,51,0,156,0,28,0,38,0,7,0,68,0,0,0,182,0,0,0,158,0,15,0,165,0,102,0,108,0);
signal scenario_full  : scenario_type := (125,31,125,30,142,31,142,30,142,29,15,31,211,31,125,31,93,31,244,31,237,31,181,31,13,31,13,30,156,31,156,30,28,31,186,31,140,31,138,31,115,31,78,31,235,31,67,31,67,30,67,29,25,31,25,30,130,31,140,31,168,31,39,31,62,31,185,31,200,31,35,31,68,31,169,31,9,31,13,31,190,31,47,31,126,31,144,31,152,31,146,31,146,30,223,31,165,31,165,30,157,31,157,30,224,31,14,31,142,31,142,30,142,29,12,31,213,31,79,31,79,30,225,31,140,31,186,31,56,31,56,30,90,31,222,31,88,31,161,31,149,31,116,31,116,30,235,31,210,31,117,31,117,30,187,31,130,31,240,31,48,31,48,30,119,31,181,31,181,30,5,31,19,31,181,31,181,30,9,31,9,30,108,31,41,31,49,31,49,30,80,31,127,31,7,31,7,30,219,31,158,31,158,30,53,31,192,31,240,31,240,30,244,31,174,31,81,31,81,30,127,31,4,31,122,31,32,31,224,31,88,31,88,30,103,31,174,31,78,31,99,31,31,31,72,31,255,31,24,31,197,31,53,31,63,31,63,30,99,31,118,31,118,30,96,31,96,30,253,31,32,31,228,31,195,31,29,31,191,31,197,31,10,31,243,31,228,31,143,31,143,30,206,31,206,30,206,29,248,31,248,30,188,31,188,30,123,31,36,31,36,30,71,31,2,31,2,30,126,31,126,30,18,31,255,31,2,31,2,30,88,31,74,31,74,30,74,29,5,31,192,31,55,31,55,30,197,31,226,31,226,30,177,31,129,31,12,31,239,31,53,31,51,31,200,31,161,31,198,31,84,31,213,31,18,31,95,31,226,31,226,30,41,31,189,31,189,30,117,31,51,31,51,30,7,31,7,30,143,31,56,31,52,31,52,30,211,31,36,31,146,31,216,31,189,31,189,30,243,31,243,30,243,29,116,31,116,30,156,31,196,31,167,31,167,30,167,29,251,31,6,31,233,31,198,31,117,31,240,31,199,31,143,31,244,31,178,31,124,31,186,31,140,31,206,31,49,31,102,31,200,31,154,31,154,30,174,31,225,31,240,31,154,31,154,30,214,31,214,30,101,31,101,30,149,31,72,31,72,30,134,31,45,31,236,31,41,31,118,31,193,31,193,30,90,31,151,31,245,31,186,31,91,31,79,31,20,31,96,31,96,30,96,29,96,28,151,31,151,30,83,31,99,31,99,30,255,31,255,30,186,31,154,31,154,30,38,31,248,31,248,30,248,29,225,31,196,31,184,31,71,31,234,31,27,31,36,31,78,31,68,31,39,31,39,30,92,31,28,31,137,31,61,31,197,31,8,31,8,30,113,31,113,30,180,31,61,31,86,31,55,31,57,31,163,31,196,31,196,30,140,31,87,31,94,31,212,31,242,31,169,31,169,30,207,31,21,31,21,30,38,31,209,31,209,30,209,29,125,31,86,31,195,31,127,31,127,30,251,31,251,30,251,29,234,31,234,30,78,31,78,30,171,31,117,31,205,31,205,30,70,31,70,30,178,31,100,31,100,30,90,31,90,30,143,31,150,31,180,31,80,31,80,31,80,30,80,29,181,31,68,31,238,31,58,31,58,31,203,31,153,31,153,30,216,31,220,31,143,31,143,30,125,31,188,31,100,31,100,30,100,29,35,31,30,31,74,31,74,30,127,31,89,31,242,31,204,31,113,31,152,31,238,31,236,31,136,31,231,31,60,31,111,31,158,31,9,31,9,30,137,31,137,30,137,29,197,31,197,30,197,29,135,31,180,31,12,31,12,30,177,31,63,31,192,31,192,30,235,31,235,30,36,31,250,31,165,31,11,31,11,30,11,29,227,31,144,31,96,31,171,31,189,31,51,31,51,30,245,31,182,31,70,31,181,31,109,31,101,31,32,31,153,31,190,31,128,31,77,31,77,30,224,31,39,31,230,31,197,31,253,31,251,31,251,30,254,31,54,31,11,31,102,31,26,31,115,31,254,31,33,31,232,31,50,31,58,31,58,30,58,29,58,28,3,31,46,31,122,31,122,30,128,31,4,31,139,31,74,31,208,31,125,31,125,30,131,31,70,31,160,31,192,31,192,30,197,31,229,31,244,31,68,31,42,31,229,31,148,31,148,30,5,31,33,31,71,31,71,30,71,29,170,31,59,31,59,30,215,31,14,31,229,31,69,31,8,31,127,31,127,30,160,31,108,31,211,31,184,31,6,31,193,31,207,31,1,31,19,31,19,30,121,31,82,31,124,31,205,31,210,31,45,31,132,31,83,31,157,31,184,31,54,31,147,31,43,31,251,31,251,30,47,31,35,31,181,31,155,31,86,31,86,30,60,31,5,31,136,31,136,30,191,31,96,31,125,31,149,31,101,31,21,31,81,31,160,31,169,31,169,30,173,31,95,31,52,31,189,31,23,31,106,31,10,31,96,31,84,31,84,30,213,31,76,31,186,31,39,31,30,31,85,31,39,31,78,31,208,31,208,30,251,31,51,31,13,31,56,31,140,31,234,31,115,31,70,31,209,31,209,30,206,31,16,31,166,31,164,31,164,30,25,31,178,31,226,31,41,31,197,31,107,31,204,31,204,30,136,31,214,31,71,31,167,31,17,31,17,30,164,31,21,31,21,30,21,29,246,31,69,31,69,30,69,29,67,31,50,31,116,31,86,31,156,31,156,30,156,29,156,28,241,31,91,31,35,31,70,31,70,30,71,31,74,31,46,31,215,31,58,31,23,31,159,31,118,31,130,31,130,30,140,31,131,31,131,30,156,31,119,31,8,31,86,31,161,31,252,31,24,31,24,30,160,31,97,31,250,31,46,31,78,31,121,31,51,31,156,31,28,31,38,31,7,31,68,31,68,30,182,31,182,30,158,31,15,31,165,31,102,31,108,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
