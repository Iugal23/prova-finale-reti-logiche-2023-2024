-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_44 is
end project_tb_44;

architecture project_tb_arch_44 of project_tb_44 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1017;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (161,0,17,0,66,0,0,0,0,0,173,0,177,0,87,0,250,0,161,0,177,0,198,0,111,0,0,0,0,0,191,0,19,0,31,0,187,0,5,0,155,0,50,0,0,0,219,0,214,0,24,0,180,0,14,0,143,0,0,0,205,0,0,0,0,0,161,0,145,0,0,0,126,0,59,0,141,0,0,0,96,0,226,0,91,0,114,0,224,0,22,0,0,0,195,0,0,0,215,0,203,0,174,0,148,0,4,0,80,0,0,0,0,0,226,0,0,0,97,0,22,0,49,0,38,0,221,0,0,0,170,0,190,0,51,0,197,0,59,0,80,0,120,0,242,0,0,0,8,0,56,0,0,0,206,0,129,0,72,0,138,0,39,0,164,0,211,0,217,0,65,0,141,0,21,0,36,0,32,0,0,0,50,0,193,0,0,0,0,0,53,0,37,0,0,0,237,0,0,0,27,0,0,0,75,0,126,0,113,0,0,0,249,0,111,0,0,0,0,0,0,0,77,0,248,0,131,0,14,0,227,0,0,0,204,0,220,0,0,0,176,0,64,0,199,0,72,0,250,0,11,0,0,0,32,0,14,0,0,0,192,0,0,0,104,0,0,0,204,0,0,0,24,0,191,0,25,0,181,0,242,0,205,0,0,0,229,0,156,0,250,0,220,0,216,0,39,0,0,0,144,0,31,0,11,0,29,0,0,0,0,0,0,0,154,0,183,0,239,0,247,0,110,0,89,0,241,0,124,0,134,0,77,0,142,0,149,0,88,0,84,0,34,0,163,0,213,0,0,0,0,0,0,0,189,0,216,0,99,0,247,0,122,0,76,0,237,0,249,0,0,0,63,0,254,0,191,0,123,0,24,0,30,0,120,0,130,0,65,0,0,0,54,0,0,0,0,0,78,0,0,0,26,0,0,0,203,0,0,0,163,0,117,0,215,0,43,0,176,0,70,0,217,0,0,0,131,0,228,0,0,0,212,0,53,0,7,0,0,0,107,0,29,0,138,0,127,0,0,0,0,0,240,0,62,0,0,0,2,0,212,0,0,0,0,0,31,0,111,0,168,0,173,0,218,0,72,0,19,0,89,0,0,0,171,0,150,0,11,0,133,0,233,0,172,0,168,0,159,0,160,0,20,0,156,0,3,0,0,0,0,0,0,0,148,0,123,0,75,0,164,0,156,0,0,0,55,0,108,0,176,0,137,0,245,0,0,0,155,0,0,0,230,0,46,0,0,0,210,0,162,0,69,0,120,0,0,0,21,0,173,0,0,0,19,0,109,0,0,0,170,0,169,0,2,0,103,0,0,0,0,0,180,0,170,0,12,0,94,0,84,0,138,0,145,0,0,0,100,0,0,0,0,0,70,0,209,0,0,0,185,0,135,0,0,0,111,0,132,0,226,0,87,0,98,0,149,0,64,0,74,0,0,0,235,0,0,0,0,0,225,0,35,0,30,0,243,0,0,0,133,0,151,0,65,0,188,0,142,0,9,0,101,0,101,0,118,0,245,0,170,0,64,0,93,0,68,0,0,0,8,0,50,0,0,0,111,0,134,0,99,0,132,0,48,0,180,0,0,0,219,0,117,0,194,0,113,0,159,0,154,0,230,0,31,0,0,0,44,0,109,0,0,0,76,0,0,0,13,0,157,0,63,0,51,0,0,0,166,0,255,0,0,0,163,0,52,0,241,0,49,0,7,0,187,0,108,0,61,0,0,0,0,0,31,0,185,0,78,0,213,0,128,0,10,0,124,0,154,0,194,0,0,0,0,0,85,0,243,0,86,0,251,0,239,0,21,0,157,0,182,0,248,0,54,0,49,0,94,0,8,0,189,0,123,0,248,0,37,0,63,0,0,0,235,0,0,0,18,0,0,0,29,0,246,0,0,0,165,0,35,0,70,0,131,0,86,0,51,0,150,0,87,0,37,0,104,0,156,0,199,0,0,0,121,0,0,0,196,0,64,0,0,0,41,0,137,0,0,0,177,0,183,0,125,0,171,0,193,0,45,0,16,0,89,0,98,0,0,0,145,0,145,0,86,0,99,0,121,0,251,0,70,0,123,0,1,0,0,0,0,0,181,0,174,0,0,0,183,0,0,0,64,0,167,0,38,0,0,0,203,0,66,0,162,0,123,0,47,0,121,0,64,0,0,0,0,0,0,0,254,0,15,0,209,0,0,0,156,0,187,0,235,0,0,0,130,0,134,0,170,0,0,0,195,0,0,0,155,0,0,0,0,0,239,0,0,0,114,0,110,0,240,0,0,0,100,0,228,0,132,0,237,0,212,0,0,0,0,0,0,0,35,0,188,0,240,0,4,0,160,0,241,0,132,0,0,0,112,0,0,0,215,0,13,0,0,0,0,0,114,0,165,0,222,0,254,0,217,0,24,0,7,0,206,0,130,0,56,0,102,0,105,0,0,0,193,0,0,0,213,0,13,0,10,0,233,0,62,0,121,0,95,0,156,0,130,0,159,0,22,0,15,0,58,0,51,0,79,0,0,0,40,0,108,0,110,0,251,0,0,0,221,0,35,0,0,0,164,0,0,0,0,0,0,0,217,0,121,0,48,0,31,0,182,0,49,0,189,0,22,0,30,0,0,0,11,0,167,0,249,0,95,0,44,0,184,0,88,0,7,0,0,0,163,0,140,0,0,0,116,0,220,0,210,0,155,0,34,0,160,0,53,0,98,0,11,0,28,0,114,0,16,0,249,0,180,0,8,0,81,0,127,0,245,0,5,0,34,0,61,0,75,0,41,0,179,0,40,0,146,0,71,0,66,0,31,0,0,0,110,0,1,0,66,0,227,0,164,0,250,0,0,0,9,0,193,0,54,0,16,0,41,0,166,0,117,0,152,0,0,0,55,0,112,0,160,0,53,0,227,0,29,0,95,0,80,0,253,0,79,0,216,0,0,0,232,0,227,0,0,0,220,0,0,0,0,0,0,0,67,0,141,0,154,0,130,0,142,0,16,0,52,0,185,0,106,0,139,0,140,0,0,0,35,0,103,0,184,0,90,0,123,0,0,0,80,0,44,0,116,0,14,0,156,0,208,0,210,0,0,0,0,0,0,0,134,0,74,0,228,0,161,0,210,0,16,0,0,0,238,0,0,0,0,0,202,0,81,0,173,0,55,0,209,0,185,0,48,0,234,0,16,0,145,0,169,0,0,0,0,0,0,0,183,0,99,0,145,0,129,0,0,0,157,0,77,0,104,0,182,0,111,0,163,0,68,0,137,0,0,0,229,0,14,0,105,0,0,0,178,0,51,0,133,0,0,0,130,0,6,0,103,0,0,0,80,0,143,0,211,0,157,0,151,0,114,0,138,0,0,0,235,0,21,0,0,0,95,0,53,0,145,0,141,0,173,0,0,0,110,0,210,0,178,0,58,0,38,0,121,0,0,0,0,0,223,0,61,0,34,0,167,0,174,0,80,0,52,0,211,0,33,0,206,0,0,0,66,0,113,0,176,0,172,0,240,0,95,0,0,0,117,0,0,0,63,0,247,0,40,0,191,0,0,0,113,0,251,0,41,0,3,0,131,0,0,0,219,0,150,0,0,0,0,0,207,0,128,0,178,0,53,0,0,0,194,0,0,0,149,0,92,0,149,0,224,0,0,0,226,0,117,0,251,0,0,0,159,0,218,0,55,0,91,0,97,0,0,0,224,0,250,0,208,0,41,0,208,0,128,0,220,0,132,0,171,0,0,0,27,0,206,0,23,0,60,0,0,0,0,0,229,0,193,0,246,0,253,0,238,0,198,0,240,0,0,0,0,0,0,0,147,0,214,0,247,0,253,0,0,0,0,0,127,0,34,0,191,0,0,0,85,0,239,0,39,0,0,0,189,0,163,0,70,0,131,0,0,0,26,0,162,0,46,0,39,0,247,0,0,0,215,0,122,0,110,0,175,0,53,0,185,0,0,0,233,0,112,0,224,0,111,0,210,0,0,0,95,0,180,0,105,0,0,0,219,0,0,0,150,0,109,0,195,0,0,0,0,0,0,0,113,0,205,0,0,0,163,0,19,0,246,0,138,0,161,0,148,0,0,0,123,0,214,0,85,0,24,0,54,0,82,0,67,0,62,0,160,0,137,0,83,0,245,0,0,0,138,0,17,0,187,0,119,0,160,0,210,0,73,0,105,0,84,0,83,0,0,0,35,0,20,0,220,0,114,0,185,0,39,0,233,0,200,0,0,0,83,0,19,0,65,0,235,0,191,0,0,0,42,0,222,0,148,0,41,0,135,0,0,0,165,0,0,0,200,0,0,0,78,0,231,0,220,0,0,0,174,0,0,0,69,0,206,0,46,0,67,0,0,0,174,0,10,0,0,0,204,0,245,0,23,0,84,0,98,0,9,0,71,0,236,0,197,0,67,0,191,0,70,0,208,0,0,0,219,0,104,0,74,0,72,0,185,0,114,0,36,0,151,0,0,0,185,0,237,0,17,0,132,0,112,0,222,0,23,0,0,0,124,0,134,0,0,0,9,0,242,0,237,0,221,0,236,0,0,0,21,0,44,0,0,0,215,0,54,0,42,0,0,0,31,0,92,0,0,0,254,0,0,0,215,0);
signal scenario_full  : scenario_type := (161,31,17,31,66,31,66,30,66,29,173,31,177,31,87,31,250,31,161,31,177,31,198,31,111,31,111,30,111,29,191,31,19,31,31,31,187,31,5,31,155,31,50,31,50,30,219,31,214,31,24,31,180,31,14,31,143,31,143,30,205,31,205,30,205,29,161,31,145,31,145,30,126,31,59,31,141,31,141,30,96,31,226,31,91,31,114,31,224,31,22,31,22,30,195,31,195,30,215,31,203,31,174,31,148,31,4,31,80,31,80,30,80,29,226,31,226,30,97,31,22,31,49,31,38,31,221,31,221,30,170,31,190,31,51,31,197,31,59,31,80,31,120,31,242,31,242,30,8,31,56,31,56,30,206,31,129,31,72,31,138,31,39,31,164,31,211,31,217,31,65,31,141,31,21,31,36,31,32,31,32,30,50,31,193,31,193,30,193,29,53,31,37,31,37,30,237,31,237,30,27,31,27,30,75,31,126,31,113,31,113,30,249,31,111,31,111,30,111,29,111,28,77,31,248,31,131,31,14,31,227,31,227,30,204,31,220,31,220,30,176,31,64,31,199,31,72,31,250,31,11,31,11,30,32,31,14,31,14,30,192,31,192,30,104,31,104,30,204,31,204,30,24,31,191,31,25,31,181,31,242,31,205,31,205,30,229,31,156,31,250,31,220,31,216,31,39,31,39,30,144,31,31,31,11,31,29,31,29,30,29,29,29,28,154,31,183,31,239,31,247,31,110,31,89,31,241,31,124,31,134,31,77,31,142,31,149,31,88,31,84,31,34,31,163,31,213,31,213,30,213,29,213,28,189,31,216,31,99,31,247,31,122,31,76,31,237,31,249,31,249,30,63,31,254,31,191,31,123,31,24,31,30,31,120,31,130,31,65,31,65,30,54,31,54,30,54,29,78,31,78,30,26,31,26,30,203,31,203,30,163,31,117,31,215,31,43,31,176,31,70,31,217,31,217,30,131,31,228,31,228,30,212,31,53,31,7,31,7,30,107,31,29,31,138,31,127,31,127,30,127,29,240,31,62,31,62,30,2,31,212,31,212,30,212,29,31,31,111,31,168,31,173,31,218,31,72,31,19,31,89,31,89,30,171,31,150,31,11,31,133,31,233,31,172,31,168,31,159,31,160,31,20,31,156,31,3,31,3,30,3,29,3,28,148,31,123,31,75,31,164,31,156,31,156,30,55,31,108,31,176,31,137,31,245,31,245,30,155,31,155,30,230,31,46,31,46,30,210,31,162,31,69,31,120,31,120,30,21,31,173,31,173,30,19,31,109,31,109,30,170,31,169,31,2,31,103,31,103,30,103,29,180,31,170,31,12,31,94,31,84,31,138,31,145,31,145,30,100,31,100,30,100,29,70,31,209,31,209,30,185,31,135,31,135,30,111,31,132,31,226,31,87,31,98,31,149,31,64,31,74,31,74,30,235,31,235,30,235,29,225,31,35,31,30,31,243,31,243,30,133,31,151,31,65,31,188,31,142,31,9,31,101,31,101,31,118,31,245,31,170,31,64,31,93,31,68,31,68,30,8,31,50,31,50,30,111,31,134,31,99,31,132,31,48,31,180,31,180,30,219,31,117,31,194,31,113,31,159,31,154,31,230,31,31,31,31,30,44,31,109,31,109,30,76,31,76,30,13,31,157,31,63,31,51,31,51,30,166,31,255,31,255,30,163,31,52,31,241,31,49,31,7,31,187,31,108,31,61,31,61,30,61,29,31,31,185,31,78,31,213,31,128,31,10,31,124,31,154,31,194,31,194,30,194,29,85,31,243,31,86,31,251,31,239,31,21,31,157,31,182,31,248,31,54,31,49,31,94,31,8,31,189,31,123,31,248,31,37,31,63,31,63,30,235,31,235,30,18,31,18,30,29,31,246,31,246,30,165,31,35,31,70,31,131,31,86,31,51,31,150,31,87,31,37,31,104,31,156,31,199,31,199,30,121,31,121,30,196,31,64,31,64,30,41,31,137,31,137,30,177,31,183,31,125,31,171,31,193,31,45,31,16,31,89,31,98,31,98,30,145,31,145,31,86,31,99,31,121,31,251,31,70,31,123,31,1,31,1,30,1,29,181,31,174,31,174,30,183,31,183,30,64,31,167,31,38,31,38,30,203,31,66,31,162,31,123,31,47,31,121,31,64,31,64,30,64,29,64,28,254,31,15,31,209,31,209,30,156,31,187,31,235,31,235,30,130,31,134,31,170,31,170,30,195,31,195,30,155,31,155,30,155,29,239,31,239,30,114,31,110,31,240,31,240,30,100,31,228,31,132,31,237,31,212,31,212,30,212,29,212,28,35,31,188,31,240,31,4,31,160,31,241,31,132,31,132,30,112,31,112,30,215,31,13,31,13,30,13,29,114,31,165,31,222,31,254,31,217,31,24,31,7,31,206,31,130,31,56,31,102,31,105,31,105,30,193,31,193,30,213,31,13,31,10,31,233,31,62,31,121,31,95,31,156,31,130,31,159,31,22,31,15,31,58,31,51,31,79,31,79,30,40,31,108,31,110,31,251,31,251,30,221,31,35,31,35,30,164,31,164,30,164,29,164,28,217,31,121,31,48,31,31,31,182,31,49,31,189,31,22,31,30,31,30,30,11,31,167,31,249,31,95,31,44,31,184,31,88,31,7,31,7,30,163,31,140,31,140,30,116,31,220,31,210,31,155,31,34,31,160,31,53,31,98,31,11,31,28,31,114,31,16,31,249,31,180,31,8,31,81,31,127,31,245,31,5,31,34,31,61,31,75,31,41,31,179,31,40,31,146,31,71,31,66,31,31,31,31,30,110,31,1,31,66,31,227,31,164,31,250,31,250,30,9,31,193,31,54,31,16,31,41,31,166,31,117,31,152,31,152,30,55,31,112,31,160,31,53,31,227,31,29,31,95,31,80,31,253,31,79,31,216,31,216,30,232,31,227,31,227,30,220,31,220,30,220,29,220,28,67,31,141,31,154,31,130,31,142,31,16,31,52,31,185,31,106,31,139,31,140,31,140,30,35,31,103,31,184,31,90,31,123,31,123,30,80,31,44,31,116,31,14,31,156,31,208,31,210,31,210,30,210,29,210,28,134,31,74,31,228,31,161,31,210,31,16,31,16,30,238,31,238,30,238,29,202,31,81,31,173,31,55,31,209,31,185,31,48,31,234,31,16,31,145,31,169,31,169,30,169,29,169,28,183,31,99,31,145,31,129,31,129,30,157,31,77,31,104,31,182,31,111,31,163,31,68,31,137,31,137,30,229,31,14,31,105,31,105,30,178,31,51,31,133,31,133,30,130,31,6,31,103,31,103,30,80,31,143,31,211,31,157,31,151,31,114,31,138,31,138,30,235,31,21,31,21,30,95,31,53,31,145,31,141,31,173,31,173,30,110,31,210,31,178,31,58,31,38,31,121,31,121,30,121,29,223,31,61,31,34,31,167,31,174,31,80,31,52,31,211,31,33,31,206,31,206,30,66,31,113,31,176,31,172,31,240,31,95,31,95,30,117,31,117,30,63,31,247,31,40,31,191,31,191,30,113,31,251,31,41,31,3,31,131,31,131,30,219,31,150,31,150,30,150,29,207,31,128,31,178,31,53,31,53,30,194,31,194,30,149,31,92,31,149,31,224,31,224,30,226,31,117,31,251,31,251,30,159,31,218,31,55,31,91,31,97,31,97,30,224,31,250,31,208,31,41,31,208,31,128,31,220,31,132,31,171,31,171,30,27,31,206,31,23,31,60,31,60,30,60,29,229,31,193,31,246,31,253,31,238,31,198,31,240,31,240,30,240,29,240,28,147,31,214,31,247,31,253,31,253,30,253,29,127,31,34,31,191,31,191,30,85,31,239,31,39,31,39,30,189,31,163,31,70,31,131,31,131,30,26,31,162,31,46,31,39,31,247,31,247,30,215,31,122,31,110,31,175,31,53,31,185,31,185,30,233,31,112,31,224,31,111,31,210,31,210,30,95,31,180,31,105,31,105,30,219,31,219,30,150,31,109,31,195,31,195,30,195,29,195,28,113,31,205,31,205,30,163,31,19,31,246,31,138,31,161,31,148,31,148,30,123,31,214,31,85,31,24,31,54,31,82,31,67,31,62,31,160,31,137,31,83,31,245,31,245,30,138,31,17,31,187,31,119,31,160,31,210,31,73,31,105,31,84,31,83,31,83,30,35,31,20,31,220,31,114,31,185,31,39,31,233,31,200,31,200,30,83,31,19,31,65,31,235,31,191,31,191,30,42,31,222,31,148,31,41,31,135,31,135,30,165,31,165,30,200,31,200,30,78,31,231,31,220,31,220,30,174,31,174,30,69,31,206,31,46,31,67,31,67,30,174,31,10,31,10,30,204,31,245,31,23,31,84,31,98,31,9,31,71,31,236,31,197,31,67,31,191,31,70,31,208,31,208,30,219,31,104,31,74,31,72,31,185,31,114,31,36,31,151,31,151,30,185,31,237,31,17,31,132,31,112,31,222,31,23,31,23,30,124,31,134,31,134,30,9,31,242,31,237,31,221,31,236,31,236,30,21,31,44,31,44,30,215,31,54,31,42,31,42,30,31,31,92,31,92,30,254,31,254,30,215,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
