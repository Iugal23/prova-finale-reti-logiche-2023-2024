-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 213;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,162,0,118,0,42,0,145,0,98,0,66,0,60,0,99,0,0,0,2,0,106,0,0,0,209,0,111,0,82,0,186,0,168,0,198,0,225,0,249,0,205,0,73,0,113,0,213,0,76,0,58,0,164,0,139,0,59,0,0,0,0,0,177,0,146,0,109,0,202,0,149,0,183,0,206,0,75,0,107,0,79,0,240,0,255,0,233,0,75,0,87,0,145,0,68,0,69,0,44,0,39,0,146,0,42,0,0,0,41,0,204,0,70,0,193,0,254,0,0,0,0,0,0,0,17,0,91,0,95,0,229,0,161,0,0,0,9,0,105,0,214,0,0,0,102,0,193,0,249,0,118,0,215,0,223,0,250,0,87,0,167,0,46,0,70,0,33,0,56,0,238,0,123,0,202,0,0,0,0,0,239,0,110,0,183,0,215,0,197,0,54,0,216,0,62,0,0,0,46,0,180,0,0,0,0,0,201,0,137,0,34,0,181,0,47,0,175,0,226,0,228,0,0,0,232,0,111,0,160,0,90,0,236,0,126,0,0,0,86,0,0,0,75,0,42,0,237,0,197,0,0,0,227,0,165,0,12,0,158,0,0,0,206,0,0,0,156,0,44,0,214,0,0,0,3,0,176,0,215,0,32,0,58,0,231,0,106,0,0,0,110,0,214,0,57,0,91,0,127,0,197,0,15,0,49,0,0,0,214,0,122,0,195,0,194,0,156,0,0,0,237,0,0,0,116,0,0,0,198,0,0,0,147,0,0,0,0,0,166,0,229,0,3,0,184,0,105,0,203,0,227,0,203,0,28,0,0,0,233,0,81,0,0,0,66,0,84,0,0,0,95,0,150,0,101,0,38,0,25,0,41,0,216,0,99,0,144,0,212,0,119,0,132,0,0,0,205,0,221,0,166,0,0,0,125,0,15,0,67,0,115,0,35,0,0,0,0,0,101,0,231,0,188,0);
signal scenario_full  : scenario_type := (0,0,162,31,118,31,42,31,145,31,98,31,66,31,60,31,99,31,99,30,2,31,106,31,106,30,209,31,111,31,82,31,186,31,168,31,198,31,225,31,249,31,205,31,73,31,113,31,213,31,76,31,58,31,164,31,139,31,59,31,59,30,59,29,177,31,146,31,109,31,202,31,149,31,183,31,206,31,75,31,107,31,79,31,240,31,255,31,233,31,75,31,87,31,145,31,68,31,69,31,44,31,39,31,146,31,42,31,42,30,41,31,204,31,70,31,193,31,254,31,254,30,254,29,254,28,17,31,91,31,95,31,229,31,161,31,161,30,9,31,105,31,214,31,214,30,102,31,193,31,249,31,118,31,215,31,223,31,250,31,87,31,167,31,46,31,70,31,33,31,56,31,238,31,123,31,202,31,202,30,202,29,239,31,110,31,183,31,215,31,197,31,54,31,216,31,62,31,62,30,46,31,180,31,180,30,180,29,201,31,137,31,34,31,181,31,47,31,175,31,226,31,228,31,228,30,232,31,111,31,160,31,90,31,236,31,126,31,126,30,86,31,86,30,75,31,42,31,237,31,197,31,197,30,227,31,165,31,12,31,158,31,158,30,206,31,206,30,156,31,44,31,214,31,214,30,3,31,176,31,215,31,32,31,58,31,231,31,106,31,106,30,110,31,214,31,57,31,91,31,127,31,197,31,15,31,49,31,49,30,214,31,122,31,195,31,194,31,156,31,156,30,237,31,237,30,116,31,116,30,198,31,198,30,147,31,147,30,147,29,166,31,229,31,3,31,184,31,105,31,203,31,227,31,203,31,28,31,28,30,233,31,81,31,81,30,66,31,84,31,84,30,95,31,150,31,101,31,38,31,25,31,41,31,216,31,99,31,144,31,212,31,119,31,132,31,132,30,205,31,221,31,166,31,166,30,125,31,15,31,67,31,115,31,35,31,35,30,35,29,101,31,231,31,188,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
