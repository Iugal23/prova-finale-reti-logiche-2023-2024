-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 523;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (107,0,0,0,63,0,122,0,0,0,189,0,9,0,0,0,0,0,0,0,210,0,109,0,0,0,0,0,57,0,22,0,0,0,147,0,0,0,154,0,85,0,130,0,166,0,0,0,83,0,0,0,192,0,9,0,175,0,55,0,217,0,63,0,0,0,219,0,223,0,0,0,186,0,0,0,174,0,184,0,84,0,108,0,229,0,180,0,191,0,202,0,0,0,0,0,164,0,0,0,249,0,0,0,35,0,183,0,121,0,0,0,0,0,203,0,4,0,98,0,62,0,153,0,0,0,185,0,167,0,153,0,3,0,62,0,19,0,13,0,94,0,137,0,181,0,149,0,127,0,234,0,32,0,0,0,46,0,0,0,47,0,208,0,143,0,173,0,0,0,174,0,27,0,141,0,50,0,0,0,162,0,96,0,12,0,195,0,0,0,199,0,101,0,102,0,82,0,202,0,95,0,44,0,155,0,178,0,162,0,110,0,157,0,247,0,140,0,0,0,134,0,155,0,191,0,39,0,142,0,139,0,201,0,24,0,123,0,203,0,231,0,80,0,58,0,242,0,157,0,43,0,217,0,160,0,135,0,53,0,183,0,0,0,24,0,247,0,62,0,234,0,43,0,105,0,0,0,232,0,0,0,32,0,134,0,15,0,211,0,181,0,0,0,44,0,11,0,214,0,36,0,61,0,113,0,204,0,0,0,25,0,244,0,178,0,239,0,4,0,0,0,239,0,0,0,253,0,23,0,41,0,0,0,245,0,78,0,41,0,0,0,239,0,0,0,44,0,39,0,66,0,47,0,187,0,234,0,85,0,0,0,117,0,19,0,94,0,228,0,50,0,91,0,0,0,129,0,7,0,180,0,213,0,0,0,73,0,23,0,63,0,125,0,44,0,0,0,2,0,236,0,114,0,3,0,142,0,108,0,1,0,43,0,130,0,0,0,183,0,139,0,8,0,51,0,167,0,5,0,36,0,85,0,0,0,235,0,171,0,22,0,0,0,2,0,189,0,85,0,245,0,83,0,217,0,97,0,0,0,13,0,167,0,168,0,244,0,150,0,196,0,165,0,192,0,81,0,0,0,109,0,190,0,0,0,41,0,214,0,191,0,194,0,150,0,246,0,0,0,121,0,211,0,74,0,95,0,154,0,147,0,250,0,83,0,34,0,254,0,162,0,188,0,146,0,231,0,0,0,36,0,52,0,151,0,28,0,221,0,155,0,78,0,149,0,0,0,38,0,0,0,100,0,176,0,0,0,78,0,0,0,35,0,243,0,237,0,0,0,162,0,177,0,224,0,168,0,78,0,0,0,86,0,13,0,0,0,182,0,41,0,97,0,145,0,162,0,120,0,227,0,142,0,160,0,139,0,204,0,185,0,0,0,77,0,29,0,111,0,0,0,0,0,1,0,100,0,229,0,48,0,0,0,18,0,0,0,158,0,50,0,82,0,36,0,0,0,0,0,0,0,0,0,140,0,202,0,218,0,76,0,213,0,248,0,147,0,11,0,88,0,68,0,114,0,221,0,103,0,161,0,206,0,66,0,0,0,58,0,206,0,0,0,116,0,127,0,0,0,38,0,145,0,100,0,237,0,95,0,152,0,101,0,0,0,130,0,0,0,0,0,222,0,154,0,248,0,208,0,230,0,92,0,129,0,194,0,0,0,46,0,5,0,44,0,0,0,136,0,233,0,120,0,242,0,134,0,0,0,156,0,0,0,101,0,219,0,89,0,154,0,87,0,173,0,113,0,31,0,186,0,152,0,222,0,62,0,251,0,189,0,0,0,0,0,0,0,0,0,91,0,0,0,168,0,250,0,18,0,77,0,3,0,10,0,3,0,239,0,0,0,42,0,101,0,0,0,0,0,73,0,134,0,126,0,148,0,168,0,36,0,222,0,222,0,24,0,252,0,80,0,231,0,106,0,183,0,190,0,255,0,69,0,20,0,111,0,107,0,0,0,103,0,46,0,122,0,168,0,155,0,0,0,0,0,240,0,148,0,247,0,0,0,197,0,156,0,108,0,243,0,115,0,0,0,192,0,130,0,252,0,0,0,53,0,0,0,64,0,0,0,60,0,216,0,0,0,239,0,108,0,0,0,180,0,0,0,0,0,115,0,237,0,11,0,218,0,88,0,0,0,0,0,112,0,64,0,23,0,114,0,0,0,178,0,24,0,0,0,62,0,0,0,245,0,10,0,0,0,99,0,0,0,26,0,234,0,237,0,84,0,38,0,0,0,186,0,78,0,16,0,10,0,207,0,23,0,185,0,122,0,156,0,241,0,39,0,169,0,221,0,75,0,0,0,70,0,104,0,230,0,0,0,124,0,242,0,65,0,55,0,66,0,144,0);
signal scenario_full  : scenario_type := (107,31,107,30,63,31,122,31,122,30,189,31,9,31,9,30,9,29,9,28,210,31,109,31,109,30,109,29,57,31,22,31,22,30,147,31,147,30,154,31,85,31,130,31,166,31,166,30,83,31,83,30,192,31,9,31,175,31,55,31,217,31,63,31,63,30,219,31,223,31,223,30,186,31,186,30,174,31,184,31,84,31,108,31,229,31,180,31,191,31,202,31,202,30,202,29,164,31,164,30,249,31,249,30,35,31,183,31,121,31,121,30,121,29,203,31,4,31,98,31,62,31,153,31,153,30,185,31,167,31,153,31,3,31,62,31,19,31,13,31,94,31,137,31,181,31,149,31,127,31,234,31,32,31,32,30,46,31,46,30,47,31,208,31,143,31,173,31,173,30,174,31,27,31,141,31,50,31,50,30,162,31,96,31,12,31,195,31,195,30,199,31,101,31,102,31,82,31,202,31,95,31,44,31,155,31,178,31,162,31,110,31,157,31,247,31,140,31,140,30,134,31,155,31,191,31,39,31,142,31,139,31,201,31,24,31,123,31,203,31,231,31,80,31,58,31,242,31,157,31,43,31,217,31,160,31,135,31,53,31,183,31,183,30,24,31,247,31,62,31,234,31,43,31,105,31,105,30,232,31,232,30,32,31,134,31,15,31,211,31,181,31,181,30,44,31,11,31,214,31,36,31,61,31,113,31,204,31,204,30,25,31,244,31,178,31,239,31,4,31,4,30,239,31,239,30,253,31,23,31,41,31,41,30,245,31,78,31,41,31,41,30,239,31,239,30,44,31,39,31,66,31,47,31,187,31,234,31,85,31,85,30,117,31,19,31,94,31,228,31,50,31,91,31,91,30,129,31,7,31,180,31,213,31,213,30,73,31,23,31,63,31,125,31,44,31,44,30,2,31,236,31,114,31,3,31,142,31,108,31,1,31,43,31,130,31,130,30,183,31,139,31,8,31,51,31,167,31,5,31,36,31,85,31,85,30,235,31,171,31,22,31,22,30,2,31,189,31,85,31,245,31,83,31,217,31,97,31,97,30,13,31,167,31,168,31,244,31,150,31,196,31,165,31,192,31,81,31,81,30,109,31,190,31,190,30,41,31,214,31,191,31,194,31,150,31,246,31,246,30,121,31,211,31,74,31,95,31,154,31,147,31,250,31,83,31,34,31,254,31,162,31,188,31,146,31,231,31,231,30,36,31,52,31,151,31,28,31,221,31,155,31,78,31,149,31,149,30,38,31,38,30,100,31,176,31,176,30,78,31,78,30,35,31,243,31,237,31,237,30,162,31,177,31,224,31,168,31,78,31,78,30,86,31,13,31,13,30,182,31,41,31,97,31,145,31,162,31,120,31,227,31,142,31,160,31,139,31,204,31,185,31,185,30,77,31,29,31,111,31,111,30,111,29,1,31,100,31,229,31,48,31,48,30,18,31,18,30,158,31,50,31,82,31,36,31,36,30,36,29,36,28,36,27,140,31,202,31,218,31,76,31,213,31,248,31,147,31,11,31,88,31,68,31,114,31,221,31,103,31,161,31,206,31,66,31,66,30,58,31,206,31,206,30,116,31,127,31,127,30,38,31,145,31,100,31,237,31,95,31,152,31,101,31,101,30,130,31,130,30,130,29,222,31,154,31,248,31,208,31,230,31,92,31,129,31,194,31,194,30,46,31,5,31,44,31,44,30,136,31,233,31,120,31,242,31,134,31,134,30,156,31,156,30,101,31,219,31,89,31,154,31,87,31,173,31,113,31,31,31,186,31,152,31,222,31,62,31,251,31,189,31,189,30,189,29,189,28,189,27,91,31,91,30,168,31,250,31,18,31,77,31,3,31,10,31,3,31,239,31,239,30,42,31,101,31,101,30,101,29,73,31,134,31,126,31,148,31,168,31,36,31,222,31,222,31,24,31,252,31,80,31,231,31,106,31,183,31,190,31,255,31,69,31,20,31,111,31,107,31,107,30,103,31,46,31,122,31,168,31,155,31,155,30,155,29,240,31,148,31,247,31,247,30,197,31,156,31,108,31,243,31,115,31,115,30,192,31,130,31,252,31,252,30,53,31,53,30,64,31,64,30,60,31,216,31,216,30,239,31,108,31,108,30,180,31,180,30,180,29,115,31,237,31,11,31,218,31,88,31,88,30,88,29,112,31,64,31,23,31,114,31,114,30,178,31,24,31,24,30,62,31,62,30,245,31,10,31,10,30,99,31,99,30,26,31,234,31,237,31,84,31,38,31,38,30,186,31,78,31,16,31,10,31,207,31,23,31,185,31,122,31,156,31,241,31,39,31,169,31,221,31,75,31,75,30,70,31,104,31,230,31,230,30,124,31,242,31,65,31,55,31,66,31,144,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
