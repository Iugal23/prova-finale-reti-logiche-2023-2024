-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 504;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,40,0,136,0,0,0,132,0,241,0,62,0,249,0,0,0,0,0,111,0,57,0,227,0,0,0,231,0,216,0,231,0,82,0,0,0,105,0,236,0,2,0,150,0,16,0,30,0,0,0,8,0,60,0,119,0,185,0,64,0,179,0,87,0,0,0,0,0,0,0,224,0,142,0,175,0,0,0,171,0,106,0,24,0,186,0,0,0,141,0,86,0,120,0,227,0,158,0,221,0,218,0,0,0,43,0,0,0,191,0,27,0,0,0,23,0,117,0,238,0,0,0,217,0,227,0,59,0,75,0,0,0,6,0,87,0,0,0,208,0,0,0,47,0,66,0,189,0,114,0,244,0,27,0,100,0,23,0,94,0,214,0,0,0,69,0,225,0,198,0,248,0,189,0,133,0,0,0,122,0,39,0,179,0,0,0,51,0,0,0,251,0,186,0,42,0,207,0,155,0,32,0,0,0,209,0,207,0,0,0,204,0,178,0,115,0,103,0,16,0,0,0,239,0,11,0,206,0,246,0,121,0,0,0,0,0,15,0,139,0,130,0,222,0,0,0,70,0,53,0,42,0,98,0,131,0,223,0,0,0,30,0,48,0,74,0,220,0,0,0,239,0,57,0,0,0,98,0,12,0,23,0,45,0,170,0,130,0,0,0,199,0,154,0,0,0,197,0,209,0,163,0,162,0,0,0,146,0,136,0,252,0,54,0,0,0,0,0,144,0,57,0,10,0,161,0,219,0,173,0,28,0,60,0,187,0,96,0,221,0,0,0,12,0,87,0,40,0,109,0,210,0,208,0,192,0,0,0,23,0,36,0,218,0,150,0,173,0,113,0,34,0,94,0,63,0,142,0,164,0,0,0,170,0,6,0,93,0,134,0,135,0,159,0,87,0,54,0,131,0,241,0,0,0,82,0,200,0,100,0,98,0,136,0,179,0,6,0,198,0,0,0,151,0,25,0,36,0,110,0,171,0,245,0,0,0,0,0,203,0,178,0,67,0,0,0,0,0,100,0,243,0,125,0,254,0,20,0,210,0,234,0,23,0,0,0,82,0,183,0,21,0,232,0,0,0,19,0,144,0,255,0,22,0,10,0,204,0,65,0,87,0,156,0,217,0,155,0,163,0,0,0,59,0,91,0,145,0,84,0,0,0,0,0,70,0,218,0,0,0,168,0,0,0,118,0,58,0,114,0,114,0,194,0,27,0,217,0,38,0,16,0,65,0,0,0,168,0,52,0,0,0,224,0,152,0,83,0,20,0,158,0,79,0,4,0,147,0,192,0,0,0,170,0,0,0,160,0,115,0,187,0,69,0,238,0,122,0,199,0,0,0,68,0,149,0,47,0,56,0,155,0,181,0,42,0,228,0,0,0,91,0,148,0,187,0,211,0,0,0,0,0,84,0,246,0,0,0,125,0,68,0,203,0,102,0,86,0,0,0,3,0,0,0,65,0,20,0,0,0,97,0,199,0,51,0,178,0,166,0,14,0,80,0,124,0,175,0,21,0,83,0,82,0,133,0,50,0,185,0,0,0,199,0,46,0,58,0,0,0,11,0,29,0,0,0,28,0,200,0,103,0,57,0,144,0,0,0,169,0,0,0,205,0,0,0,0,0,0,0,0,0,212,0,37,0,0,0,183,0,0,0,0,0,156,0,60,0,138,0,3,0,139,0,233,0,142,0,147,0,215,0,224,0,251,0,116,0,189,0,46,0,13,0,134,0,163,0,122,0,0,0,0,0,182,0,154,0,160,0,50,0,163,0,13,0,231,0,0,0,133,0,94,0,177,0,77,0,95,0,219,0,139,0,187,0,60,0,15,0,144,0,219,0,147,0,230,0,154,0,60,0,0,0,0,0,0,0,0,0,0,0,237,0,90,0,61,0,0,0,98,0,0,0,0,0,0,0,16,0,15,0,142,0,246,0,0,0,55,0,139,0,199,0,0,0,210,0,183,0,128,0,63,0,0,0,171,0,115,0,191,0,144,0,61,0,221,0,175,0,96,0,123,0,226,0,98,0,1,0,214,0,2,0,0,0,142,0,166,0,128,0,205,0,138,0,202,0,85,0,92,0,68,0,113,0,226,0,72,0,107,0,0,0,211,0,115,0,19,0,4,0,0,0,24,0,0,0,110,0,138,0,231,0,179,0,141,0,252,0,224,0,213,0,0,0,47,0,0,0,0,0,156,0,0,0,38,0,137,0,225,0,196,0,149,0,80,0,239,0,175,0,161,0,0,0,0,0,0,0,234,0,0,0,242,0);
signal scenario_full  : scenario_type := (0,0,40,31,136,31,136,30,132,31,241,31,62,31,249,31,249,30,249,29,111,31,57,31,227,31,227,30,231,31,216,31,231,31,82,31,82,30,105,31,236,31,2,31,150,31,16,31,30,31,30,30,8,31,60,31,119,31,185,31,64,31,179,31,87,31,87,30,87,29,87,28,224,31,142,31,175,31,175,30,171,31,106,31,24,31,186,31,186,30,141,31,86,31,120,31,227,31,158,31,221,31,218,31,218,30,43,31,43,30,191,31,27,31,27,30,23,31,117,31,238,31,238,30,217,31,227,31,59,31,75,31,75,30,6,31,87,31,87,30,208,31,208,30,47,31,66,31,189,31,114,31,244,31,27,31,100,31,23,31,94,31,214,31,214,30,69,31,225,31,198,31,248,31,189,31,133,31,133,30,122,31,39,31,179,31,179,30,51,31,51,30,251,31,186,31,42,31,207,31,155,31,32,31,32,30,209,31,207,31,207,30,204,31,178,31,115,31,103,31,16,31,16,30,239,31,11,31,206,31,246,31,121,31,121,30,121,29,15,31,139,31,130,31,222,31,222,30,70,31,53,31,42,31,98,31,131,31,223,31,223,30,30,31,48,31,74,31,220,31,220,30,239,31,57,31,57,30,98,31,12,31,23,31,45,31,170,31,130,31,130,30,199,31,154,31,154,30,197,31,209,31,163,31,162,31,162,30,146,31,136,31,252,31,54,31,54,30,54,29,144,31,57,31,10,31,161,31,219,31,173,31,28,31,60,31,187,31,96,31,221,31,221,30,12,31,87,31,40,31,109,31,210,31,208,31,192,31,192,30,23,31,36,31,218,31,150,31,173,31,113,31,34,31,94,31,63,31,142,31,164,31,164,30,170,31,6,31,93,31,134,31,135,31,159,31,87,31,54,31,131,31,241,31,241,30,82,31,200,31,100,31,98,31,136,31,179,31,6,31,198,31,198,30,151,31,25,31,36,31,110,31,171,31,245,31,245,30,245,29,203,31,178,31,67,31,67,30,67,29,100,31,243,31,125,31,254,31,20,31,210,31,234,31,23,31,23,30,82,31,183,31,21,31,232,31,232,30,19,31,144,31,255,31,22,31,10,31,204,31,65,31,87,31,156,31,217,31,155,31,163,31,163,30,59,31,91,31,145,31,84,31,84,30,84,29,70,31,218,31,218,30,168,31,168,30,118,31,58,31,114,31,114,31,194,31,27,31,217,31,38,31,16,31,65,31,65,30,168,31,52,31,52,30,224,31,152,31,83,31,20,31,158,31,79,31,4,31,147,31,192,31,192,30,170,31,170,30,160,31,115,31,187,31,69,31,238,31,122,31,199,31,199,30,68,31,149,31,47,31,56,31,155,31,181,31,42,31,228,31,228,30,91,31,148,31,187,31,211,31,211,30,211,29,84,31,246,31,246,30,125,31,68,31,203,31,102,31,86,31,86,30,3,31,3,30,65,31,20,31,20,30,97,31,199,31,51,31,178,31,166,31,14,31,80,31,124,31,175,31,21,31,83,31,82,31,133,31,50,31,185,31,185,30,199,31,46,31,58,31,58,30,11,31,29,31,29,30,28,31,200,31,103,31,57,31,144,31,144,30,169,31,169,30,205,31,205,30,205,29,205,28,205,27,212,31,37,31,37,30,183,31,183,30,183,29,156,31,60,31,138,31,3,31,139,31,233,31,142,31,147,31,215,31,224,31,251,31,116,31,189,31,46,31,13,31,134,31,163,31,122,31,122,30,122,29,182,31,154,31,160,31,50,31,163,31,13,31,231,31,231,30,133,31,94,31,177,31,77,31,95,31,219,31,139,31,187,31,60,31,15,31,144,31,219,31,147,31,230,31,154,31,60,31,60,30,60,29,60,28,60,27,60,26,237,31,90,31,61,31,61,30,98,31,98,30,98,29,98,28,16,31,15,31,142,31,246,31,246,30,55,31,139,31,199,31,199,30,210,31,183,31,128,31,63,31,63,30,171,31,115,31,191,31,144,31,61,31,221,31,175,31,96,31,123,31,226,31,98,31,1,31,214,31,2,31,2,30,142,31,166,31,128,31,205,31,138,31,202,31,85,31,92,31,68,31,113,31,226,31,72,31,107,31,107,30,211,31,115,31,19,31,4,31,4,30,24,31,24,30,110,31,138,31,231,31,179,31,141,31,252,31,224,31,213,31,213,30,47,31,47,30,47,29,156,31,156,30,38,31,137,31,225,31,196,31,149,31,80,31,239,31,175,31,161,31,161,30,161,29,161,28,234,31,234,30,242,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
