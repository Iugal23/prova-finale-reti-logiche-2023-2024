-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 475;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (7,0,39,0,54,0,0,0,0,0,199,0,191,0,70,0,41,0,96,0,42,0,97,0,64,0,247,0,180,0,255,0,0,0,56,0,69,0,173,0,220,0,56,0,124,0,132,0,0,0,214,0,137,0,72,0,31,0,0,0,88,0,0,0,135,0,0,0,201,0,218,0,222,0,47,0,58,0,168,0,0,0,213,0,65,0,126,0,0,0,0,0,111,0,218,0,134,0,56,0,18,0,0,0,56,0,246,0,136,0,0,0,154,0,5,0,0,0,159,0,142,0,0,0,0,0,163,0,15,0,128,0,204,0,133,0,32,0,108,0,0,0,203,0,236,0,192,0,87,0,0,0,158,0,72,0,34,0,18,0,125,0,27,0,41,0,174,0,61,0,0,0,191,0,60,0,129,0,99,0,0,0,0,0,93,0,160,0,251,0,6,0,146,0,251,0,0,0,45,0,183,0,226,0,107,0,198,0,175,0,93,0,205,0,154,0,0,0,156,0,195,0,12,0,210,0,43,0,236,0,53,0,220,0,193,0,164,0,120,0,4,0,23,0,105,0,243,0,18,0,145,0,12,0,0,0,243,0,0,0,71,0,0,0,8,0,0,0,120,0,4,0,83,0,174,0,36,0,159,0,227,0,148,0,196,0,217,0,130,0,28,0,137,0,201,0,2,0,0,0,0,0,130,0,242,0,207,0,87,0,92,0,227,0,192,0,60,0,89,0,96,0,237,0,190,0,0,0,247,0,178,0,101,0,129,0,251,0,201,0,0,0,0,0,12,0,0,0,0,0,97,0,21,0,220,0,199,0,88,0,252,0,18,0,0,0,5,0,0,0,57,0,0,0,112,0,173,0,66,0,225,0,77,0,0,0,41,0,220,0,33,0,166,0,86,0,0,0,0,0,94,0,0,0,226,0,229,0,166,0,0,0,64,0,66,0,44,0,184,0,27,0,177,0,152,0,37,0,6,0,0,0,83,0,0,0,26,0,0,0,35,0,128,0,69,0,248,0,0,0,91,0,38,0,27,0,60,0,124,0,106,0,136,0,157,0,197,0,53,0,218,0,168,0,144,0,90,0,43,0,97,0,239,0,50,0,96,0,227,0,34,0,9,0,0,0,0,0,244,0,157,0,113,0,0,0,172,0,156,0,61,0,0,0,131,0,0,0,0,0,0,0,39,0,94,0,157,0,105,0,0,0,218,0,68,0,213,0,50,0,134,0,108,0,240,0,121,0,203,0,228,0,17,0,0,0,225,0,92,0,73,0,0,0,0,0,224,0,106,0,0,0,26,0,22,0,80,0,0,0,0,0,48,0,101,0,146,0,195,0,240,0,29,0,117,0,250,0,0,0,151,0,253,0,172,0,0,0,48,0,31,0,0,0,77,0,206,0,0,0,0,0,253,0,211,0,159,0,255,0,95,0,42,0,0,0,195,0,0,0,103,0,107,0,159,0,166,0,245,0,176,0,219,0,157,0,161,0,107,0,169,0,12,0,201,0,149,0,161,0,228,0,228,0,0,0,170,0,244,0,44,0,155,0,0,0,240,0,66,0,174,0,0,0,0,0,0,0,173,0,114,0,0,0,61,0,236,0,29,0,0,0,0,0,196,0,107,0,240,0,196,0,165,0,109,0,42,0,173,0,223,0,157,0,56,0,10,0,127,0,103,0,73,0,179,0,123,0,3,0,175,0,164,0,0,0,146,0,236,0,0,0,0,0,227,0,212,0,186,0,5,0,167,0,169,0,114,0,55,0,202,0,0,0,148,0,3,0,87,0,113,0,7,0,225,0,0,0,0,0,0,0,109,0,236,0,250,0,119,0,249,0,115,0,252,0,195,0,74,0,21,0,119,0,0,0,186,0,0,0,190,0,228,0,174,0,167,0,0,0,26,0,221,0,111,0,50,0,117,0,169,0,150,0,124,0,151,0,155,0,159,0,180,0,0,0,37,0,0,0,29,0,121,0,221,0,0,0,0,0,72,0,254,0,0,0,0,0,104,0,34,0,0,0,251,0,205,0,27,0,38,0,63,0,98,0,127,0,131,0,82,0,63,0,122,0,98,0,0,0,246,0,33,0,20,0,115,0,241,0,0,0,0,0,237,0,155,0,233,0,92,0,115,0,226,0,55,0,22,0);
signal scenario_full  : scenario_type := (7,31,39,31,54,31,54,30,54,29,199,31,191,31,70,31,41,31,96,31,42,31,97,31,64,31,247,31,180,31,255,31,255,30,56,31,69,31,173,31,220,31,56,31,124,31,132,31,132,30,214,31,137,31,72,31,31,31,31,30,88,31,88,30,135,31,135,30,201,31,218,31,222,31,47,31,58,31,168,31,168,30,213,31,65,31,126,31,126,30,126,29,111,31,218,31,134,31,56,31,18,31,18,30,56,31,246,31,136,31,136,30,154,31,5,31,5,30,159,31,142,31,142,30,142,29,163,31,15,31,128,31,204,31,133,31,32,31,108,31,108,30,203,31,236,31,192,31,87,31,87,30,158,31,72,31,34,31,18,31,125,31,27,31,41,31,174,31,61,31,61,30,191,31,60,31,129,31,99,31,99,30,99,29,93,31,160,31,251,31,6,31,146,31,251,31,251,30,45,31,183,31,226,31,107,31,198,31,175,31,93,31,205,31,154,31,154,30,156,31,195,31,12,31,210,31,43,31,236,31,53,31,220,31,193,31,164,31,120,31,4,31,23,31,105,31,243,31,18,31,145,31,12,31,12,30,243,31,243,30,71,31,71,30,8,31,8,30,120,31,4,31,83,31,174,31,36,31,159,31,227,31,148,31,196,31,217,31,130,31,28,31,137,31,201,31,2,31,2,30,2,29,130,31,242,31,207,31,87,31,92,31,227,31,192,31,60,31,89,31,96,31,237,31,190,31,190,30,247,31,178,31,101,31,129,31,251,31,201,31,201,30,201,29,12,31,12,30,12,29,97,31,21,31,220,31,199,31,88,31,252,31,18,31,18,30,5,31,5,30,57,31,57,30,112,31,173,31,66,31,225,31,77,31,77,30,41,31,220,31,33,31,166,31,86,31,86,30,86,29,94,31,94,30,226,31,229,31,166,31,166,30,64,31,66,31,44,31,184,31,27,31,177,31,152,31,37,31,6,31,6,30,83,31,83,30,26,31,26,30,35,31,128,31,69,31,248,31,248,30,91,31,38,31,27,31,60,31,124,31,106,31,136,31,157,31,197,31,53,31,218,31,168,31,144,31,90,31,43,31,97,31,239,31,50,31,96,31,227,31,34,31,9,31,9,30,9,29,244,31,157,31,113,31,113,30,172,31,156,31,61,31,61,30,131,31,131,30,131,29,131,28,39,31,94,31,157,31,105,31,105,30,218,31,68,31,213,31,50,31,134,31,108,31,240,31,121,31,203,31,228,31,17,31,17,30,225,31,92,31,73,31,73,30,73,29,224,31,106,31,106,30,26,31,22,31,80,31,80,30,80,29,48,31,101,31,146,31,195,31,240,31,29,31,117,31,250,31,250,30,151,31,253,31,172,31,172,30,48,31,31,31,31,30,77,31,206,31,206,30,206,29,253,31,211,31,159,31,255,31,95,31,42,31,42,30,195,31,195,30,103,31,107,31,159,31,166,31,245,31,176,31,219,31,157,31,161,31,107,31,169,31,12,31,201,31,149,31,161,31,228,31,228,31,228,30,170,31,244,31,44,31,155,31,155,30,240,31,66,31,174,31,174,30,174,29,174,28,173,31,114,31,114,30,61,31,236,31,29,31,29,30,29,29,196,31,107,31,240,31,196,31,165,31,109,31,42,31,173,31,223,31,157,31,56,31,10,31,127,31,103,31,73,31,179,31,123,31,3,31,175,31,164,31,164,30,146,31,236,31,236,30,236,29,227,31,212,31,186,31,5,31,167,31,169,31,114,31,55,31,202,31,202,30,148,31,3,31,87,31,113,31,7,31,225,31,225,30,225,29,225,28,109,31,236,31,250,31,119,31,249,31,115,31,252,31,195,31,74,31,21,31,119,31,119,30,186,31,186,30,190,31,228,31,174,31,167,31,167,30,26,31,221,31,111,31,50,31,117,31,169,31,150,31,124,31,151,31,155,31,159,31,180,31,180,30,37,31,37,30,29,31,121,31,221,31,221,30,221,29,72,31,254,31,254,30,254,29,104,31,34,31,34,30,251,31,205,31,27,31,38,31,63,31,98,31,127,31,131,31,82,31,63,31,122,31,98,31,98,30,246,31,33,31,20,31,115,31,241,31,241,30,241,29,237,31,155,31,233,31,92,31,115,31,226,31,55,31,22,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
