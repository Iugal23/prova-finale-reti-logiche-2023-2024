-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_121 is
end project_tb_121;

architecture project_tb_arch_121 of project_tb_121 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 823;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (27,0,0,0,0,0,226,0,150,0,115,0,19,0,14,0,30,0,216,0,0,0,135,0,251,0,145,0,65,0,0,0,151,0,38,0,0,0,7,0,50,0,221,0,152,0,49,0,40,0,87,0,2,0,223,0,141,0,163,0,36,0,224,0,0,0,236,0,204,0,164,0,155,0,0,0,5,0,164,0,13,0,49,0,152,0,102,0,249,0,229,0,63,0,0,0,58,0,176,0,59,0,201,0,0,0,0,0,2,0,135,0,170,0,21,0,25,0,171,0,47,0,0,0,158,0,0,0,242,0,0,0,59,0,135,0,0,0,7,0,0,0,0,0,123,0,0,0,0,0,0,0,169,0,0,0,46,0,205,0,232,0,42,0,205,0,149,0,16,0,35,0,145,0,0,0,50,0,0,0,0,0,140,0,0,0,229,0,0,0,142,0,247,0,110,0,0,0,82,0,189,0,84,0,199,0,67,0,9,0,210,0,0,0,20,0,243,0,156,0,227,0,0,0,131,0,155,0,214,0,237,0,38,0,0,0,104,0,150,0,221,0,102,0,211,0,11,0,185,0,190,0,87,0,39,0,237,0,39,0,67,0,70,0,173,0,0,0,0,0,197,0,230,0,0,0,39,0,76,0,95,0,0,0,0,0,151,0,155,0,70,0,23,0,214,0,158,0,46,0,0,0,0,0,0,0,112,0,114,0,0,0,171,0,211,0,79,0,32,0,124,0,29,0,0,0,196,0,132,0,105,0,0,0,115,0,71,0,62,0,194,0,0,0,0,0,45,0,0,0,231,0,232,0,0,0,154,0,0,0,14,0,169,0,26,0,0,0,240,0,150,0,34,0,127,0,113,0,182,0,212,0,0,0,0,0,95,0,0,0,236,0,233,0,0,0,0,0,223,0,65,0,229,0,0,0,5,0,147,0,0,0,175,0,197,0,174,0,55,0,67,0,183,0,26,0,82,0,144,0,167,0,74,0,102,0,0,0,0,0,221,0,229,0,162,0,178,0,224,0,93,0,175,0,170,0,245,0,0,0,231,0,0,0,28,0,255,0,193,0,138,0,127,0,131,0,143,0,0,0,109,0,126,0,86,0,94,0,172,0,139,0,172,0,208,0,21,0,147,0,113,0,169,0,183,0,0,0,88,0,135,0,204,0,34,0,201,0,41,0,109,0,145,0,27,0,200,0,0,0,146,0,252,0,172,0,161,0,43,0,247,0,37,0,37,0,0,0,199,0,184,0,0,0,171,0,92,0,107,0,0,0,6,0,50,0,242,0,0,0,105,0,111,0,39,0,47,0,0,0,0,0,44,0,127,0,237,0,149,0,230,0,80,0,0,0,0,0,0,0,26,0,70,0,191,0,92,0,229,0,74,0,0,0,0,0,210,0,59,0,193,0,0,0,140,0,99,0,82,0,223,0,179,0,223,0,93,0,0,0,2,0,173,0,215,0,0,0,219,0,116,0,230,0,42,0,0,0,194,0,123,0,139,0,119,0,139,0,83,0,38,0,0,0,10,0,248,0,164,0,0,0,217,0,37,0,93,0,117,0,254,0,158,0,70,0,153,0,208,0,216,0,40,0,0,0,148,0,214,0,100,0,55,0,95,0,101,0,184,0,0,0,168,0,171,0,0,0,0,0,34,0,0,0,66,0,189,0,237,0,112,0,158,0,249,0,184,0,239,0,0,0,0,0,146,0,79,0,186,0,215,0,66,0,46,0,0,0,203,0,11,0,15,0,19,0,250,0,40,0,0,0,0,0,0,0,77,0,20,0,155,0,138,0,22,0,246,0,225,0,69,0,227,0,198,0,9,0,0,0,121,0,125,0,0,0,0,0,131,0,41,0,102,0,0,0,225,0,62,0,4,0,182,0,41,0,50,0,229,0,60,0,49,0,221,0,66,0,76,0,125,0,188,0,226,0,68,0,57,0,217,0,86,0,105,0,212,0,198,0,0,0,0,0,100,0,198,0,39,0,207,0,10,0,162,0,40,0,0,0,0,0,147,0,178,0,193,0,40,0,221,0,242,0,226,0,35,0,85,0,209,0,0,0,144,0,11,0,92,0,237,0,13,0,220,0,65,0,135,0,20,0,9,0,190,0,97,0,238,0,132,0,102,0,0,0,192,0,219,0,16,0,72,0,206,0,0,0,22,0,117,0,24,0,74,0,206,0,0,0,33,0,78,0,109,0,196,0,91,0,20,0,175,0,189,0,47,0,165,0,95,0,0,0,75,0,0,0,0,0,118,0,250,0,0,0,247,0,97,0,130,0,54,0,223,0,63,0,88,0,217,0,141,0,107,0,0,0,0,0,142,0,0,0,26,0,42,0,55,0,229,0,40,0,0,0,156,0,0,0,0,0,74,0,0,0,0,0,0,0,217,0,117,0,210,0,32,0,77,0,131,0,13,0,135,0,110,0,0,0,84,0,84,0,142,0,0,0,43,0,0,0,87,0,183,0,54,0,78,0,173,0,247,0,35,0,0,0,253,0,25,0,102,0,67,0,39,0,0,0,0,0,151,0,1,0,213,0,2,0,152,0,66,0,26,0,147,0,77,0,82,0,38,0,157,0,145,0,0,0,101,0,15,0,189,0,192,0,129,0,70,0,0,0,241,0,133,0,252,0,0,0,70,0,77,0,0,0,219,0,250,0,37,0,235,0,3,0,0,0,149,0,0,0,194,0,0,0,50,0,210,0,73,0,59,0,44,0,116,0,0,0,16,0,0,0,136,0,123,0,31,0,95,0,88,0,0,0,0,0,161,0,36,0,35,0,21,0,229,0,140,0,7,0,48,0,123,0,83,0,177,0,0,0,179,0,251,0,28,0,170,0,133,0,0,0,12,0,34,0,205,0,90,0,17,0,44,0,15,0,62,0,124,0,136,0,193,0,98,0,0,0,101,0,0,0,88,0,0,0,172,0,89,0,90,0,0,0,79,0,230,0,173,0,9,0,35,0,44,0,191,0,201,0,172,0,104,0,213,0,28,0,88,0,37,0,164,0,48,0,114,0,175,0,96,0,132,0,0,0,191,0,144,0,72,0,11,0,112,0,196,0,33,0,8,0,153,0,199,0,217,0,201,0,0,0,93,0,136,0,134,0,0,0,0,0,205,0,12,0,122,0,242,0,152,0,154,0,117,0,155,0,126,0,0,0,56,0,57,0,153,0,155,0,116,0,0,0,0,0,181,0,203,0,7,0,94,0,252,0,175,0,230,0,0,0,29,0,247,0,130,0,180,0,132,0,70,0,215,0,0,0,129,0,137,0,229,0,0,0,33,0,0,0,241,0,251,0,146,0,124,0,0,0,130,0,171,0,138,0,0,0,0,0,56,0,0,0,231,0,15,0,24,0,0,0,57,0,60,0,141,0,47,0,162,0,114,0,96,0,0,0,0,0,0,0,60,0,7,0,0,0,246,0,121,0,144,0,135,0,0,0,7,0,0,0,0,0,245,0,0,0,114,0,116,0,0,0,183,0,229,0,207,0,0,0,75,0,145,0,24,0,140,0,99,0,179,0,102,0,108,0,247,0,0,0,0,0,0,0,215,0,0,0,243,0,9,0,122,0,0,0,58,0,74,0,0,0,124,0,243,0,179,0,0,0,101,0,173,0,220,0,14,0,71,0,190,0,5,0,124,0,60,0,143,0,0,0,149,0,197,0,112,0,2,0,183,0,0,0,54,0,0,0,237,0);
signal scenario_full  : scenario_type := (27,31,27,30,27,29,226,31,150,31,115,31,19,31,14,31,30,31,216,31,216,30,135,31,251,31,145,31,65,31,65,30,151,31,38,31,38,30,7,31,50,31,221,31,152,31,49,31,40,31,87,31,2,31,223,31,141,31,163,31,36,31,224,31,224,30,236,31,204,31,164,31,155,31,155,30,5,31,164,31,13,31,49,31,152,31,102,31,249,31,229,31,63,31,63,30,58,31,176,31,59,31,201,31,201,30,201,29,2,31,135,31,170,31,21,31,25,31,171,31,47,31,47,30,158,31,158,30,242,31,242,30,59,31,135,31,135,30,7,31,7,30,7,29,123,31,123,30,123,29,123,28,169,31,169,30,46,31,205,31,232,31,42,31,205,31,149,31,16,31,35,31,145,31,145,30,50,31,50,30,50,29,140,31,140,30,229,31,229,30,142,31,247,31,110,31,110,30,82,31,189,31,84,31,199,31,67,31,9,31,210,31,210,30,20,31,243,31,156,31,227,31,227,30,131,31,155,31,214,31,237,31,38,31,38,30,104,31,150,31,221,31,102,31,211,31,11,31,185,31,190,31,87,31,39,31,237,31,39,31,67,31,70,31,173,31,173,30,173,29,197,31,230,31,230,30,39,31,76,31,95,31,95,30,95,29,151,31,155,31,70,31,23,31,214,31,158,31,46,31,46,30,46,29,46,28,112,31,114,31,114,30,171,31,211,31,79,31,32,31,124,31,29,31,29,30,196,31,132,31,105,31,105,30,115,31,71,31,62,31,194,31,194,30,194,29,45,31,45,30,231,31,232,31,232,30,154,31,154,30,14,31,169,31,26,31,26,30,240,31,150,31,34,31,127,31,113,31,182,31,212,31,212,30,212,29,95,31,95,30,236,31,233,31,233,30,233,29,223,31,65,31,229,31,229,30,5,31,147,31,147,30,175,31,197,31,174,31,55,31,67,31,183,31,26,31,82,31,144,31,167,31,74,31,102,31,102,30,102,29,221,31,229,31,162,31,178,31,224,31,93,31,175,31,170,31,245,31,245,30,231,31,231,30,28,31,255,31,193,31,138,31,127,31,131,31,143,31,143,30,109,31,126,31,86,31,94,31,172,31,139,31,172,31,208,31,21,31,147,31,113,31,169,31,183,31,183,30,88,31,135,31,204,31,34,31,201,31,41,31,109,31,145,31,27,31,200,31,200,30,146,31,252,31,172,31,161,31,43,31,247,31,37,31,37,31,37,30,199,31,184,31,184,30,171,31,92,31,107,31,107,30,6,31,50,31,242,31,242,30,105,31,111,31,39,31,47,31,47,30,47,29,44,31,127,31,237,31,149,31,230,31,80,31,80,30,80,29,80,28,26,31,70,31,191,31,92,31,229,31,74,31,74,30,74,29,210,31,59,31,193,31,193,30,140,31,99,31,82,31,223,31,179,31,223,31,93,31,93,30,2,31,173,31,215,31,215,30,219,31,116,31,230,31,42,31,42,30,194,31,123,31,139,31,119,31,139,31,83,31,38,31,38,30,10,31,248,31,164,31,164,30,217,31,37,31,93,31,117,31,254,31,158,31,70,31,153,31,208,31,216,31,40,31,40,30,148,31,214,31,100,31,55,31,95,31,101,31,184,31,184,30,168,31,171,31,171,30,171,29,34,31,34,30,66,31,189,31,237,31,112,31,158,31,249,31,184,31,239,31,239,30,239,29,146,31,79,31,186,31,215,31,66,31,46,31,46,30,203,31,11,31,15,31,19,31,250,31,40,31,40,30,40,29,40,28,77,31,20,31,155,31,138,31,22,31,246,31,225,31,69,31,227,31,198,31,9,31,9,30,121,31,125,31,125,30,125,29,131,31,41,31,102,31,102,30,225,31,62,31,4,31,182,31,41,31,50,31,229,31,60,31,49,31,221,31,66,31,76,31,125,31,188,31,226,31,68,31,57,31,217,31,86,31,105,31,212,31,198,31,198,30,198,29,100,31,198,31,39,31,207,31,10,31,162,31,40,31,40,30,40,29,147,31,178,31,193,31,40,31,221,31,242,31,226,31,35,31,85,31,209,31,209,30,144,31,11,31,92,31,237,31,13,31,220,31,65,31,135,31,20,31,9,31,190,31,97,31,238,31,132,31,102,31,102,30,192,31,219,31,16,31,72,31,206,31,206,30,22,31,117,31,24,31,74,31,206,31,206,30,33,31,78,31,109,31,196,31,91,31,20,31,175,31,189,31,47,31,165,31,95,31,95,30,75,31,75,30,75,29,118,31,250,31,250,30,247,31,97,31,130,31,54,31,223,31,63,31,88,31,217,31,141,31,107,31,107,30,107,29,142,31,142,30,26,31,42,31,55,31,229,31,40,31,40,30,156,31,156,30,156,29,74,31,74,30,74,29,74,28,217,31,117,31,210,31,32,31,77,31,131,31,13,31,135,31,110,31,110,30,84,31,84,31,142,31,142,30,43,31,43,30,87,31,183,31,54,31,78,31,173,31,247,31,35,31,35,30,253,31,25,31,102,31,67,31,39,31,39,30,39,29,151,31,1,31,213,31,2,31,152,31,66,31,26,31,147,31,77,31,82,31,38,31,157,31,145,31,145,30,101,31,15,31,189,31,192,31,129,31,70,31,70,30,241,31,133,31,252,31,252,30,70,31,77,31,77,30,219,31,250,31,37,31,235,31,3,31,3,30,149,31,149,30,194,31,194,30,50,31,210,31,73,31,59,31,44,31,116,31,116,30,16,31,16,30,136,31,123,31,31,31,95,31,88,31,88,30,88,29,161,31,36,31,35,31,21,31,229,31,140,31,7,31,48,31,123,31,83,31,177,31,177,30,179,31,251,31,28,31,170,31,133,31,133,30,12,31,34,31,205,31,90,31,17,31,44,31,15,31,62,31,124,31,136,31,193,31,98,31,98,30,101,31,101,30,88,31,88,30,172,31,89,31,90,31,90,30,79,31,230,31,173,31,9,31,35,31,44,31,191,31,201,31,172,31,104,31,213,31,28,31,88,31,37,31,164,31,48,31,114,31,175,31,96,31,132,31,132,30,191,31,144,31,72,31,11,31,112,31,196,31,33,31,8,31,153,31,199,31,217,31,201,31,201,30,93,31,136,31,134,31,134,30,134,29,205,31,12,31,122,31,242,31,152,31,154,31,117,31,155,31,126,31,126,30,56,31,57,31,153,31,155,31,116,31,116,30,116,29,181,31,203,31,7,31,94,31,252,31,175,31,230,31,230,30,29,31,247,31,130,31,180,31,132,31,70,31,215,31,215,30,129,31,137,31,229,31,229,30,33,31,33,30,241,31,251,31,146,31,124,31,124,30,130,31,171,31,138,31,138,30,138,29,56,31,56,30,231,31,15,31,24,31,24,30,57,31,60,31,141,31,47,31,162,31,114,31,96,31,96,30,96,29,96,28,60,31,7,31,7,30,246,31,121,31,144,31,135,31,135,30,7,31,7,30,7,29,245,31,245,30,114,31,116,31,116,30,183,31,229,31,207,31,207,30,75,31,145,31,24,31,140,31,99,31,179,31,102,31,108,31,247,31,247,30,247,29,247,28,215,31,215,30,243,31,9,31,122,31,122,30,58,31,74,31,74,30,124,31,243,31,179,31,179,30,101,31,173,31,220,31,14,31,71,31,190,31,5,31,124,31,60,31,143,31,143,30,149,31,197,31,112,31,2,31,183,31,183,30,54,31,54,30,237,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
