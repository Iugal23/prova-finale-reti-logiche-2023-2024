-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 352;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (232,0,194,0,0,0,247,0,0,0,0,0,88,0,28,0,127,0,0,0,177,0,248,0,21,0,76,0,0,0,175,0,46,0,195,0,200,0,16,0,0,0,163,0,0,0,78,0,0,0,183,0,0,0,106,0,0,0,231,0,0,0,22,0,0,0,0,0,18,0,182,0,145,0,187,0,33,0,201,0,150,0,161,0,216,0,139,0,131,0,38,0,248,0,92,0,84,0,74,0,199,0,241,0,0,0,147,0,184,0,178,0,49,0,0,0,76,0,122,0,124,0,242,0,184,0,239,0,25,0,58,0,2,0,219,0,0,0,145,0,115,0,239,0,0,0,131,0,255,0,167,0,204,0,92,0,189,0,0,0,11,0,2,0,76,0,143,0,97,0,39,0,241,0,0,0,205,0,0,0,0,0,0,0,30,0,85,0,11,0,39,0,52,0,20,0,147,0,74,0,120,0,186,0,177,0,49,0,236,0,0,0,0,0,0,0,164,0,126,0,239,0,71,0,10,0,8,0,152,0,127,0,158,0,0,0,18,0,0,0,0,0,101,0,0,0,212,0,83,0,0,0,132,0,44,0,80,0,37,0,0,0,75,0,220,0,239,0,228,0,31,0,0,0,4,0,0,0,240,0,0,0,140,0,0,0,105,0,167,0,37,0,0,0,221,0,0,0,162,0,190,0,41,0,130,0,22,0,56,0,178,0,120,0,0,0,219,0,85,0,95,0,108,0,219,0,251,0,35,0,108,0,92,0,0,0,115,0,254,0,41,0,17,0,154,0,0,0,0,0,168,0,170,0,120,0,0,0,115,0,101,0,211,0,206,0,17,0,136,0,21,0,8,0,215,0,209,0,210,0,176,0,0,0,247,0,0,0,139,0,8,0,0,0,86,0,254,0,141,0,99,0,7,0,199,0,102,0,181,0,0,0,220,0,0,0,66,0,0,0,0,0,239,0,115,0,0,0,0,0,53,0,0,0,153,0,225,0,240,0,97,0,70,0,209,0,197,0,112,0,121,0,0,0,32,0,0,0,0,0,47,0,0,0,241,0,0,0,51,0,5,0,227,0,81,0,179,0,142,0,0,0,15,0,153,0,181,0,0,0,0,0,198,0,242,0,13,0,55,0,108,0,61,0,56,0,0,0,140,0,153,0,161,0,5,0,0,0,0,0,58,0,61,0,22,0,165,0,194,0,46,0,138,0,150,0,12,0,0,0,95,0,0,0,52,0,148,0,0,0,0,0,92,0,210,0,75,0,215,0,139,0,0,0,53,0,204,0,24,0,11,0,169,0,154,0,186,0,0,0,162,0,0,0,106,0,126,0,179,0,108,0,229,0,0,0,61,0,4,0,220,0,25,0,114,0,68,0,38,0,41,0,0,0,189,0,197,0,196,0,43,0,0,0,26,0,210,0,115,0,165,0,0,0,0,0,41,0,68,0,235,0,0,0,241,0,188,0,137,0,0,0,51,0,161,0,192,0,88,0,28,0,0,0,0,0,175,0,232,0,0,0,53,0,163,0,108,0,15,0,37,0,175,0,164,0,67,0,157,0,2,0,0,0,67,0,168,0,36,0,48,0,63,0);
signal scenario_full  : scenario_type := (232,31,194,31,194,30,247,31,247,30,247,29,88,31,28,31,127,31,127,30,177,31,248,31,21,31,76,31,76,30,175,31,46,31,195,31,200,31,16,31,16,30,163,31,163,30,78,31,78,30,183,31,183,30,106,31,106,30,231,31,231,30,22,31,22,30,22,29,18,31,182,31,145,31,187,31,33,31,201,31,150,31,161,31,216,31,139,31,131,31,38,31,248,31,92,31,84,31,74,31,199,31,241,31,241,30,147,31,184,31,178,31,49,31,49,30,76,31,122,31,124,31,242,31,184,31,239,31,25,31,58,31,2,31,219,31,219,30,145,31,115,31,239,31,239,30,131,31,255,31,167,31,204,31,92,31,189,31,189,30,11,31,2,31,76,31,143,31,97,31,39,31,241,31,241,30,205,31,205,30,205,29,205,28,30,31,85,31,11,31,39,31,52,31,20,31,147,31,74,31,120,31,186,31,177,31,49,31,236,31,236,30,236,29,236,28,164,31,126,31,239,31,71,31,10,31,8,31,152,31,127,31,158,31,158,30,18,31,18,30,18,29,101,31,101,30,212,31,83,31,83,30,132,31,44,31,80,31,37,31,37,30,75,31,220,31,239,31,228,31,31,31,31,30,4,31,4,30,240,31,240,30,140,31,140,30,105,31,167,31,37,31,37,30,221,31,221,30,162,31,190,31,41,31,130,31,22,31,56,31,178,31,120,31,120,30,219,31,85,31,95,31,108,31,219,31,251,31,35,31,108,31,92,31,92,30,115,31,254,31,41,31,17,31,154,31,154,30,154,29,168,31,170,31,120,31,120,30,115,31,101,31,211,31,206,31,17,31,136,31,21,31,8,31,215,31,209,31,210,31,176,31,176,30,247,31,247,30,139,31,8,31,8,30,86,31,254,31,141,31,99,31,7,31,199,31,102,31,181,31,181,30,220,31,220,30,66,31,66,30,66,29,239,31,115,31,115,30,115,29,53,31,53,30,153,31,225,31,240,31,97,31,70,31,209,31,197,31,112,31,121,31,121,30,32,31,32,30,32,29,47,31,47,30,241,31,241,30,51,31,5,31,227,31,81,31,179,31,142,31,142,30,15,31,153,31,181,31,181,30,181,29,198,31,242,31,13,31,55,31,108,31,61,31,56,31,56,30,140,31,153,31,161,31,5,31,5,30,5,29,58,31,61,31,22,31,165,31,194,31,46,31,138,31,150,31,12,31,12,30,95,31,95,30,52,31,148,31,148,30,148,29,92,31,210,31,75,31,215,31,139,31,139,30,53,31,204,31,24,31,11,31,169,31,154,31,186,31,186,30,162,31,162,30,106,31,126,31,179,31,108,31,229,31,229,30,61,31,4,31,220,31,25,31,114,31,68,31,38,31,41,31,41,30,189,31,197,31,196,31,43,31,43,30,26,31,210,31,115,31,165,31,165,30,165,29,41,31,68,31,235,31,235,30,241,31,188,31,137,31,137,30,51,31,161,31,192,31,88,31,28,31,28,30,28,29,175,31,232,31,232,30,53,31,163,31,108,31,15,31,37,31,175,31,164,31,67,31,157,31,2,31,2,30,67,31,168,31,36,31,48,31,63,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
