-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_502 is
end project_tb_502;

architecture project_tb_arch_502 of project_tb_502 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 798;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,0,0,0,0,110,0,196,0,90,0,97,0,143,0,0,0,128,0,56,0,88,0,56,0,1,0,94,0,61,0,211,0,0,0,229,0,12,0,32,0,106,0,0,0,159,0,233,0,0,0,201,0,123,0,0,0,42,0,184,0,120,0,0,0,24,0,14,0,0,0,0,0,0,0,70,0,209,0,247,0,174,0,127,0,0,0,3,0,0,0,224,0,1,0,0,0,191,0,253,0,0,0,22,0,202,0,204,0,191,0,107,0,215,0,0,0,0,0,156,0,136,0,24,0,207,0,244,0,50,0,135,0,228,0,0,0,252,0,0,0,0,0,186,0,152,0,215,0,0,0,167,0,12,0,117,0,4,0,0,0,155,0,19,0,166,0,33,0,1,0,0,0,113,0,169,0,231,0,141,0,131,0,9,0,53,0,40,0,148,0,203,0,0,0,104,0,0,0,0,0,104,0,104,0,255,0,131,0,245,0,0,0,229,0,199,0,68,0,74,0,84,0,0,0,134,0,203,0,162,0,0,0,12,0,27,0,61,0,140,0,0,0,237,0,189,0,249,0,0,0,77,0,112,0,111,0,166,0,110,0,214,0,105,0,77,0,0,0,45,0,226,0,46,0,66,0,140,0,0,0,123,0,217,0,0,0,48,0,99,0,140,0,0,0,0,0,113,0,0,0,129,0,29,0,40,0,82,0,68,0,217,0,220,0,79,0,250,0,32,0,10,0,43,0,237,0,194,0,213,0,156,0,0,0,123,0,6,0,0,0,235,0,0,0,0,0,139,0,225,0,0,0,81,0,150,0,212,0,223,0,87,0,52,0,55,0,218,0,197,0,169,0,60,0,236,0,135,0,15,0,218,0,21,0,248,0,6,0,0,0,122,0,76,0,113,0,207,0,17,0,5,0,198,0,190,0,5,0,76,0,138,0,169,0,0,0,150,0,40,0,38,0,0,0,0,0,138,0,20,0,94,0,47,0,96,0,95,0,212,0,102,0,251,0,0,0,58,0,220,0,198,0,141,0,139,0,31,0,94,0,62,0,118,0,0,0,150,0,247,0,150,0,25,0,245,0,10,0,160,0,0,0,248,0,0,0,133,0,124,0,179,0,39,0,0,0,240,0,0,0,129,0,124,0,36,0,40,0,20,0,0,0,55,0,201,0,143,0,246,0,116,0,192,0,130,0,114,0,8,0,0,0,224,0,0,0,241,0,51,0,29,0,0,0,174,0,34,0,255,0,39,0,0,0,0,0,95,0,0,0,0,0,231,0,79,0,235,0,130,0,33,0,236,0,171,0,155,0,25,0,188,0,0,0,0,0,0,0,0,0,69,0,176,0,59,0,0,0,246,0,187,0,77,0,0,0,176,0,220,0,43,0,208,0,57,0,40,0,0,0,166,0,189,0,165,0,0,0,141,0,65,0,120,0,101,0,175,0,32,0,0,0,195,0,0,0,168,0,239,0,0,0,10,0,56,0,208,0,0,0,214,0,0,0,105,0,127,0,0,0,61,0,150,0,0,0,102,0,92,0,83,0,253,0,72,0,0,0,0,0,0,0,73,0,192,0,28,0,62,0,131,0,0,0,0,0,101,0,0,0,0,0,0,0,39,0,0,0,97,0,160,0,229,0,154,0,176,0,100,0,100,0,255,0,217,0,224,0,212,0,3,0,94,0,137,0,24,0,6,0,98,0,79,0,100,0,124,0,14,0,32,0,0,0,0,0,30,0,7,0,23,0,146,0,108,0,0,0,252,0,90,0,133,0,182,0,7,0,115,0,39,0,146,0,195,0,27,0,1,0,149,0,128,0,24,0,27,0,25,0,10,0,208,0,142,0,18,0,0,0,0,0,87,0,0,0,3,0,138,0,26,0,196,0,88,0,0,0,0,0,0,0,33,0,128,0,77,0,87,0,0,0,213,0,221,0,51,0,0,0,0,0,0,0,82,0,132,0,0,0,0,0,192,0,97,0,230,0,56,0,213,0,143,0,123,0,102,0,248,0,141,0,42,0,50,0,135,0,6,0,185,0,0,0,24,0,237,0,31,0,0,0,182,0,84,0,0,0,0,0,182,0,191,0,0,0,214,0,115,0,105,0,93,0,62,0,145,0,0,0,0,0,13,0,64,0,183,0,40,0,10,0,250,0,127,0,105,0,188,0,106,0,0,0,218,0,34,0,93,0,234,0,126,0,145,0,208,0,80,0,126,0,83,0,0,0,0,0,137,0,239,0,145,0,83,0,12,0,101,0,100,0,9,0,20,0,0,0,0,0,154,0,107,0,0,0,113,0,80,0,0,0,138,0,206,0,174,0,49,0,0,0,0,0,46,0,162,0,62,0,239,0,26,0,0,0,0,0,102,0,0,0,0,0,104,0,0,0,89,0,0,0,68,0,77,0,0,0,156,0,210,0,10,0,196,0,0,0,122,0,93,0,254,0,162,0,204,0,42,0,9,0,0,0,240,0,241,0,219,0,0,0,167,0,255,0,39,0,229,0,22,0,120,0,0,0,133,0,137,0,234,0,0,0,60,0,179,0,0,0,133,0,0,0,0,0,134,0,0,0,29,0,138,0,216,0,107,0,215,0,161,0,111,0,156,0,147,0,188,0,15,0,89,0,56,0,229,0,69,0,148,0,172,0,0,0,133,0,197,0,75,0,125,0,115,0,171,0,0,0,154,0,0,0,0,0,224,0,28,0,42,0,198,0,129,0,101,0,86,0,0,0,0,0,54,0,217,0,58,0,2,0,104,0,176,0,166,0,80,0,0,0,7,0,185,0,55,0,201,0,0,0,203,0,0,0,82,0,0,0,4,0,0,0,0,0,254,0,1,0,96,0,23,0,135,0,168,0,203,0,98,0,0,0,189,0,77,0,19,0,11,0,41,0,100,0,71,0,204,0,23,0,0,0,122,0,71,0,25,0,0,0,0,0,87,0,250,0,207,0,0,0,0,0,137,0,113,0,152,0,62,0,0,0,102,0,7,0,0,0,148,0,72,0,167,0,9,0,11,0,33,0,227,0,96,0,0,0,191,0,225,0,0,0,0,0,75,0,65,0,141,0,88,0,147,0,70,0,125,0,216,0,203,0,0,0,30,0,71,0,227,0,0,0,0,0,18,0,21,0,186,0,0,0,199,0,144,0,173,0,57,0,179,0,16,0,0,0,0,0,0,0,0,0,48,0,112,0,0,0,0,0,209,0,118,0,146,0,0,0,119,0,139,0,114,0,231,0,227,0,25,0,17,0,0,0,30,0,240,0,122,0,24,0,130,0,43,0,158,0,225,0,63,0,116,0,148,0,127,0,83,0,208,0,147,0,0,0,87,0,0,0,17,0,219,0,152,0,137,0,69,0,250,0,189,0,63,0,0,0,74,0,76,0,30,0,11,0,224,0,70,0,0,0,0,0,143,0,7,0,203,0,211,0,154,0,229,0,0,0,0,0,229,0,47,0,122,0,108,0,0,0,0,0,0,0,247,0,139,0,35,0,180,0,94,0,153,0,107,0,0,0,127,0,30,0,0,0,54,0,118,0,64,0,213,0,144,0,0,0,200,0,78,0,76,0,201,0,111,0,172,0);
signal scenario_full  : scenario_type := (0,0,0,0,0,0,0,0,110,31,196,31,90,31,97,31,143,31,143,30,128,31,56,31,88,31,56,31,1,31,94,31,61,31,211,31,211,30,229,31,12,31,32,31,106,31,106,30,159,31,233,31,233,30,201,31,123,31,123,30,42,31,184,31,120,31,120,30,24,31,14,31,14,30,14,29,14,28,70,31,209,31,247,31,174,31,127,31,127,30,3,31,3,30,224,31,1,31,1,30,191,31,253,31,253,30,22,31,202,31,204,31,191,31,107,31,215,31,215,30,215,29,156,31,136,31,24,31,207,31,244,31,50,31,135,31,228,31,228,30,252,31,252,30,252,29,186,31,152,31,215,31,215,30,167,31,12,31,117,31,4,31,4,30,155,31,19,31,166,31,33,31,1,31,1,30,113,31,169,31,231,31,141,31,131,31,9,31,53,31,40,31,148,31,203,31,203,30,104,31,104,30,104,29,104,31,104,31,255,31,131,31,245,31,245,30,229,31,199,31,68,31,74,31,84,31,84,30,134,31,203,31,162,31,162,30,12,31,27,31,61,31,140,31,140,30,237,31,189,31,249,31,249,30,77,31,112,31,111,31,166,31,110,31,214,31,105,31,77,31,77,30,45,31,226,31,46,31,66,31,140,31,140,30,123,31,217,31,217,30,48,31,99,31,140,31,140,30,140,29,113,31,113,30,129,31,29,31,40,31,82,31,68,31,217,31,220,31,79,31,250,31,32,31,10,31,43,31,237,31,194,31,213,31,156,31,156,30,123,31,6,31,6,30,235,31,235,30,235,29,139,31,225,31,225,30,81,31,150,31,212,31,223,31,87,31,52,31,55,31,218,31,197,31,169,31,60,31,236,31,135,31,15,31,218,31,21,31,248,31,6,31,6,30,122,31,76,31,113,31,207,31,17,31,5,31,198,31,190,31,5,31,76,31,138,31,169,31,169,30,150,31,40,31,38,31,38,30,38,29,138,31,20,31,94,31,47,31,96,31,95,31,212,31,102,31,251,31,251,30,58,31,220,31,198,31,141,31,139,31,31,31,94,31,62,31,118,31,118,30,150,31,247,31,150,31,25,31,245,31,10,31,160,31,160,30,248,31,248,30,133,31,124,31,179,31,39,31,39,30,240,31,240,30,129,31,124,31,36,31,40,31,20,31,20,30,55,31,201,31,143,31,246,31,116,31,192,31,130,31,114,31,8,31,8,30,224,31,224,30,241,31,51,31,29,31,29,30,174,31,34,31,255,31,39,31,39,30,39,29,95,31,95,30,95,29,231,31,79,31,235,31,130,31,33,31,236,31,171,31,155,31,25,31,188,31,188,30,188,29,188,28,188,27,69,31,176,31,59,31,59,30,246,31,187,31,77,31,77,30,176,31,220,31,43,31,208,31,57,31,40,31,40,30,166,31,189,31,165,31,165,30,141,31,65,31,120,31,101,31,175,31,32,31,32,30,195,31,195,30,168,31,239,31,239,30,10,31,56,31,208,31,208,30,214,31,214,30,105,31,127,31,127,30,61,31,150,31,150,30,102,31,92,31,83,31,253,31,72,31,72,30,72,29,72,28,73,31,192,31,28,31,62,31,131,31,131,30,131,29,101,31,101,30,101,29,101,28,39,31,39,30,97,31,160,31,229,31,154,31,176,31,100,31,100,31,255,31,217,31,224,31,212,31,3,31,94,31,137,31,24,31,6,31,98,31,79,31,100,31,124,31,14,31,32,31,32,30,32,29,30,31,7,31,23,31,146,31,108,31,108,30,252,31,90,31,133,31,182,31,7,31,115,31,39,31,146,31,195,31,27,31,1,31,149,31,128,31,24,31,27,31,25,31,10,31,208,31,142,31,18,31,18,30,18,29,87,31,87,30,3,31,138,31,26,31,196,31,88,31,88,30,88,29,88,28,33,31,128,31,77,31,87,31,87,30,213,31,221,31,51,31,51,30,51,29,51,28,82,31,132,31,132,30,132,29,192,31,97,31,230,31,56,31,213,31,143,31,123,31,102,31,248,31,141,31,42,31,50,31,135,31,6,31,185,31,185,30,24,31,237,31,31,31,31,30,182,31,84,31,84,30,84,29,182,31,191,31,191,30,214,31,115,31,105,31,93,31,62,31,145,31,145,30,145,29,13,31,64,31,183,31,40,31,10,31,250,31,127,31,105,31,188,31,106,31,106,30,218,31,34,31,93,31,234,31,126,31,145,31,208,31,80,31,126,31,83,31,83,30,83,29,137,31,239,31,145,31,83,31,12,31,101,31,100,31,9,31,20,31,20,30,20,29,154,31,107,31,107,30,113,31,80,31,80,30,138,31,206,31,174,31,49,31,49,30,49,29,46,31,162,31,62,31,239,31,26,31,26,30,26,29,102,31,102,30,102,29,104,31,104,30,89,31,89,30,68,31,77,31,77,30,156,31,210,31,10,31,196,31,196,30,122,31,93,31,254,31,162,31,204,31,42,31,9,31,9,30,240,31,241,31,219,31,219,30,167,31,255,31,39,31,229,31,22,31,120,31,120,30,133,31,137,31,234,31,234,30,60,31,179,31,179,30,133,31,133,30,133,29,134,31,134,30,29,31,138,31,216,31,107,31,215,31,161,31,111,31,156,31,147,31,188,31,15,31,89,31,56,31,229,31,69,31,148,31,172,31,172,30,133,31,197,31,75,31,125,31,115,31,171,31,171,30,154,31,154,30,154,29,224,31,28,31,42,31,198,31,129,31,101,31,86,31,86,30,86,29,54,31,217,31,58,31,2,31,104,31,176,31,166,31,80,31,80,30,7,31,185,31,55,31,201,31,201,30,203,31,203,30,82,31,82,30,4,31,4,30,4,29,254,31,1,31,96,31,23,31,135,31,168,31,203,31,98,31,98,30,189,31,77,31,19,31,11,31,41,31,100,31,71,31,204,31,23,31,23,30,122,31,71,31,25,31,25,30,25,29,87,31,250,31,207,31,207,30,207,29,137,31,113,31,152,31,62,31,62,30,102,31,7,31,7,30,148,31,72,31,167,31,9,31,11,31,33,31,227,31,96,31,96,30,191,31,225,31,225,30,225,29,75,31,65,31,141,31,88,31,147,31,70,31,125,31,216,31,203,31,203,30,30,31,71,31,227,31,227,30,227,29,18,31,21,31,186,31,186,30,199,31,144,31,173,31,57,31,179,31,16,31,16,30,16,29,16,28,16,27,48,31,112,31,112,30,112,29,209,31,118,31,146,31,146,30,119,31,139,31,114,31,231,31,227,31,25,31,17,31,17,30,30,31,240,31,122,31,24,31,130,31,43,31,158,31,225,31,63,31,116,31,148,31,127,31,83,31,208,31,147,31,147,30,87,31,87,30,17,31,219,31,152,31,137,31,69,31,250,31,189,31,63,31,63,30,74,31,76,31,30,31,11,31,224,31,70,31,70,30,70,29,143,31,7,31,203,31,211,31,154,31,229,31,229,30,229,29,229,31,47,31,122,31,108,31,108,30,108,29,108,28,247,31,139,31,35,31,180,31,94,31,153,31,107,31,107,30,127,31,30,31,30,30,54,31,118,31,64,31,213,31,144,31,144,30,200,31,78,31,76,31,201,31,111,31,172,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
