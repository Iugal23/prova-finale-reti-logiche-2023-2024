-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 716;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (48,0,56,0,224,0,66,0,211,0,230,0,160,0,169,0,143,0,8,0,0,0,127,0,10,0,93,0,18,0,88,0,125,0,241,0,0,0,197,0,0,0,0,0,179,0,121,0,0,0,0,0,19,0,0,0,2,0,175,0,0,0,154,0,178,0,89,0,87,0,0,0,65,0,0,0,248,0,30,0,241,0,0,0,44,0,42,0,151,0,0,0,238,0,216,0,202,0,0,0,16,0,19,0,104,0,219,0,0,0,45,0,231,0,146,0,77,0,195,0,130,0,0,0,149,0,46,0,102,0,0,0,203,0,59,0,72,0,45,0,239,0,159,0,143,0,186,0,99,0,160,0,0,0,37,0,118,0,7,0,239,0,198,0,236,0,134,0,151,0,48,0,23,0,0,0,152,0,38,0,142,0,184,0,94,0,114,0,241,0,56,0,0,0,0,0,0,0,152,0,231,0,78,0,40,0,120,0,0,0,0,0,0,0,143,0,0,0,42,0,63,0,36,0,70,0,102,0,154,0,83,0,137,0,242,0,196,0,48,0,16,0,78,0,0,0,220,0,162,0,0,0,166,0,224,0,253,0,220,0,36,0,157,0,155,0,182,0,0,0,0,0,76,0,135,0,195,0,2,0,0,0,244,0,58,0,96,0,157,0,0,0,0,0,147,0,0,0,0,0,0,0,252,0,236,0,251,0,0,0,117,0,0,0,82,0,13,0,189,0,68,0,230,0,0,0,58,0,159,0,0,0,55,0,0,0,0,0,178,0,208,0,0,0,194,0,103,0,101,0,24,0,0,0,148,0,99,0,81,0,176,0,5,0,59,0,217,0,114,0,14,0,205,0,36,0,159,0,98,0,73,0,90,0,232,0,24,0,192,0,1,0,134,0,135,0,96,0,144,0,243,0,2,0,176,0,0,0,235,0,203,0,252,0,13,0,0,0,0,0,71,0,159,0,205,0,63,0,230,0,154,0,235,0,140,0,221,0,238,0,0,0,101,0,234,0,0,0,23,0,114,0,32,0,218,0,0,0,0,0,223,0,105,0,4,0,31,0,54,0,123,0,0,0,178,0,0,0,105,0,68,0,40,0,2,0,32,0,53,0,2,0,18,0,134,0,183,0,54,0,0,0,234,0,108,0,172,0,47,0,228,0,177,0,24,0,127,0,176,0,0,0,0,0,21,0,142,0,43,0,153,0,0,0,0,0,176,0,70,0,193,0,0,0,225,0,237,0,236,0,213,0,125,0,178,0,120,0,250,0,219,0,62,0,228,0,12,0,35,0,29,0,89,0,186,0,28,0,0,0,0,0,34,0,29,0,45,0,93,0,96,0,23,0,29,0,248,0,0,0,0,0,229,0,168,0,0,0,165,0,0,0,206,0,245,0,229,0,114,0,87,0,11,0,0,0,1,0,66,0,196,0,87,0,0,0,114,0,185,0,161,0,243,0,120,0,74,0,217,0,72,0,14,0,156,0,64,0,147,0,107,0,241,0,83,0,233,0,73,0,114,0,54,0,49,0,183,0,185,0,29,0,115,0,23,0,181,0,161,0,71,0,166,0,31,0,0,0,0,0,73,0,0,0,0,0,34,0,128,0,28,0,0,0,124,0,0,0,143,0,7,0,170,0,0,0,0,0,0,0,238,0,76,0,166,0,155,0,187,0,113,0,0,0,94,0,43,0,40,0,204,0,59,0,0,0,0,0,0,0,169,0,122,0,0,0,0,0,103,0,88,0,50,0,52,0,211,0,218,0,248,0,42,0,0,0,8,0,1,0,111,0,206,0,29,0,95,0,95,0,155,0,242,0,252,0,88,0,208,0,62,0,211,0,0,0,209,0,32,0,120,0,231,0,117,0,79,0,63,0,137,0,35,0,57,0,157,0,214,0,185,0,104,0,5,0,0,0,107,0,60,0,0,0,68,0,53,0,149,0,51,0,50,0,155,0,65,0,108,0,253,0,117,0,197,0,0,0,0,0,0,0,125,0,206,0,181,0,184,0,98,0,174,0,0,0,101,0,72,0,0,0,81,0,251,0,0,0,13,0,0,0,238,0,29,0,178,0,181,0,32,0,32,0,12,0,0,0,161,0,197,0,0,0,176,0,183,0,66,0,79,0,153,0,0,0,228,0,219,0,116,0,0,0,55,0,0,0,74,0,44,0,138,0,40,0,192,0,112,0,162,0,207,0,196,0,190,0,72,0,128,0,34,0,43,0,0,0,0,0,16,0,0,0,19,0,129,0,241,0,167,0,121,0,179,0,250,0,6,0,87,0,0,0,114,0,8,0,63,0,115,0,23,0,55,0,205,0,0,0,200,0,74,0,0,0,0,0,212,0,55,0,118,0,0,0,0,0,0,0,158,0,156,0,201,0,91,0,0,0,138,0,5,0,97,0,41,0,144,0,0,0,200,0,231,0,160,0,0,0,136,0,0,0,199,0,67,0,0,0,154,0,202,0,0,0,92,0,54,0,105,0,112,0,179,0,55,0,0,0,41,0,0,0,87,0,198,0,6,0,252,0,0,0,0,0,71,0,110,0,113,0,86,0,0,0,45,0,146,0,0,0,190,0,24,0,0,0,83,0,14,0,123,0,123,0,0,0,239,0,3,0,0,0,122,0,228,0,176,0,15,0,239,0,0,0,151,0,18,0,64,0,0,0,117,0,19,0,186,0,204,0,54,0,183,0,0,0,0,0,151,0,7,0,135,0,102,0,72,0,182,0,69,0,0,0,184,0,110,0,0,0,6,0,126,0,224,0,0,0,222,0,50,0,0,0,0,0,61,0,139,0,0,0,72,0,223,0,119,0,44,0,130,0,218,0,82,0,4,0,0,0,0,0,71,0,116,0,81,0,15,0,188,0,170,0,0,0,62,0,47,0,21,0,0,0,160,0,220,0,222,0,0,0,107,0,235,0,109,0,85,0,0,0,161,0,11,0,193,0,219,0,223,0,138,0,105,0,156,0,178,0,136,0,138,0,36,0,45,0,0,0,0,0,66,0,91,0,0,0,230,0,0,0,0,0,71,0,95,0,105,0,66,0,91,0,207,0,205,0,0,0,0,0,109,0,27,0,142,0,96,0,0,0,111,0,132,0,0,0,229,0,240,0,253,0,127,0,223,0,164,0,0,0,0,0,0,0,0,0,228,0,132,0,201,0,211,0,58,0,4,0,0,0,0,0,71,0,40,0,0,0,162,0,175,0,0,0,0,0,88,0);
signal scenario_full  : scenario_type := (48,31,56,31,224,31,66,31,211,31,230,31,160,31,169,31,143,31,8,31,8,30,127,31,10,31,93,31,18,31,88,31,125,31,241,31,241,30,197,31,197,30,197,29,179,31,121,31,121,30,121,29,19,31,19,30,2,31,175,31,175,30,154,31,178,31,89,31,87,31,87,30,65,31,65,30,248,31,30,31,241,31,241,30,44,31,42,31,151,31,151,30,238,31,216,31,202,31,202,30,16,31,19,31,104,31,219,31,219,30,45,31,231,31,146,31,77,31,195,31,130,31,130,30,149,31,46,31,102,31,102,30,203,31,59,31,72,31,45,31,239,31,159,31,143,31,186,31,99,31,160,31,160,30,37,31,118,31,7,31,239,31,198,31,236,31,134,31,151,31,48,31,23,31,23,30,152,31,38,31,142,31,184,31,94,31,114,31,241,31,56,31,56,30,56,29,56,28,152,31,231,31,78,31,40,31,120,31,120,30,120,29,120,28,143,31,143,30,42,31,63,31,36,31,70,31,102,31,154,31,83,31,137,31,242,31,196,31,48,31,16,31,78,31,78,30,220,31,162,31,162,30,166,31,224,31,253,31,220,31,36,31,157,31,155,31,182,31,182,30,182,29,76,31,135,31,195,31,2,31,2,30,244,31,58,31,96,31,157,31,157,30,157,29,147,31,147,30,147,29,147,28,252,31,236,31,251,31,251,30,117,31,117,30,82,31,13,31,189,31,68,31,230,31,230,30,58,31,159,31,159,30,55,31,55,30,55,29,178,31,208,31,208,30,194,31,103,31,101,31,24,31,24,30,148,31,99,31,81,31,176,31,5,31,59,31,217,31,114,31,14,31,205,31,36,31,159,31,98,31,73,31,90,31,232,31,24,31,192,31,1,31,134,31,135,31,96,31,144,31,243,31,2,31,176,31,176,30,235,31,203,31,252,31,13,31,13,30,13,29,71,31,159,31,205,31,63,31,230,31,154,31,235,31,140,31,221,31,238,31,238,30,101,31,234,31,234,30,23,31,114,31,32,31,218,31,218,30,218,29,223,31,105,31,4,31,31,31,54,31,123,31,123,30,178,31,178,30,105,31,68,31,40,31,2,31,32,31,53,31,2,31,18,31,134,31,183,31,54,31,54,30,234,31,108,31,172,31,47,31,228,31,177,31,24,31,127,31,176,31,176,30,176,29,21,31,142,31,43,31,153,31,153,30,153,29,176,31,70,31,193,31,193,30,225,31,237,31,236,31,213,31,125,31,178,31,120,31,250,31,219,31,62,31,228,31,12,31,35,31,29,31,89,31,186,31,28,31,28,30,28,29,34,31,29,31,45,31,93,31,96,31,23,31,29,31,248,31,248,30,248,29,229,31,168,31,168,30,165,31,165,30,206,31,245,31,229,31,114,31,87,31,11,31,11,30,1,31,66,31,196,31,87,31,87,30,114,31,185,31,161,31,243,31,120,31,74,31,217,31,72,31,14,31,156,31,64,31,147,31,107,31,241,31,83,31,233,31,73,31,114,31,54,31,49,31,183,31,185,31,29,31,115,31,23,31,181,31,161,31,71,31,166,31,31,31,31,30,31,29,73,31,73,30,73,29,34,31,128,31,28,31,28,30,124,31,124,30,143,31,7,31,170,31,170,30,170,29,170,28,238,31,76,31,166,31,155,31,187,31,113,31,113,30,94,31,43,31,40,31,204,31,59,31,59,30,59,29,59,28,169,31,122,31,122,30,122,29,103,31,88,31,50,31,52,31,211,31,218,31,248,31,42,31,42,30,8,31,1,31,111,31,206,31,29,31,95,31,95,31,155,31,242,31,252,31,88,31,208,31,62,31,211,31,211,30,209,31,32,31,120,31,231,31,117,31,79,31,63,31,137,31,35,31,57,31,157,31,214,31,185,31,104,31,5,31,5,30,107,31,60,31,60,30,68,31,53,31,149,31,51,31,50,31,155,31,65,31,108,31,253,31,117,31,197,31,197,30,197,29,197,28,125,31,206,31,181,31,184,31,98,31,174,31,174,30,101,31,72,31,72,30,81,31,251,31,251,30,13,31,13,30,238,31,29,31,178,31,181,31,32,31,32,31,12,31,12,30,161,31,197,31,197,30,176,31,183,31,66,31,79,31,153,31,153,30,228,31,219,31,116,31,116,30,55,31,55,30,74,31,44,31,138,31,40,31,192,31,112,31,162,31,207,31,196,31,190,31,72,31,128,31,34,31,43,31,43,30,43,29,16,31,16,30,19,31,129,31,241,31,167,31,121,31,179,31,250,31,6,31,87,31,87,30,114,31,8,31,63,31,115,31,23,31,55,31,205,31,205,30,200,31,74,31,74,30,74,29,212,31,55,31,118,31,118,30,118,29,118,28,158,31,156,31,201,31,91,31,91,30,138,31,5,31,97,31,41,31,144,31,144,30,200,31,231,31,160,31,160,30,136,31,136,30,199,31,67,31,67,30,154,31,202,31,202,30,92,31,54,31,105,31,112,31,179,31,55,31,55,30,41,31,41,30,87,31,198,31,6,31,252,31,252,30,252,29,71,31,110,31,113,31,86,31,86,30,45,31,146,31,146,30,190,31,24,31,24,30,83,31,14,31,123,31,123,31,123,30,239,31,3,31,3,30,122,31,228,31,176,31,15,31,239,31,239,30,151,31,18,31,64,31,64,30,117,31,19,31,186,31,204,31,54,31,183,31,183,30,183,29,151,31,7,31,135,31,102,31,72,31,182,31,69,31,69,30,184,31,110,31,110,30,6,31,126,31,224,31,224,30,222,31,50,31,50,30,50,29,61,31,139,31,139,30,72,31,223,31,119,31,44,31,130,31,218,31,82,31,4,31,4,30,4,29,71,31,116,31,81,31,15,31,188,31,170,31,170,30,62,31,47,31,21,31,21,30,160,31,220,31,222,31,222,30,107,31,235,31,109,31,85,31,85,30,161,31,11,31,193,31,219,31,223,31,138,31,105,31,156,31,178,31,136,31,138,31,36,31,45,31,45,30,45,29,66,31,91,31,91,30,230,31,230,30,230,29,71,31,95,31,105,31,66,31,91,31,207,31,205,31,205,30,205,29,109,31,27,31,142,31,96,31,96,30,111,31,132,31,132,30,229,31,240,31,253,31,127,31,223,31,164,31,164,30,164,29,164,28,164,27,228,31,132,31,201,31,211,31,58,31,4,31,4,30,4,29,71,31,40,31,40,30,162,31,175,31,175,30,175,29,88,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
