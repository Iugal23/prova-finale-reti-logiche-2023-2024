-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 380;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (129,0,213,0,0,0,210,0,89,0,149,0,102,0,251,0,208,0,234,0,0,0,198,0,0,0,104,0,0,0,152,0,0,0,231,0,193,0,219,0,0,0,108,0,230,0,136,0,0,0,19,0,0,0,212,0,33,0,103,0,135,0,13,0,16,0,0,0,253,0,83,0,218,0,253,0,67,0,212,0,0,0,235,0,142,0,10,0,119,0,85,0,98,0,12,0,137,0,79,0,214,0,0,0,81,0,88,0,222,0,249,0,220,0,26,0,0,0,20,0,73,0,0,0,31,0,58,0,0,0,101,0,0,0,238,0,223,0,216,0,151,0,183,0,120,0,185,0,3,0,25,0,8,0,181,0,0,0,172,0,0,0,68,0,155,0,170,0,202,0,0,0,0,0,48,0,90,0,0,0,0,0,243,0,213,0,134,0,0,0,90,0,204,0,151,0,0,0,217,0,0,0,123,0,248,0,0,0,97,0,183,0,131,0,14,0,130,0,120,0,243,0,150,0,0,0,29,0,99,0,0,0,28,0,131,0,241,0,180,0,204,0,107,0,60,0,178,0,118,0,189,0,0,0,149,0,185,0,195,0,78,0,164,0,0,0,0,0,14,0,77,0,211,0,104,0,14,0,92,0,15,0,80,0,21,0,168,0,25,0,87,0,0,0,228,0,90,0,62,0,100,0,191,0,89,0,207,0,27,0,0,0,130,0,161,0,55,0,224,0,186,0,0,0,223,0,79,0,214,0,148,0,55,0,100,0,0,0,0,0,12,0,174,0,0,0,102,0,18,0,100,0,6,0,31,0,16,0,57,0,0,0,112,0,88,0,104,0,0,0,0,0,23,0,122,0,154,0,0,0,176,0,184,0,126,0,127,0,0,0,77,0,132,0,0,0,0,0,192,0,250,0,83,0,225,0,74,0,17,0,0,0,11,0,149,0,80,0,0,0,0,0,0,0,86,0,15,0,194,0,149,0,153,0,63,0,0,0,74,0,0,0,42,0,0,0,80,0,221,0,190,0,182,0,228,0,45,0,223,0,115,0,71,0,0,0,234,0,30,0,134,0,55,0,168,0,211,0,36,0,29,0,84,0,210,0,146,0,36,0,238,0,0,0,0,0,28,0,208,0,156,0,1,0,23,0,77,0,0,0,219,0,153,0,28,0,95,0,26,0,223,0,63,0,0,0,54,0,129,0,160,0,8,0,26,0,151,0,0,0,0,0,70,0,39,0,0,0,206,0,38,0,0,0,63,0,0,0,0,0,0,0,120,0,68,0,105,0,0,0,45,0,29,0,135,0,17,0,0,0,0,0,0,0,238,0,173,0,117,0,252,0,134,0,109,0,105,0,39,0,15,0,152,0,226,0,0,0,0,0,0,0,0,0,235,0,178,0,243,0,251,0,134,0,10,0,0,0,182,0,28,0,36,0,101,0,25,0,78,0,0,0,0,0,4,0,236,0,94,0,153,0,65,0,0,0,232,0,20,0,0,0,198,0,205,0,0,0,134,0,185,0,27,0,0,0,0,0,51,0,78,0,172,0,182,0,0,0,140,0,28,0,137,0,0,0,239,0,101,0,0,0,0,0,22,0,188,0,220,0,0,0,120,0,82,0,234,0,116,0,0,0,37,0,255,0,165,0,139,0,235,0,0,0,126,0,180,0,0,0,248,0,80,0,126,0,136,0,226,0,141,0,0,0,121,0,0,0,0,0);
signal scenario_full  : scenario_type := (129,31,213,31,213,30,210,31,89,31,149,31,102,31,251,31,208,31,234,31,234,30,198,31,198,30,104,31,104,30,152,31,152,30,231,31,193,31,219,31,219,30,108,31,230,31,136,31,136,30,19,31,19,30,212,31,33,31,103,31,135,31,13,31,16,31,16,30,253,31,83,31,218,31,253,31,67,31,212,31,212,30,235,31,142,31,10,31,119,31,85,31,98,31,12,31,137,31,79,31,214,31,214,30,81,31,88,31,222,31,249,31,220,31,26,31,26,30,20,31,73,31,73,30,31,31,58,31,58,30,101,31,101,30,238,31,223,31,216,31,151,31,183,31,120,31,185,31,3,31,25,31,8,31,181,31,181,30,172,31,172,30,68,31,155,31,170,31,202,31,202,30,202,29,48,31,90,31,90,30,90,29,243,31,213,31,134,31,134,30,90,31,204,31,151,31,151,30,217,31,217,30,123,31,248,31,248,30,97,31,183,31,131,31,14,31,130,31,120,31,243,31,150,31,150,30,29,31,99,31,99,30,28,31,131,31,241,31,180,31,204,31,107,31,60,31,178,31,118,31,189,31,189,30,149,31,185,31,195,31,78,31,164,31,164,30,164,29,14,31,77,31,211,31,104,31,14,31,92,31,15,31,80,31,21,31,168,31,25,31,87,31,87,30,228,31,90,31,62,31,100,31,191,31,89,31,207,31,27,31,27,30,130,31,161,31,55,31,224,31,186,31,186,30,223,31,79,31,214,31,148,31,55,31,100,31,100,30,100,29,12,31,174,31,174,30,102,31,18,31,100,31,6,31,31,31,16,31,57,31,57,30,112,31,88,31,104,31,104,30,104,29,23,31,122,31,154,31,154,30,176,31,184,31,126,31,127,31,127,30,77,31,132,31,132,30,132,29,192,31,250,31,83,31,225,31,74,31,17,31,17,30,11,31,149,31,80,31,80,30,80,29,80,28,86,31,15,31,194,31,149,31,153,31,63,31,63,30,74,31,74,30,42,31,42,30,80,31,221,31,190,31,182,31,228,31,45,31,223,31,115,31,71,31,71,30,234,31,30,31,134,31,55,31,168,31,211,31,36,31,29,31,84,31,210,31,146,31,36,31,238,31,238,30,238,29,28,31,208,31,156,31,1,31,23,31,77,31,77,30,219,31,153,31,28,31,95,31,26,31,223,31,63,31,63,30,54,31,129,31,160,31,8,31,26,31,151,31,151,30,151,29,70,31,39,31,39,30,206,31,38,31,38,30,63,31,63,30,63,29,63,28,120,31,68,31,105,31,105,30,45,31,29,31,135,31,17,31,17,30,17,29,17,28,238,31,173,31,117,31,252,31,134,31,109,31,105,31,39,31,15,31,152,31,226,31,226,30,226,29,226,28,226,27,235,31,178,31,243,31,251,31,134,31,10,31,10,30,182,31,28,31,36,31,101,31,25,31,78,31,78,30,78,29,4,31,236,31,94,31,153,31,65,31,65,30,232,31,20,31,20,30,198,31,205,31,205,30,134,31,185,31,27,31,27,30,27,29,51,31,78,31,172,31,182,31,182,30,140,31,28,31,137,31,137,30,239,31,101,31,101,30,101,29,22,31,188,31,220,31,220,30,120,31,82,31,234,31,116,31,116,30,37,31,255,31,165,31,139,31,235,31,235,30,126,31,180,31,180,30,248,31,80,31,126,31,136,31,226,31,141,31,141,30,121,31,121,30,121,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
