-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_406 is
end project_tb_406;

architecture project_tb_arch_406 of project_tb_406 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 341;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (28,0,245,0,0,0,170,0,220,0,147,0,165,0,137,0,130,0,203,0,0,0,233,0,164,0,51,0,236,0,103,0,62,0,254,0,0,0,224,0,146,0,44,0,137,0,92,0,144,0,0,0,50,0,200,0,107,0,0,0,198,0,1,0,164,0,62,0,70,0,173,0,219,0,66,0,0,0,3,0,241,0,0,0,0,0,60,0,0,0,0,0,92,0,0,0,12,0,213,0,108,0,36,0,211,0,212,0,168,0,68,0,0,0,69,0,209,0,79,0,61,0,140,0,26,0,60,0,203,0,105,0,137,0,141,0,42,0,82,0,72,0,222,0,22,0,161,0,84,0,0,0,110,0,42,0,100,0,203,0,164,0,95,0,73,0,42,0,0,0,102,0,96,0,16,0,178,0,181,0,139,0,247,0,158,0,168,0,166,0,202,0,19,0,6,0,62,0,56,0,42,0,59,0,0,0,0,0,192,0,254,0,222,0,206,0,254,0,66,0,80,0,115,0,141,0,13,0,44,0,250,0,179,0,1,0,166,0,233,0,61,0,0,0,187,0,52,0,89,0,88,0,241,0,192,0,0,0,204,0,1,0,162,0,224,0,237,0,0,0,223,0,148,0,128,0,0,0,202,0,0,0,156,0,0,0,57,0,101,0,87,0,45,0,58,0,236,0,0,0,183,0,124,0,33,0,0,0,2,0,75,0,24,0,203,0,191,0,178,0,53,0,0,0,70,0,0,0,227,0,232,0,0,0,0,0,114,0,160,0,137,0,15,0,131,0,146,0,0,0,71,0,198,0,0,0,157,0,72,0,144,0,0,0,224,0,0,0,150,0,56,0,75,0,51,0,185,0,0,0,85,0,176,0,0,0,226,0,20,0,0,0,133,0,108,0,160,0,39,0,200,0,43,0,53,0,245,0,250,0,78,0,176,0,0,0,68,0,221,0,72,0,0,0,111,0,168,0,0,0,190,0,26,0,0,0,122,0,225,0,0,0,0,0,70,0,201,0,227,0,170,0,45,0,162,0,0,0,0,0,150,0,232,0,90,0,172,0,109,0,39,0,0,0,106,0,200,0,144,0,158,0,0,0,249,0,80,0,35,0,182,0,142,0,45,0,94,0,33,0,190,0,2,0,0,0,234,0,39,0,0,0,28,0,157,0,131,0,52,0,234,0,244,0,204,0,214,0,14,0,103,0,74,0,70,0,208,0,0,0,0,0,241,0,77,0,108,0,90,0,200,0,171,0,166,0,104,0,232,0,0,0,0,0,116,0,81,0,0,0,7,0,0,0,56,0,0,0,0,0,204,0,146,0,211,0,227,0,103,0,0,0,154,0,57,0,123,0,0,0,0,0,217,0,222,0,102,0,0,0,210,0,90,0,0,0,40,0,87,0,179,0,0,0,71,0,167,0,119,0,232,0,132,0,129,0,71,0,225,0,0,0,0,0,36,0,213,0,249,0,153,0,60,0,9,0,0,0,0,0,114,0,224,0,235,0,94,0,0,0,77,0,56,0,183,0,59,0,189,0,36,0);
signal scenario_full  : scenario_type := (28,31,245,31,245,30,170,31,220,31,147,31,165,31,137,31,130,31,203,31,203,30,233,31,164,31,51,31,236,31,103,31,62,31,254,31,254,30,224,31,146,31,44,31,137,31,92,31,144,31,144,30,50,31,200,31,107,31,107,30,198,31,1,31,164,31,62,31,70,31,173,31,219,31,66,31,66,30,3,31,241,31,241,30,241,29,60,31,60,30,60,29,92,31,92,30,12,31,213,31,108,31,36,31,211,31,212,31,168,31,68,31,68,30,69,31,209,31,79,31,61,31,140,31,26,31,60,31,203,31,105,31,137,31,141,31,42,31,82,31,72,31,222,31,22,31,161,31,84,31,84,30,110,31,42,31,100,31,203,31,164,31,95,31,73,31,42,31,42,30,102,31,96,31,16,31,178,31,181,31,139,31,247,31,158,31,168,31,166,31,202,31,19,31,6,31,62,31,56,31,42,31,59,31,59,30,59,29,192,31,254,31,222,31,206,31,254,31,66,31,80,31,115,31,141,31,13,31,44,31,250,31,179,31,1,31,166,31,233,31,61,31,61,30,187,31,52,31,89,31,88,31,241,31,192,31,192,30,204,31,1,31,162,31,224,31,237,31,237,30,223,31,148,31,128,31,128,30,202,31,202,30,156,31,156,30,57,31,101,31,87,31,45,31,58,31,236,31,236,30,183,31,124,31,33,31,33,30,2,31,75,31,24,31,203,31,191,31,178,31,53,31,53,30,70,31,70,30,227,31,232,31,232,30,232,29,114,31,160,31,137,31,15,31,131,31,146,31,146,30,71,31,198,31,198,30,157,31,72,31,144,31,144,30,224,31,224,30,150,31,56,31,75,31,51,31,185,31,185,30,85,31,176,31,176,30,226,31,20,31,20,30,133,31,108,31,160,31,39,31,200,31,43,31,53,31,245,31,250,31,78,31,176,31,176,30,68,31,221,31,72,31,72,30,111,31,168,31,168,30,190,31,26,31,26,30,122,31,225,31,225,30,225,29,70,31,201,31,227,31,170,31,45,31,162,31,162,30,162,29,150,31,232,31,90,31,172,31,109,31,39,31,39,30,106,31,200,31,144,31,158,31,158,30,249,31,80,31,35,31,182,31,142,31,45,31,94,31,33,31,190,31,2,31,2,30,234,31,39,31,39,30,28,31,157,31,131,31,52,31,234,31,244,31,204,31,214,31,14,31,103,31,74,31,70,31,208,31,208,30,208,29,241,31,77,31,108,31,90,31,200,31,171,31,166,31,104,31,232,31,232,30,232,29,116,31,81,31,81,30,7,31,7,30,56,31,56,30,56,29,204,31,146,31,211,31,227,31,103,31,103,30,154,31,57,31,123,31,123,30,123,29,217,31,222,31,102,31,102,30,210,31,90,31,90,30,40,31,87,31,179,31,179,30,71,31,167,31,119,31,232,31,132,31,129,31,71,31,225,31,225,30,225,29,36,31,213,31,249,31,153,31,60,31,9,31,9,30,9,29,114,31,224,31,235,31,94,31,94,30,77,31,56,31,183,31,59,31,189,31,36,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
