-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_771 is
end project_tb_771;

architecture project_tb_arch_771 of project_tb_771 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 664;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (185,0,74,0,244,0,0,0,21,0,29,0,0,0,190,0,17,0,160,0,197,0,38,0,7,0,148,0,106,0,120,0,130,0,0,0,112,0,161,0,134,0,0,0,245,0,105,0,72,0,32,0,0,0,0,0,0,0,107,0,93,0,0,0,103,0,244,0,61,0,45,0,0,0,68,0,150,0,81,0,134,0,0,0,129,0,0,0,0,0,111,0,0,0,0,0,33,0,249,0,0,0,174,0,0,0,110,0,0,0,87,0,55,0,189,0,157,0,230,0,0,0,27,0,0,0,46,0,221,0,0,0,14,0,220,0,57,0,25,0,0,0,0,0,10,0,210,0,95,0,67,0,111,0,45,0,92,0,241,0,218,0,56,0,190,0,246,0,0,0,64,0,187,0,242,0,80,0,147,0,162,0,186,0,38,0,72,0,147,0,0,0,164,0,116,0,214,0,0,0,39,0,0,0,222,0,0,0,179,0,0,0,117,0,174,0,8,0,0,0,249,0,41,0,52,0,51,0,154,0,244,0,37,0,129,0,174,0,244,0,108,0,217,0,94,0,52,0,122,0,249,0,113,0,94,0,60,0,36,0,142,0,0,0,254,0,166,0,0,0,0,0,249,0,0,0,0,0,212,0,195,0,212,0,65,0,9,0,0,0,113,0,53,0,4,0,195,0,0,0,218,0,135,0,86,0,27,0,255,0,173,0,91,0,132,0,159,0,157,0,127,0,115,0,217,0,107,0,151,0,0,0,126,0,121,0,106,0,241,0,70,0,92,0,0,0,73,0,195,0,192,0,251,0,22,0,9,0,74,0,226,0,0,0,238,0,0,0,98,0,63,0,0,0,105,0,0,0,217,0,178,0,52,0,47,0,0,0,41,0,115,0,0,0,226,0,127,0,120,0,211,0,236,0,0,0,127,0,81,0,97,0,0,0,0,0,133,0,66,0,0,0,40,0,0,0,200,0,124,0,9,0,0,0,2,0,0,0,114,0,0,0,89,0,247,0,136,0,1,0,93,0,226,0,35,0,75,0,0,0,105,0,77,0,0,0,0,0,102,0,121,0,85,0,127,0,0,0,207,0,0,0,0,0,0,0,0,0,0,0,57,0,13,0,107,0,0,0,0,0,201,0,0,0,170,0,115,0,0,0,166,0,158,0,33,0,127,0,97,0,166,0,40,0,0,0,0,0,6,0,11,0,11,0,85,0,80,0,235,0,102,0,74,0,65,0,11,0,225,0,156,0,140,0,125,0,0,0,128,0,19,0,235,0,51,0,172,0,27,0,0,0,76,0,90,0,108,0,79,0,0,0,0,0,204,0,152,0,166,0,42,0,12,0,123,0,0,0,48,0,199,0,0,0,229,0,0,0,0,0,101,0,187,0,27,0,90,0,185,0,73,0,81,0,214,0,0,0,36,0,11,0,35,0,195,0,177,0,72,0,230,0,109,0,0,0,52,0,228,0,174,0,98,0,6,0,174,0,0,0,223,0,224,0,137,0,0,0,71,0,251,0,246,0,174,0,202,0,140,0,224,0,244,0,149,0,0,0,253,0,245,0,0,0,164,0,0,0,254,0,180,0,191,0,213,0,83,0,177,0,185,0,238,0,1,0,215,0,201,0,0,0,0,0,68,0,102,0,0,0,220,0,0,0,235,0,144,0,0,0,137,0,0,0,223,0,240,0,35,0,67,0,8,0,160,0,198,0,139,0,186,0,151,0,184,0,185,0,0,0,79,0,175,0,0,0,16,0,179,0,132,0,125,0,247,0,108,0,11,0,32,0,199,0,65,0,146,0,114,0,196,0,0,0,143,0,239,0,54,0,104,0,9,0,29,0,85,0,114,0,170,0,92,0,238,0,220,0,221,0,98,0,153,0,0,0,71,0,126,0,36,0,148,0,216,0,73,0,0,0,195,0,174,0,125,0,217,0,61,0,0,0,76,0,203,0,59,0,156,0,144,0,0,0,142,0,62,0,233,0,187,0,128,0,0,0,0,0,43,0,186,0,91,0,0,0,0,0,110,0,243,0,16,0,233,0,88,0,50,0,34,0,103,0,102,0,218,0,89,0,17,0,99,0,197,0,139,0,114,0,0,0,0,0,122,0,124,0,139,0,65,0,181,0,8,0,0,0,55,0,59,0,116,0,248,0,1,0,198,0,0,0,125,0,147,0,105,0,180,0,0,0,162,0,77,0,239,0,239,0,4,0,0,0,0,0,146,0,155,0,0,0,0,0,124,0,0,0,57,0,77,0,171,0,8,0,222,0,134,0,250,0,31,0,188,0,102,0,71,0,80,0,160,0,31,0,0,0,42,0,59,0,0,0,233,0,23,0,240,0,112,0,58,0,97,0,168,0,24,0,149,0,83,0,0,0,38,0,48,0,244,0,129,0,112,0,199,0,126,0,241,0,25,0,0,0,121,0,71,0,119,0,64,0,0,0,189,0,47,0,138,0,0,0,180,0,48,0,0,0,37,0,24,0,0,0,89,0,187,0,149,0,142,0,180,0,244,0,0,0,154,0,183,0,10,0,77,0,249,0,0,0,169,0,0,0,45,0,81,0,232,0,87,0,0,0,0,0,134,0,0,0,188,0,4,0,7,0,79,0,77,0,0,0,84,0,205,0,0,0,233,0,207,0,50,0,238,0,0,0,116,0,137,0,208,0,0,0,0,0,14,0,78,0,158,0,25,0,127,0,239,0,175,0,239,0,53,0,152,0,110,0,227,0,0,0,25,0,0,0,179,0,149,0,39,0,86,0,238,0,0,0,132,0,98,0,252,0,48,0,77,0,0,0,248,0,228,0,0,0,167,0,21,0,184,0,29,0,7,0,0,0,111,0,0,0,237,0,122,0,137,0,89,0,238,0,0,0,0,0,55,0,83,0,102,0,0,0,138,0,9,0,0,0,0,0,0,0,119,0,236,0,76,0,78,0,192,0,39,0,153,0,160,0,0,0,0,0,207,0,249,0,1,0,0,0,0,0);
signal scenario_full  : scenario_type := (185,31,74,31,244,31,244,30,21,31,29,31,29,30,190,31,17,31,160,31,197,31,38,31,7,31,148,31,106,31,120,31,130,31,130,30,112,31,161,31,134,31,134,30,245,31,105,31,72,31,32,31,32,30,32,29,32,28,107,31,93,31,93,30,103,31,244,31,61,31,45,31,45,30,68,31,150,31,81,31,134,31,134,30,129,31,129,30,129,29,111,31,111,30,111,29,33,31,249,31,249,30,174,31,174,30,110,31,110,30,87,31,55,31,189,31,157,31,230,31,230,30,27,31,27,30,46,31,221,31,221,30,14,31,220,31,57,31,25,31,25,30,25,29,10,31,210,31,95,31,67,31,111,31,45,31,92,31,241,31,218,31,56,31,190,31,246,31,246,30,64,31,187,31,242,31,80,31,147,31,162,31,186,31,38,31,72,31,147,31,147,30,164,31,116,31,214,31,214,30,39,31,39,30,222,31,222,30,179,31,179,30,117,31,174,31,8,31,8,30,249,31,41,31,52,31,51,31,154,31,244,31,37,31,129,31,174,31,244,31,108,31,217,31,94,31,52,31,122,31,249,31,113,31,94,31,60,31,36,31,142,31,142,30,254,31,166,31,166,30,166,29,249,31,249,30,249,29,212,31,195,31,212,31,65,31,9,31,9,30,113,31,53,31,4,31,195,31,195,30,218,31,135,31,86,31,27,31,255,31,173,31,91,31,132,31,159,31,157,31,127,31,115,31,217,31,107,31,151,31,151,30,126,31,121,31,106,31,241,31,70,31,92,31,92,30,73,31,195,31,192,31,251,31,22,31,9,31,74,31,226,31,226,30,238,31,238,30,98,31,63,31,63,30,105,31,105,30,217,31,178,31,52,31,47,31,47,30,41,31,115,31,115,30,226,31,127,31,120,31,211,31,236,31,236,30,127,31,81,31,97,31,97,30,97,29,133,31,66,31,66,30,40,31,40,30,200,31,124,31,9,31,9,30,2,31,2,30,114,31,114,30,89,31,247,31,136,31,1,31,93,31,226,31,35,31,75,31,75,30,105,31,77,31,77,30,77,29,102,31,121,31,85,31,127,31,127,30,207,31,207,30,207,29,207,28,207,27,207,26,57,31,13,31,107,31,107,30,107,29,201,31,201,30,170,31,115,31,115,30,166,31,158,31,33,31,127,31,97,31,166,31,40,31,40,30,40,29,6,31,11,31,11,31,85,31,80,31,235,31,102,31,74,31,65,31,11,31,225,31,156,31,140,31,125,31,125,30,128,31,19,31,235,31,51,31,172,31,27,31,27,30,76,31,90,31,108,31,79,31,79,30,79,29,204,31,152,31,166,31,42,31,12,31,123,31,123,30,48,31,199,31,199,30,229,31,229,30,229,29,101,31,187,31,27,31,90,31,185,31,73,31,81,31,214,31,214,30,36,31,11,31,35,31,195,31,177,31,72,31,230,31,109,31,109,30,52,31,228,31,174,31,98,31,6,31,174,31,174,30,223,31,224,31,137,31,137,30,71,31,251,31,246,31,174,31,202,31,140,31,224,31,244,31,149,31,149,30,253,31,245,31,245,30,164,31,164,30,254,31,180,31,191,31,213,31,83,31,177,31,185,31,238,31,1,31,215,31,201,31,201,30,201,29,68,31,102,31,102,30,220,31,220,30,235,31,144,31,144,30,137,31,137,30,223,31,240,31,35,31,67,31,8,31,160,31,198,31,139,31,186,31,151,31,184,31,185,31,185,30,79,31,175,31,175,30,16,31,179,31,132,31,125,31,247,31,108,31,11,31,32,31,199,31,65,31,146,31,114,31,196,31,196,30,143,31,239,31,54,31,104,31,9,31,29,31,85,31,114,31,170,31,92,31,238,31,220,31,221,31,98,31,153,31,153,30,71,31,126,31,36,31,148,31,216,31,73,31,73,30,195,31,174,31,125,31,217,31,61,31,61,30,76,31,203,31,59,31,156,31,144,31,144,30,142,31,62,31,233,31,187,31,128,31,128,30,128,29,43,31,186,31,91,31,91,30,91,29,110,31,243,31,16,31,233,31,88,31,50,31,34,31,103,31,102,31,218,31,89,31,17,31,99,31,197,31,139,31,114,31,114,30,114,29,122,31,124,31,139,31,65,31,181,31,8,31,8,30,55,31,59,31,116,31,248,31,1,31,198,31,198,30,125,31,147,31,105,31,180,31,180,30,162,31,77,31,239,31,239,31,4,31,4,30,4,29,146,31,155,31,155,30,155,29,124,31,124,30,57,31,77,31,171,31,8,31,222,31,134,31,250,31,31,31,188,31,102,31,71,31,80,31,160,31,31,31,31,30,42,31,59,31,59,30,233,31,23,31,240,31,112,31,58,31,97,31,168,31,24,31,149,31,83,31,83,30,38,31,48,31,244,31,129,31,112,31,199,31,126,31,241,31,25,31,25,30,121,31,71,31,119,31,64,31,64,30,189,31,47,31,138,31,138,30,180,31,48,31,48,30,37,31,24,31,24,30,89,31,187,31,149,31,142,31,180,31,244,31,244,30,154,31,183,31,10,31,77,31,249,31,249,30,169,31,169,30,45,31,81,31,232,31,87,31,87,30,87,29,134,31,134,30,188,31,4,31,7,31,79,31,77,31,77,30,84,31,205,31,205,30,233,31,207,31,50,31,238,31,238,30,116,31,137,31,208,31,208,30,208,29,14,31,78,31,158,31,25,31,127,31,239,31,175,31,239,31,53,31,152,31,110,31,227,31,227,30,25,31,25,30,179,31,149,31,39,31,86,31,238,31,238,30,132,31,98,31,252,31,48,31,77,31,77,30,248,31,228,31,228,30,167,31,21,31,184,31,29,31,7,31,7,30,111,31,111,30,237,31,122,31,137,31,89,31,238,31,238,30,238,29,55,31,83,31,102,31,102,30,138,31,9,31,9,30,9,29,9,28,119,31,236,31,76,31,78,31,192,31,39,31,153,31,160,31,160,30,160,29,207,31,249,31,1,31,1,30,1,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
