-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_238 is
end project_tb_238;

architecture project_tb_arch_238 of project_tb_238 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 874;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (17,0,31,0,221,0,65,0,148,0,119,0,181,0,60,0,0,0,0,0,228,0,0,0,72,0,0,0,0,0,224,0,223,0,12,0,0,0,0,0,27,0,226,0,0,0,236,0,132,0,0,0,0,0,138,0,59,0,52,0,87,0,247,0,0,0,117,0,0,0,0,0,247,0,0,0,64,0,198,0,12,0,174,0,89,0,162,0,17,0,0,0,0,0,0,0,170,0,164,0,0,0,193,0,126,0,5,0,194,0,19,0,0,0,114,0,0,0,122,0,245,0,99,0,50,0,8,0,113,0,21,0,58,0,149,0,0,0,9,0,175,0,216,0,31,0,166,0,167,0,134,0,39,0,0,0,151,0,119,0,184,0,0,0,0,0,102,0,219,0,221,0,139,0,228,0,212,0,233,0,100,0,0,0,72,0,0,0,184,0,164,0,200,0,230,0,137,0,0,0,251,0,21,0,36,0,237,0,0,0,163,0,53,0,88,0,0,0,0,0,225,0,42,0,86,0,0,0,0,0,0,0,145,0,73,0,25,0,180,0,87,0,232,0,104,0,204,0,53,0,233,0,121,0,62,0,0,0,19,0,173,0,179,0,185,0,0,0,230,0,80,0,39,0,27,0,119,0,46,0,69,0,156,0,205,0,0,0,33,0,228,0,32,0,103,0,214,0,0,0,127,0,49,0,247,0,194,0,211,0,251,0,138,0,0,0,159,0,146,0,213,0,0,0,0,0,8,0,242,0,29,0,235,0,0,0,101,0,177,0,120,0,34,0,212,0,98,0,174,0,202,0,90,0,241,0,13,0,20,0,35,0,0,0,233,0,223,0,202,0,201,0,77,0,28,0,0,0,11,0,36,0,87,0,225,0,189,0,181,0,0,0,0,0,8,0,253,0,83,0,165,0,149,0,55,0,0,0,95,0,105,0,116,0,28,0,34,0,243,0,147,0,164,0,0,0,60,0,116,0,0,0,132,0,141,0,144,0,0,0,48,0,76,0,249,0,211,0,15,0,190,0,100,0,137,0,203,0,183,0,223,0,202,0,162,0,0,0,174,0,231,0,5,0,208,0,133,0,202,0,12,0,196,0,97,0,240,0,99,0,0,0,221,0,58,0,225,0,242,0,6,0,0,0,248,0,162,0,0,0,3,0,109,0,75,0,192,0,36,0,0,0,87,0,242,0,0,0,167,0,0,0,221,0,0,0,163,0,174,0,110,0,174,0,206,0,242,0,234,0,49,0,171,0,190,0,235,0,39,0,133,0,57,0,0,0,42,0,18,0,242,0,22,0,130,0,153,0,179,0,247,0,245,0,100,0,142,0,11,0,40,0,153,0,234,0,118,0,38,0,78,0,87,0,75,0,45,0,7,0,86,0,21,0,86,0,139,0,69,0,74,0,43,0,45,0,185,0,42,0,187,0,1,0,69,0,95,0,0,0,7,0,0,0,0,0,0,0,179,0,125,0,169,0,238,0,173,0,0,0,97,0,26,0,18,0,223,0,121,0,140,0,26,0,199,0,213,0,234,0,0,0,149,0,1,0,54,0,116,0,112,0,159,0,42,0,73,0,227,0,48,0,248,0,0,0,0,0,0,0,22,0,208,0,109,0,190,0,23,0,140,0,177,0,47,0,137,0,200,0,162,0,170,0,162,0,87,0,0,0,135,0,93,0,0,0,0,0,252,0,125,0,249,0,0,0,0,0,193,0,58,0,0,0,0,0,91,0,176,0,204,0,64,0,27,0,221,0,61,0,204,0,152,0,105,0,3,0,0,0,121,0,43,0,1,0,247,0,0,0,21,0,91,0,144,0,59,0,0,0,0,0,131,0,2,0,143,0,183,0,234,0,0,0,141,0,105,0,0,0,95,0,101,0,185,0,219,0,216,0,221,0,196,0,224,0,78,0,125,0,240,0,209,0,48,0,62,0,229,0,27,0,0,0,84,0,89,0,138,0,0,0,168,0,0,0,203,0,68,0,19,0,121,0,0,0,250,0,0,0,165,0,20,0,57,0,0,0,93,0,25,0,0,0,134,0,211,0,213,0,0,0,242,0,92,0,245,0,11,0,150,0,121,0,1,0,9,0,179,0,12,0,0,0,183,0,219,0,0,0,9,0,122,0,0,0,126,0,0,0,7,0,213,0,81,0,8,0,93,0,139,0,0,0,20,0,15,0,147,0,59,0,0,0,176,0,67,0,79,0,168,0,110,0,58,0,177,0,233,0,159,0,18,0,250,0,90,0,0,0,185,0,55,0,38,0,77,0,222,0,175,0,145,0,108,0,159,0,0,0,34,0,164,0,238,0,97,0,31,0,151,0,34,0,177,0,241,0,127,0,7,0,9,0,154,0,150,0,1,0,126,0,140,0,231,0,120,0,0,0,249,0,8,0,117,0,89,0,253,0,156,0,215,0,106,0,79,0,203,0,211,0,214,0,129,0,0,0,120,0,0,0,78,0,239,0,114,0,227,0,35,0,124,0,191,0,46,0,229,0,194,0,0,0,0,0,121,0,0,0,50,0,199,0,31,0,74,0,189,0,71,0,0,0,90,0,0,0,225,0,0,0,162,0,18,0,18,0,109,0,0,0,0,0,198,0,178,0,49,0,0,0,0,0,0,0,97,0,232,0,82,0,107,0,187,0,0,0,1,0,130,0,225,0,69,0,228,0,105,0,211,0,122,0,8,0,47,0,47,0,0,0,88,0,49,0,0,0,230,0,0,0,209,0,182,0,235,0,13,0,87,0,109,0,0,0,203,0,163,0,152,0,39,0,137,0,0,0,106,0,117,0,22,0,87,0,0,0,0,0,15,0,180,0,41,0,144,0,190,0,255,0,0,0,87,0,189,0,76,0,81,0,68,0,227,0,156,0,122,0,228,0,0,0,187,0,167,0,55,0,60,0,16,0,0,0,51,0,0,0,192,0,212,0,0,0,211,0,113,0,23,0,0,0,38,0,54,0,0,0,229,0,0,0,0,0,50,0,25,0,119,0,150,0,0,0,158,0,211,0,0,0,242,0,38,0,50,0,0,0,233,0,159,0,18,0,233,0,0,0,4,0,241,0,13,0,192,0,0,0,235,0,222,0,0,0,138,0,148,0,25,0,235,0,151,0,103,0,111,0,0,0,123,0,10,0,239,0,198,0,27,0,144,0,0,0,210,0,218,0,193,0,110,0,254,0,184,0,55,0,136,0,0,0,216,0,83,0,86,0,242,0,224,0,0,0,0,0,190,0,152,0,67,0,242,0,206,0,14,0,162,0,40,0,15,0,0,0,142,0,47,0,99,0,0,0,184,0,35,0,195,0,27,0,90,0,2,0,0,0,9,0,30,0,80,0,94,0,251,0,208,0,0,0,109,0,149,0,7,0,0,0,252,0,30,0,134,0,230,0,178,0,245,0,231,0,60,0,0,0,169,0,238,0,125,0,121,0,164,0,229,0,116,0,0,0,111,0,50,0,89,0,204,0,0,0,0,0,56,0,104,0,238,0,2,0,171,0,53,0,193,0,123,0,71,0,47,0,249,0,22,0,164,0,171,0,0,0,0,0,0,0,8,0,126,0,174,0,180,0,43,0,0,0,0,0,213,0,0,0,242,0,0,0,224,0,163,0,159,0,229,0,0,0,225,0,141,0,243,0,210,0,47,0,0,0,0,0,239,0,225,0,24,0,116,0,65,0,0,0,30,0,138,0,120,0,20,0,105,0,216,0,0,0,201,0,0,0,69,0,194,0,162,0,239,0,195,0,128,0,0,0,0,0,0,0,234,0,35,0,222,0,79,0,135,0,124,0,116,0,249,0,81,0,84,0,233,0,0,0,169,0,78,0,223,0,41,0,240,0,123,0,133,0,97,0,248,0,187,0,82,0,69,0,0,0,136,0,0,0,87,0,0,0,0,0,0,0,18,0,176,0,180,0,0,0,238,0);
signal scenario_full  : scenario_type := (17,31,31,31,221,31,65,31,148,31,119,31,181,31,60,31,60,30,60,29,228,31,228,30,72,31,72,30,72,29,224,31,223,31,12,31,12,30,12,29,27,31,226,31,226,30,236,31,132,31,132,30,132,29,138,31,59,31,52,31,87,31,247,31,247,30,117,31,117,30,117,29,247,31,247,30,64,31,198,31,12,31,174,31,89,31,162,31,17,31,17,30,17,29,17,28,170,31,164,31,164,30,193,31,126,31,5,31,194,31,19,31,19,30,114,31,114,30,122,31,245,31,99,31,50,31,8,31,113,31,21,31,58,31,149,31,149,30,9,31,175,31,216,31,31,31,166,31,167,31,134,31,39,31,39,30,151,31,119,31,184,31,184,30,184,29,102,31,219,31,221,31,139,31,228,31,212,31,233,31,100,31,100,30,72,31,72,30,184,31,164,31,200,31,230,31,137,31,137,30,251,31,21,31,36,31,237,31,237,30,163,31,53,31,88,31,88,30,88,29,225,31,42,31,86,31,86,30,86,29,86,28,145,31,73,31,25,31,180,31,87,31,232,31,104,31,204,31,53,31,233,31,121,31,62,31,62,30,19,31,173,31,179,31,185,31,185,30,230,31,80,31,39,31,27,31,119,31,46,31,69,31,156,31,205,31,205,30,33,31,228,31,32,31,103,31,214,31,214,30,127,31,49,31,247,31,194,31,211,31,251,31,138,31,138,30,159,31,146,31,213,31,213,30,213,29,8,31,242,31,29,31,235,31,235,30,101,31,177,31,120,31,34,31,212,31,98,31,174,31,202,31,90,31,241,31,13,31,20,31,35,31,35,30,233,31,223,31,202,31,201,31,77,31,28,31,28,30,11,31,36,31,87,31,225,31,189,31,181,31,181,30,181,29,8,31,253,31,83,31,165,31,149,31,55,31,55,30,95,31,105,31,116,31,28,31,34,31,243,31,147,31,164,31,164,30,60,31,116,31,116,30,132,31,141,31,144,31,144,30,48,31,76,31,249,31,211,31,15,31,190,31,100,31,137,31,203,31,183,31,223,31,202,31,162,31,162,30,174,31,231,31,5,31,208,31,133,31,202,31,12,31,196,31,97,31,240,31,99,31,99,30,221,31,58,31,225,31,242,31,6,31,6,30,248,31,162,31,162,30,3,31,109,31,75,31,192,31,36,31,36,30,87,31,242,31,242,30,167,31,167,30,221,31,221,30,163,31,174,31,110,31,174,31,206,31,242,31,234,31,49,31,171,31,190,31,235,31,39,31,133,31,57,31,57,30,42,31,18,31,242,31,22,31,130,31,153,31,179,31,247,31,245,31,100,31,142,31,11,31,40,31,153,31,234,31,118,31,38,31,78,31,87,31,75,31,45,31,7,31,86,31,21,31,86,31,139,31,69,31,74,31,43,31,45,31,185,31,42,31,187,31,1,31,69,31,95,31,95,30,7,31,7,30,7,29,7,28,179,31,125,31,169,31,238,31,173,31,173,30,97,31,26,31,18,31,223,31,121,31,140,31,26,31,199,31,213,31,234,31,234,30,149,31,1,31,54,31,116,31,112,31,159,31,42,31,73,31,227,31,48,31,248,31,248,30,248,29,248,28,22,31,208,31,109,31,190,31,23,31,140,31,177,31,47,31,137,31,200,31,162,31,170,31,162,31,87,31,87,30,135,31,93,31,93,30,93,29,252,31,125,31,249,31,249,30,249,29,193,31,58,31,58,30,58,29,91,31,176,31,204,31,64,31,27,31,221,31,61,31,204,31,152,31,105,31,3,31,3,30,121,31,43,31,1,31,247,31,247,30,21,31,91,31,144,31,59,31,59,30,59,29,131,31,2,31,143,31,183,31,234,31,234,30,141,31,105,31,105,30,95,31,101,31,185,31,219,31,216,31,221,31,196,31,224,31,78,31,125,31,240,31,209,31,48,31,62,31,229,31,27,31,27,30,84,31,89,31,138,31,138,30,168,31,168,30,203,31,68,31,19,31,121,31,121,30,250,31,250,30,165,31,20,31,57,31,57,30,93,31,25,31,25,30,134,31,211,31,213,31,213,30,242,31,92,31,245,31,11,31,150,31,121,31,1,31,9,31,179,31,12,31,12,30,183,31,219,31,219,30,9,31,122,31,122,30,126,31,126,30,7,31,213,31,81,31,8,31,93,31,139,31,139,30,20,31,15,31,147,31,59,31,59,30,176,31,67,31,79,31,168,31,110,31,58,31,177,31,233,31,159,31,18,31,250,31,90,31,90,30,185,31,55,31,38,31,77,31,222,31,175,31,145,31,108,31,159,31,159,30,34,31,164,31,238,31,97,31,31,31,151,31,34,31,177,31,241,31,127,31,7,31,9,31,154,31,150,31,1,31,126,31,140,31,231,31,120,31,120,30,249,31,8,31,117,31,89,31,253,31,156,31,215,31,106,31,79,31,203,31,211,31,214,31,129,31,129,30,120,31,120,30,78,31,239,31,114,31,227,31,35,31,124,31,191,31,46,31,229,31,194,31,194,30,194,29,121,31,121,30,50,31,199,31,31,31,74,31,189,31,71,31,71,30,90,31,90,30,225,31,225,30,162,31,18,31,18,31,109,31,109,30,109,29,198,31,178,31,49,31,49,30,49,29,49,28,97,31,232,31,82,31,107,31,187,31,187,30,1,31,130,31,225,31,69,31,228,31,105,31,211,31,122,31,8,31,47,31,47,31,47,30,88,31,49,31,49,30,230,31,230,30,209,31,182,31,235,31,13,31,87,31,109,31,109,30,203,31,163,31,152,31,39,31,137,31,137,30,106,31,117,31,22,31,87,31,87,30,87,29,15,31,180,31,41,31,144,31,190,31,255,31,255,30,87,31,189,31,76,31,81,31,68,31,227,31,156,31,122,31,228,31,228,30,187,31,167,31,55,31,60,31,16,31,16,30,51,31,51,30,192,31,212,31,212,30,211,31,113,31,23,31,23,30,38,31,54,31,54,30,229,31,229,30,229,29,50,31,25,31,119,31,150,31,150,30,158,31,211,31,211,30,242,31,38,31,50,31,50,30,233,31,159,31,18,31,233,31,233,30,4,31,241,31,13,31,192,31,192,30,235,31,222,31,222,30,138,31,148,31,25,31,235,31,151,31,103,31,111,31,111,30,123,31,10,31,239,31,198,31,27,31,144,31,144,30,210,31,218,31,193,31,110,31,254,31,184,31,55,31,136,31,136,30,216,31,83,31,86,31,242,31,224,31,224,30,224,29,190,31,152,31,67,31,242,31,206,31,14,31,162,31,40,31,15,31,15,30,142,31,47,31,99,31,99,30,184,31,35,31,195,31,27,31,90,31,2,31,2,30,9,31,30,31,80,31,94,31,251,31,208,31,208,30,109,31,149,31,7,31,7,30,252,31,30,31,134,31,230,31,178,31,245,31,231,31,60,31,60,30,169,31,238,31,125,31,121,31,164,31,229,31,116,31,116,30,111,31,50,31,89,31,204,31,204,30,204,29,56,31,104,31,238,31,2,31,171,31,53,31,193,31,123,31,71,31,47,31,249,31,22,31,164,31,171,31,171,30,171,29,171,28,8,31,126,31,174,31,180,31,43,31,43,30,43,29,213,31,213,30,242,31,242,30,224,31,163,31,159,31,229,31,229,30,225,31,141,31,243,31,210,31,47,31,47,30,47,29,239,31,225,31,24,31,116,31,65,31,65,30,30,31,138,31,120,31,20,31,105,31,216,31,216,30,201,31,201,30,69,31,194,31,162,31,239,31,195,31,128,31,128,30,128,29,128,28,234,31,35,31,222,31,79,31,135,31,124,31,116,31,249,31,81,31,84,31,233,31,233,30,169,31,78,31,223,31,41,31,240,31,123,31,133,31,97,31,248,31,187,31,82,31,69,31,69,30,136,31,136,30,87,31,87,30,87,29,87,28,18,31,176,31,180,31,180,30,238,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
