-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_321 is
end project_tb_321;

architecture project_tb_arch_321 of project_tb_321 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 739;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (251,0,12,0,228,0,83,0,180,0,80,0,251,0,72,0,0,0,0,0,153,0,181,0,0,0,133,0,172,0,209,0,30,0,245,0,164,0,0,0,207,0,205,0,38,0,0,0,147,0,71,0,148,0,0,0,76,0,31,0,0,0,121,0,89,0,153,0,17,0,35,0,0,0,115,0,0,0,101,0,0,0,68,0,123,0,0,0,156,0,39,0,153,0,148,0,0,0,226,0,239,0,186,0,42,0,176,0,191,0,229,0,138,0,87,0,162,0,0,0,138,0,233,0,140,0,0,0,161,0,142,0,0,0,0,0,248,0,45,0,254,0,0,0,210,0,107,0,182,0,35,0,76,0,72,0,83,0,16,0,0,0,128,0,71,0,89,0,0,0,144,0,71,0,0,0,233,0,192,0,142,0,5,0,153,0,111,0,206,0,82,0,130,0,226,0,0,0,16,0,0,0,7,0,58,0,0,0,17,0,139,0,0,0,50,0,202,0,220,0,105,0,0,0,98,0,10,0,122,0,75,0,97,0,27,0,199,0,154,0,153,0,5,0,92,0,237,0,0,0,244,0,103,0,160,0,193,0,84,0,32,0,36,0,76,0,160,0,20,0,0,0,250,0,68,0,0,0,137,0,24,0,84,0,64,0,0,0,106,0,0,0,170,0,0,0,0,0,0,0,83,0,0,0,77,0,7,0,145,0,0,0,112,0,0,0,215,0,96,0,0,0,64,0,27,0,0,0,42,0,237,0,144,0,240,0,249,0,202,0,123,0,161,0,175,0,31,0,147,0,71,0,254,0,96,0,65,0,193,0,0,0,165,0,7,0,98,0,23,0,219,0,122,0,120,0,25,0,210,0,75,0,0,0,197,0,183,0,2,0,2,0,87,0,147,0,189,0,78,0,245,0,157,0,0,0,223,0,51,0,104,0,0,0,235,0,0,0,227,0,219,0,0,0,126,0,93,0,201,0,0,0,130,0,0,0,235,0,163,0,147,0,68,0,0,0,0,0,83,0,172,0,130,0,40,0,131,0,150,0,71,0,0,0,240,0,58,0,72,0,0,0,0,0,111,0,250,0,125,0,96,0,6,0,162,0,87,0,0,0,150,0,3,0,145,0,176,0,114,0,203,0,0,0,65,0,150,0,119,0,0,0,237,0,75,0,90,0,193,0,116,0,0,0,33,0,221,0,28,0,104,0,115,0,97,0,145,0,166,0,26,0,47,0,0,0,111,0,1,0,236,0,58,0,0,0,0,0,176,0,94,0,180,0,189,0,205,0,169,0,0,0,1,0,245,0,49,0,241,0,224,0,141,0,2,0,101,0,226,0,234,0,122,0,0,0,194,0,167,0,128,0,250,0,0,0,76,0,163,0,11,0,203,0,0,0,111,0,229,0,43,0,123,0,77,0,159,0,0,0,240,0,31,0,208,0,182,0,103,0,0,0,0,0,132,0,109,0,37,0,51,0,204,0,238,0,209,0,0,0,242,0,225,0,147,0,41,0,101,0,226,0,0,0,51,0,140,0,159,0,40,0,109,0,0,0,31,0,0,0,0,0,74,0,254,0,61,0,238,0,83,0,0,0,70,0,163,0,0,0,170,0,143,0,106,0,0,0,164,0,115,0,180,0,53,0,15,0,249,0,250,0,75,0,235,0,174,0,0,0,41,0,0,0,0,0,135,0,0,0,93,0,213,0,94,0,116,0,0,0,191,0,167,0,56,0,215,0,196,0,191,0,251,0,29,0,235,0,0,0,160,0,39,0,0,0,14,0,195,0,231,0,153,0,87,0,87,0,190,0,112,0,0,0,16,0,238,0,199,0,246,0,255,0,3,0,15,0,109,0,30,0,82,0,186,0,0,0,118,0,156,0,160,0,12,0,86,0,16,0,146,0,214,0,51,0,9,0,223,0,231,0,234,0,200,0,0,0,212,0,71,0,0,0,167,0,88,0,232,0,49,0,0,0,223,0,43,0,33,0,80,0,0,0,126,0,0,0,36,0,111,0,41,0,41,0,161,0,0,0,0,0,201,0,253,0,179,0,93,0,0,0,155,0,0,0,227,0,0,0,112,0,226,0,0,0,155,0,192,0,197,0,195,0,31,0,5,0,140,0,162,0,38,0,0,0,127,0,159,0,58,0,144,0,0,0,46,0,43,0,6,0,81,0,93,0,0,0,163,0,0,0,93,0,129,0,229,0,0,0,139,0,94,0,120,0,15,0,198,0,59,0,141,0,183,0,10,0,61,0,0,0,206,0,87,0,204,0,0,0,54,0,153,0,243,0,0,0,62,0,174,0,0,0,6,0,108,0,0,0,0,0,0,0,218,0,0,0,51,0,192,0,207,0,4,0,0,0,150,0,123,0,111,0,53,0,216,0,37,0,67,0,78,0,153,0,0,0,6,0,24,0,68,0,0,0,238,0,104,0,93,0,189,0,237,0,222,0,207,0,36,0,107,0,106,0,0,0,29,0,87,0,0,0,67,0,112,0,0,0,117,0,45,0,54,0,174,0,74,0,131,0,128,0,235,0,186,0,54,0,128,0,0,0,175,0,118,0,138,0,42,0,226,0,29,0,212,0,191,0,240,0,78,0,128,0,6,0,0,0,230,0,112,0,0,0,169,0,119,0,246,0,10,0,13,0,166,0,89,0,205,0,85,0,245,0,100,0,227,0,241,0,169,0,234,0,219,0,161,0,158,0,0,0,67,0,200,0,134,0,128,0,7,0,252,0,0,0,9,0,154,0,74,0,109,0,0,0,239,0,217,0,204,0,0,0,75,0,58,0,221,0,131,0,231,0,0,0,111,0,0,0,145,0,227,0,9,0,138,0,31,0,253,0,179,0,161,0,0,0,20,0,168,0,41,0,179,0,180,0,207,0,186,0,0,0,0,0,55,0,145,0,243,0,133,0,67,0,236,0,244,0,87,0,164,0,90,0,87,0,37,0,32,0,202,0,118,0,33,0,0,0,0,0,0,0,80,0,94,0,193,0,32,0,136,0,114,0,129,0,68,0,0,0,120,0,1,0,233,0,0,0,4,0,0,0,142,0,142,0,38,0,85,0,235,0,155,0,17,0,0,0,0,0,0,0,237,0,0,0,0,0,0,0,225,0,209,0,173,0,100,0,133,0,243,0,229,0,132,0,9,0,78,0,69,0,0,0,101,0,41,0,218,0,244,0,163,0,0,0,29,0,161,0,220,0,0,0,38,0,0,0,41,0,180,0,179,0,8,0,0,0,73,0,118,0,191,0,204,0,187,0,105,0,110,0,0,0,74,0,36,0,31,0,0,0,110,0,0,0,41,0,0,0,182,0,10,0);
signal scenario_full  : scenario_type := (251,31,12,31,228,31,83,31,180,31,80,31,251,31,72,31,72,30,72,29,153,31,181,31,181,30,133,31,172,31,209,31,30,31,245,31,164,31,164,30,207,31,205,31,38,31,38,30,147,31,71,31,148,31,148,30,76,31,31,31,31,30,121,31,89,31,153,31,17,31,35,31,35,30,115,31,115,30,101,31,101,30,68,31,123,31,123,30,156,31,39,31,153,31,148,31,148,30,226,31,239,31,186,31,42,31,176,31,191,31,229,31,138,31,87,31,162,31,162,30,138,31,233,31,140,31,140,30,161,31,142,31,142,30,142,29,248,31,45,31,254,31,254,30,210,31,107,31,182,31,35,31,76,31,72,31,83,31,16,31,16,30,128,31,71,31,89,31,89,30,144,31,71,31,71,30,233,31,192,31,142,31,5,31,153,31,111,31,206,31,82,31,130,31,226,31,226,30,16,31,16,30,7,31,58,31,58,30,17,31,139,31,139,30,50,31,202,31,220,31,105,31,105,30,98,31,10,31,122,31,75,31,97,31,27,31,199,31,154,31,153,31,5,31,92,31,237,31,237,30,244,31,103,31,160,31,193,31,84,31,32,31,36,31,76,31,160,31,20,31,20,30,250,31,68,31,68,30,137,31,24,31,84,31,64,31,64,30,106,31,106,30,170,31,170,30,170,29,170,28,83,31,83,30,77,31,7,31,145,31,145,30,112,31,112,30,215,31,96,31,96,30,64,31,27,31,27,30,42,31,237,31,144,31,240,31,249,31,202,31,123,31,161,31,175,31,31,31,147,31,71,31,254,31,96,31,65,31,193,31,193,30,165,31,7,31,98,31,23,31,219,31,122,31,120,31,25,31,210,31,75,31,75,30,197,31,183,31,2,31,2,31,87,31,147,31,189,31,78,31,245,31,157,31,157,30,223,31,51,31,104,31,104,30,235,31,235,30,227,31,219,31,219,30,126,31,93,31,201,31,201,30,130,31,130,30,235,31,163,31,147,31,68,31,68,30,68,29,83,31,172,31,130,31,40,31,131,31,150,31,71,31,71,30,240,31,58,31,72,31,72,30,72,29,111,31,250,31,125,31,96,31,6,31,162,31,87,31,87,30,150,31,3,31,145,31,176,31,114,31,203,31,203,30,65,31,150,31,119,31,119,30,237,31,75,31,90,31,193,31,116,31,116,30,33,31,221,31,28,31,104,31,115,31,97,31,145,31,166,31,26,31,47,31,47,30,111,31,1,31,236,31,58,31,58,30,58,29,176,31,94,31,180,31,189,31,205,31,169,31,169,30,1,31,245,31,49,31,241,31,224,31,141,31,2,31,101,31,226,31,234,31,122,31,122,30,194,31,167,31,128,31,250,31,250,30,76,31,163,31,11,31,203,31,203,30,111,31,229,31,43,31,123,31,77,31,159,31,159,30,240,31,31,31,208,31,182,31,103,31,103,30,103,29,132,31,109,31,37,31,51,31,204,31,238,31,209,31,209,30,242,31,225,31,147,31,41,31,101,31,226,31,226,30,51,31,140,31,159,31,40,31,109,31,109,30,31,31,31,30,31,29,74,31,254,31,61,31,238,31,83,31,83,30,70,31,163,31,163,30,170,31,143,31,106,31,106,30,164,31,115,31,180,31,53,31,15,31,249,31,250,31,75,31,235,31,174,31,174,30,41,31,41,30,41,29,135,31,135,30,93,31,213,31,94,31,116,31,116,30,191,31,167,31,56,31,215,31,196,31,191,31,251,31,29,31,235,31,235,30,160,31,39,31,39,30,14,31,195,31,231,31,153,31,87,31,87,31,190,31,112,31,112,30,16,31,238,31,199,31,246,31,255,31,3,31,15,31,109,31,30,31,82,31,186,31,186,30,118,31,156,31,160,31,12,31,86,31,16,31,146,31,214,31,51,31,9,31,223,31,231,31,234,31,200,31,200,30,212,31,71,31,71,30,167,31,88,31,232,31,49,31,49,30,223,31,43,31,33,31,80,31,80,30,126,31,126,30,36,31,111,31,41,31,41,31,161,31,161,30,161,29,201,31,253,31,179,31,93,31,93,30,155,31,155,30,227,31,227,30,112,31,226,31,226,30,155,31,192,31,197,31,195,31,31,31,5,31,140,31,162,31,38,31,38,30,127,31,159,31,58,31,144,31,144,30,46,31,43,31,6,31,81,31,93,31,93,30,163,31,163,30,93,31,129,31,229,31,229,30,139,31,94,31,120,31,15,31,198,31,59,31,141,31,183,31,10,31,61,31,61,30,206,31,87,31,204,31,204,30,54,31,153,31,243,31,243,30,62,31,174,31,174,30,6,31,108,31,108,30,108,29,108,28,218,31,218,30,51,31,192,31,207,31,4,31,4,30,150,31,123,31,111,31,53,31,216,31,37,31,67,31,78,31,153,31,153,30,6,31,24,31,68,31,68,30,238,31,104,31,93,31,189,31,237,31,222,31,207,31,36,31,107,31,106,31,106,30,29,31,87,31,87,30,67,31,112,31,112,30,117,31,45,31,54,31,174,31,74,31,131,31,128,31,235,31,186,31,54,31,128,31,128,30,175,31,118,31,138,31,42,31,226,31,29,31,212,31,191,31,240,31,78,31,128,31,6,31,6,30,230,31,112,31,112,30,169,31,119,31,246,31,10,31,13,31,166,31,89,31,205,31,85,31,245,31,100,31,227,31,241,31,169,31,234,31,219,31,161,31,158,31,158,30,67,31,200,31,134,31,128,31,7,31,252,31,252,30,9,31,154,31,74,31,109,31,109,30,239,31,217,31,204,31,204,30,75,31,58,31,221,31,131,31,231,31,231,30,111,31,111,30,145,31,227,31,9,31,138,31,31,31,253,31,179,31,161,31,161,30,20,31,168,31,41,31,179,31,180,31,207,31,186,31,186,30,186,29,55,31,145,31,243,31,133,31,67,31,236,31,244,31,87,31,164,31,90,31,87,31,37,31,32,31,202,31,118,31,33,31,33,30,33,29,33,28,80,31,94,31,193,31,32,31,136,31,114,31,129,31,68,31,68,30,120,31,1,31,233,31,233,30,4,31,4,30,142,31,142,31,38,31,85,31,235,31,155,31,17,31,17,30,17,29,17,28,237,31,237,30,237,29,237,28,225,31,209,31,173,31,100,31,133,31,243,31,229,31,132,31,9,31,78,31,69,31,69,30,101,31,41,31,218,31,244,31,163,31,163,30,29,31,161,31,220,31,220,30,38,31,38,30,41,31,180,31,179,31,8,31,8,30,73,31,118,31,191,31,204,31,187,31,105,31,110,31,110,30,74,31,36,31,31,31,31,30,110,31,110,30,41,31,41,30,182,31,10,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
