-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_724 is
end project_tb_724;

architecture project_tb_arch_724 of project_tb_724 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1014;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (147,0,126,0,0,0,0,0,210,0,91,0,245,0,0,0,0,0,245,0,238,0,0,0,148,0,9,0,72,0,106,0,28,0,34,0,41,0,230,0,127,0,22,0,172,0,195,0,224,0,8,0,103,0,0,0,185,0,103,0,249,0,240,0,0,0,149,0,248,0,84,0,0,0,9,0,205,0,11,0,0,0,140,0,234,0,223,0,8,0,123,0,0,0,98,0,0,0,86,0,198,0,185,0,131,0,81,0,44,0,84,0,15,0,0,0,182,0,15,0,55,0,0,0,92,0,25,0,109,0,28,0,161,0,47,0,0,0,0,0,237,0,176,0,0,0,0,0,72,0,0,0,39,0,64,0,0,0,0,0,164,0,221,0,208,0,204,0,82,0,29,0,0,0,104,0,243,0,0,0,167,0,0,0,23,0,0,0,168,0,18,0,252,0,217,0,25,0,130,0,0,0,244,0,0,0,122,0,226,0,50,0,0,0,39,0,110,0,121,0,10,0,65,0,111,0,122,0,183,0,15,0,144,0,190,0,0,0,111,0,165,0,0,0,0,0,161,0,0,0,149,0,130,0,76,0,131,0,232,0,27,0,192,0,195,0,0,0,230,0,246,0,250,0,207,0,122,0,51,0,0,0,0,0,232,0,176,0,37,0,233,0,116,0,16,0,248,0,25,0,168,0,15,0,0,0,188,0,0,0,104,0,229,0,0,0,0,0,0,0,0,0,94,0,74,0,150,0,79,0,33,0,0,0,230,0,179,0,108,0,184,0,0,0,235,0,0,0,165,0,137,0,47,0,183,0,12,0,37,0,2,0,163,0,241,0,200,0,50,0,55,0,191,0,178,0,112,0,0,0,0,0,0,0,0,0,251,0,162,0,204,0,0,0,202,0,173,0,224,0,158,0,88,0,178,0,39,0,174,0,0,0,249,0,25,0,171,0,187,0,0,0,8,0,29,0,7,0,77,0,22,0,251,0,215,0,193,0,115,0,177,0,0,0,242,0,144,0,181,0,54,0,0,0,0,0,235,0,0,0,116,0,66,0,75,0,0,0,0,0,164,0,81,0,74,0,0,0,220,0,127,0,178,0,0,0,201,0,13,0,101,0,82,0,150,0,42,0,108,0,35,0,184,0,209,0,9,0,9,0,35,0,83,0,67,0,171,0,141,0,35,0,81,0,24,0,201,0,152,0,55,0,0,0,0,0,133,0,2,0,123,0,195,0,237,0,127,0,43,0,94,0,0,0,237,0,200,0,84,0,0,0,156,0,238,0,0,0,159,0,69,0,234,0,168,0,222,0,219,0,146,0,229,0,78,0,251,0,114,0,139,0,114,0,2,0,254,0,172,0,0,0,0,0,211,0,18,0,234,0,117,0,74,0,76,0,214,0,181,0,218,0,146,0,76,0,0,0,0,0,136,0,9,0,45,0,190,0,46,0,37,0,191,0,164,0,54,0,33,0,33,0,144,0,104,0,250,0,2,0,208,0,134,0,165,0,4,0,241,0,108,0,23,0,254,0,83,0,187,0,41,0,150,0,210,0,166,0,137,0,0,0,190,0,18,0,88,0,211,0,213,0,21,0,56,0,215,0,203,0,222,0,33,0,0,0,148,0,224,0,211,0,85,0,157,0,165,0,164,0,215,0,0,0,167,0,114,0,0,0,34,0,94,0,0,0,0,0,117,0,0,0,215,0,60,0,71,0,214,0,36,0,156,0,218,0,62,0,111,0,36,0,52,0,0,0,152,0,40,0,6,0,0,0,4,0,15,0,0,0,102,0,43,0,0,0,74,0,173,0,111,0,6,0,0,0,198,0,41,0,111,0,0,0,196,0,113,0,120,0,190,0,218,0,46,0,0,0,180,0,43,0,39,0,53,0,245,0,197,0,0,0,102,0,0,0,223,0,89,0,34,0,199,0,199,0,150,0,67,0,235,0,162,0,0,0,137,0,249,0,172,0,6,0,235,0,252,0,74,0,218,0,45,0,0,0,128,0,0,0,136,0,55,0,116,0,42,0,118,0,90,0,234,0,0,0,247,0,43,0,66,0,82,0,41,0,126,0,0,0,0,0,99,0,222,0,242,0,166,0,237,0,202,0,0,0,103,0,74,0,50,0,161,0,195,0,186,0,0,0,11,0,0,0,84,0,230,0,0,0,31,0,195,0,201,0,49,0,124,0,68,0,93,0,31,0,0,0,0,0,0,0,0,0,228,0,227,0,71,0,16,0,20,0,72,0,254,0,18,0,135,0,21,0,26,0,0,0,144,0,116,0,35,0,0,0,139,0,80,0,0,0,0,0,195,0,187,0,93,0,66,0,225,0,239,0,0,0,113,0,101,0,231,0,0,0,155,0,92,0,169,0,168,0,189,0,195,0,0,0,135,0,61,0,0,0,0,0,243,0,45,0,241,0,39,0,98,0,58,0,39,0,231,0,86,0,21,0,192,0,17,0,0,0,109,0,146,0,26,0,254,0,217,0,106,0,142,0,146,0,0,0,39,0,86,0,42,0,35,0,131,0,31,0,152,0,29,0,124,0,0,0,194,0,132,0,225,0,137,0,204,0,186,0,0,0,247,0,251,0,8,0,133,0,85,0,155,0,210,0,0,0,34,0,106,0,0,0,211,0,172,0,230,0,0,0,45,0,33,0,193,0,0,0,253,0,53,0,255,0,0,0,145,0,242,0,202,0,171,0,230,0,122,0,196,0,89,0,0,0,163,0,0,0,112,0,250,0,0,0,220,0,143,0,187,0,96,0,0,0,253,0,98,0,0,0,218,0,38,0,25,0,208,0,143,0,18,0,62,0,222,0,191,0,0,0,85,0,39,0,126,0,44,0,180,0,0,0,151,0,221,0,248,0,67,0,191,0,0,0,0,0,144,0,240,0,150,0,100,0,110,0,248,0,127,0,78,0,210,0,230,0,160,0,175,0,145,0,28,0,242,0,61,0,125,0,64,0,0,0,0,0,0,0,15,0,72,0,207,0,173,0,80,0,23,0,101,0,0,0,222,0,0,0,40,0,66,0,213,0,23,0,17,0,194,0,26,0,0,0,174,0,210,0,61,0,0,0,101,0,42,0,48,0,0,0,117,0,197,0,74,0,0,0,106,0,248,0,0,0,0,0,46,0,51,0,0,0,18,0,190,0,101,0,0,0,199,0,0,0,0,0,21,0,123,0,204,0,0,0,14,0,44,0,0,0,232,0,98,0,77,0,138,0,112,0,34,0,119,0,232,0,48,0,0,0,72,0,156,0,66,0,209,0,163,0,1,0,0,0,155,0,121,0,125,0,251,0,0,0,159,0,250,0,0,0,135,0,181,0,116,0,54,0,49,0,34,0,94,0,191,0,88,0,74,0,144,0,67,0,21,0,86,0,19,0,181,0,65,0,63,0,72,0,0,0,104,0,0,0,0,0,147,0,0,0,123,0,203,0,71,0,104,0,46,0,53,0,50,0,239,0,55,0,204,0,0,0,0,0,218,0,200,0,0,0,196,0,61,0,0,0,58,0,50,0,35,0,213,0,17,0,173,0,98,0,116,0,230,0,0,0,150,0,77,0,150,0,204,0,67,0,0,0,235,0,33,0,234,0,28,0,0,0,0,0,70,0,100,0,223,0,115,0,250,0,30,0,175,0,214,0,7,0,0,0,2,0,0,0,130,0,99,0,72,0,14,0,39,0,192,0,187,0,35,0,179,0,50,0,0,0,75,0,0,0,0,0,98,0,44,0,9,0,23,0,0,0,160,0,108,0,48,0,51,0,67,0,6,0,252,0,76,0,157,0,66,0,103,0,158,0,0,0,164,0,95,0,0,0,173,0,229,0,160,0,141,0,238,0,160,0,111,0,0,0,161,0,159,0,24,0,253,0,0,0,148,0,168,0,245,0,250,0,203,0,149,0,61,0,19,0,0,0,80,0,61,0,232,0,0,0,225,0,0,0,181,0,24,0,84,0,0,0,131,0,230,0,46,0,0,0,254,0,174,0,0,0,198,0,123,0,17,0,0,0,0,0,37,0,243,0,10,0,184,0,143,0,33,0,7,0,26,0,0,0,195,0,56,0,200,0,196,0,232,0,0,0,0,0,0,0,111,0,0,0,122,0,118,0,180,0,0,0,92,0,71,0,10,0,74,0,74,0,215,0,17,0,0,0,0,0,0,0,113,0,0,0,58,0,47,0,123,0,0,0,0,0,186,0,128,0,159,0,232,0,253,0,83,0,205,0,119,0,174,0,174,0,50,0,195,0,0,0,0,0,85,0,111,0,35,0,0,0,25,0,106,0,212,0,122,0,13,0,191,0,13,0,103,0,65,0,140,0,147,0,155,0,245,0,7,0,10,0,134,0,210,0,151,0,69,0,187,0,163,0,247,0,187,0,81,0,234,0,186,0,237,0,205,0,144,0,0,0,253,0,201,0,17,0,0,0,67,0,142,0,112,0,0,0,198,0,0,0,0,0,112,0,73,0,75,0,92,0,0,0,112,0,39,0,230,0,0,0,0,0,246,0,0,0,168,0,33,0,163,0,69,0,69,0,191,0,0,0,70,0,171,0);
signal scenario_full  : scenario_type := (147,31,126,31,126,30,126,29,210,31,91,31,245,31,245,30,245,29,245,31,238,31,238,30,148,31,9,31,72,31,106,31,28,31,34,31,41,31,230,31,127,31,22,31,172,31,195,31,224,31,8,31,103,31,103,30,185,31,103,31,249,31,240,31,240,30,149,31,248,31,84,31,84,30,9,31,205,31,11,31,11,30,140,31,234,31,223,31,8,31,123,31,123,30,98,31,98,30,86,31,198,31,185,31,131,31,81,31,44,31,84,31,15,31,15,30,182,31,15,31,55,31,55,30,92,31,25,31,109,31,28,31,161,31,47,31,47,30,47,29,237,31,176,31,176,30,176,29,72,31,72,30,39,31,64,31,64,30,64,29,164,31,221,31,208,31,204,31,82,31,29,31,29,30,104,31,243,31,243,30,167,31,167,30,23,31,23,30,168,31,18,31,252,31,217,31,25,31,130,31,130,30,244,31,244,30,122,31,226,31,50,31,50,30,39,31,110,31,121,31,10,31,65,31,111,31,122,31,183,31,15,31,144,31,190,31,190,30,111,31,165,31,165,30,165,29,161,31,161,30,149,31,130,31,76,31,131,31,232,31,27,31,192,31,195,31,195,30,230,31,246,31,250,31,207,31,122,31,51,31,51,30,51,29,232,31,176,31,37,31,233,31,116,31,16,31,248,31,25,31,168,31,15,31,15,30,188,31,188,30,104,31,229,31,229,30,229,29,229,28,229,27,94,31,74,31,150,31,79,31,33,31,33,30,230,31,179,31,108,31,184,31,184,30,235,31,235,30,165,31,137,31,47,31,183,31,12,31,37,31,2,31,163,31,241,31,200,31,50,31,55,31,191,31,178,31,112,31,112,30,112,29,112,28,112,27,251,31,162,31,204,31,204,30,202,31,173,31,224,31,158,31,88,31,178,31,39,31,174,31,174,30,249,31,25,31,171,31,187,31,187,30,8,31,29,31,7,31,77,31,22,31,251,31,215,31,193,31,115,31,177,31,177,30,242,31,144,31,181,31,54,31,54,30,54,29,235,31,235,30,116,31,66,31,75,31,75,30,75,29,164,31,81,31,74,31,74,30,220,31,127,31,178,31,178,30,201,31,13,31,101,31,82,31,150,31,42,31,108,31,35,31,184,31,209,31,9,31,9,31,35,31,83,31,67,31,171,31,141,31,35,31,81,31,24,31,201,31,152,31,55,31,55,30,55,29,133,31,2,31,123,31,195,31,237,31,127,31,43,31,94,31,94,30,237,31,200,31,84,31,84,30,156,31,238,31,238,30,159,31,69,31,234,31,168,31,222,31,219,31,146,31,229,31,78,31,251,31,114,31,139,31,114,31,2,31,254,31,172,31,172,30,172,29,211,31,18,31,234,31,117,31,74,31,76,31,214,31,181,31,218,31,146,31,76,31,76,30,76,29,136,31,9,31,45,31,190,31,46,31,37,31,191,31,164,31,54,31,33,31,33,31,144,31,104,31,250,31,2,31,208,31,134,31,165,31,4,31,241,31,108,31,23,31,254,31,83,31,187,31,41,31,150,31,210,31,166,31,137,31,137,30,190,31,18,31,88,31,211,31,213,31,21,31,56,31,215,31,203,31,222,31,33,31,33,30,148,31,224,31,211,31,85,31,157,31,165,31,164,31,215,31,215,30,167,31,114,31,114,30,34,31,94,31,94,30,94,29,117,31,117,30,215,31,60,31,71,31,214,31,36,31,156,31,218,31,62,31,111,31,36,31,52,31,52,30,152,31,40,31,6,31,6,30,4,31,15,31,15,30,102,31,43,31,43,30,74,31,173,31,111,31,6,31,6,30,198,31,41,31,111,31,111,30,196,31,113,31,120,31,190,31,218,31,46,31,46,30,180,31,43,31,39,31,53,31,245,31,197,31,197,30,102,31,102,30,223,31,89,31,34,31,199,31,199,31,150,31,67,31,235,31,162,31,162,30,137,31,249,31,172,31,6,31,235,31,252,31,74,31,218,31,45,31,45,30,128,31,128,30,136,31,55,31,116,31,42,31,118,31,90,31,234,31,234,30,247,31,43,31,66,31,82,31,41,31,126,31,126,30,126,29,99,31,222,31,242,31,166,31,237,31,202,31,202,30,103,31,74,31,50,31,161,31,195,31,186,31,186,30,11,31,11,30,84,31,230,31,230,30,31,31,195,31,201,31,49,31,124,31,68,31,93,31,31,31,31,30,31,29,31,28,31,27,228,31,227,31,71,31,16,31,20,31,72,31,254,31,18,31,135,31,21,31,26,31,26,30,144,31,116,31,35,31,35,30,139,31,80,31,80,30,80,29,195,31,187,31,93,31,66,31,225,31,239,31,239,30,113,31,101,31,231,31,231,30,155,31,92,31,169,31,168,31,189,31,195,31,195,30,135,31,61,31,61,30,61,29,243,31,45,31,241,31,39,31,98,31,58,31,39,31,231,31,86,31,21,31,192,31,17,31,17,30,109,31,146,31,26,31,254,31,217,31,106,31,142,31,146,31,146,30,39,31,86,31,42,31,35,31,131,31,31,31,152,31,29,31,124,31,124,30,194,31,132,31,225,31,137,31,204,31,186,31,186,30,247,31,251,31,8,31,133,31,85,31,155,31,210,31,210,30,34,31,106,31,106,30,211,31,172,31,230,31,230,30,45,31,33,31,193,31,193,30,253,31,53,31,255,31,255,30,145,31,242,31,202,31,171,31,230,31,122,31,196,31,89,31,89,30,163,31,163,30,112,31,250,31,250,30,220,31,143,31,187,31,96,31,96,30,253,31,98,31,98,30,218,31,38,31,25,31,208,31,143,31,18,31,62,31,222,31,191,31,191,30,85,31,39,31,126,31,44,31,180,31,180,30,151,31,221,31,248,31,67,31,191,31,191,30,191,29,144,31,240,31,150,31,100,31,110,31,248,31,127,31,78,31,210,31,230,31,160,31,175,31,145,31,28,31,242,31,61,31,125,31,64,31,64,30,64,29,64,28,15,31,72,31,207,31,173,31,80,31,23,31,101,31,101,30,222,31,222,30,40,31,66,31,213,31,23,31,17,31,194,31,26,31,26,30,174,31,210,31,61,31,61,30,101,31,42,31,48,31,48,30,117,31,197,31,74,31,74,30,106,31,248,31,248,30,248,29,46,31,51,31,51,30,18,31,190,31,101,31,101,30,199,31,199,30,199,29,21,31,123,31,204,31,204,30,14,31,44,31,44,30,232,31,98,31,77,31,138,31,112,31,34,31,119,31,232,31,48,31,48,30,72,31,156,31,66,31,209,31,163,31,1,31,1,30,155,31,121,31,125,31,251,31,251,30,159,31,250,31,250,30,135,31,181,31,116,31,54,31,49,31,34,31,94,31,191,31,88,31,74,31,144,31,67,31,21,31,86,31,19,31,181,31,65,31,63,31,72,31,72,30,104,31,104,30,104,29,147,31,147,30,123,31,203,31,71,31,104,31,46,31,53,31,50,31,239,31,55,31,204,31,204,30,204,29,218,31,200,31,200,30,196,31,61,31,61,30,58,31,50,31,35,31,213,31,17,31,173,31,98,31,116,31,230,31,230,30,150,31,77,31,150,31,204,31,67,31,67,30,235,31,33,31,234,31,28,31,28,30,28,29,70,31,100,31,223,31,115,31,250,31,30,31,175,31,214,31,7,31,7,30,2,31,2,30,130,31,99,31,72,31,14,31,39,31,192,31,187,31,35,31,179,31,50,31,50,30,75,31,75,30,75,29,98,31,44,31,9,31,23,31,23,30,160,31,108,31,48,31,51,31,67,31,6,31,252,31,76,31,157,31,66,31,103,31,158,31,158,30,164,31,95,31,95,30,173,31,229,31,160,31,141,31,238,31,160,31,111,31,111,30,161,31,159,31,24,31,253,31,253,30,148,31,168,31,245,31,250,31,203,31,149,31,61,31,19,31,19,30,80,31,61,31,232,31,232,30,225,31,225,30,181,31,24,31,84,31,84,30,131,31,230,31,46,31,46,30,254,31,174,31,174,30,198,31,123,31,17,31,17,30,17,29,37,31,243,31,10,31,184,31,143,31,33,31,7,31,26,31,26,30,195,31,56,31,200,31,196,31,232,31,232,30,232,29,232,28,111,31,111,30,122,31,118,31,180,31,180,30,92,31,71,31,10,31,74,31,74,31,215,31,17,31,17,30,17,29,17,28,113,31,113,30,58,31,47,31,123,31,123,30,123,29,186,31,128,31,159,31,232,31,253,31,83,31,205,31,119,31,174,31,174,31,50,31,195,31,195,30,195,29,85,31,111,31,35,31,35,30,25,31,106,31,212,31,122,31,13,31,191,31,13,31,103,31,65,31,140,31,147,31,155,31,245,31,7,31,10,31,134,31,210,31,151,31,69,31,187,31,163,31,247,31,187,31,81,31,234,31,186,31,237,31,205,31,144,31,144,30,253,31,201,31,17,31,17,30,67,31,142,31,112,31,112,30,198,31,198,30,198,29,112,31,73,31,75,31,92,31,92,30,112,31,39,31,230,31,230,30,230,29,246,31,246,30,168,31,33,31,163,31,69,31,69,31,191,31,191,30,70,31,171,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
