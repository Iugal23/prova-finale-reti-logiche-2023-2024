-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_84 is
end project_tb_84;

architecture project_tb_arch_84 of project_tb_84 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 898;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (26,0,81,0,160,0,169,0,176,0,0,0,44,0,254,0,0,0,87,0,19,0,16,0,131,0,10,0,53,0,96,0,0,0,146,0,150,0,163,0,43,0,0,0,209,0,133,0,73,0,116,0,211,0,209,0,189,0,0,0,241,0,218,0,115,0,134,0,12,0,31,0,0,0,39,0,31,0,0,0,94,0,119,0,14,0,104,0,107,0,251,0,152,0,255,0,163,0,97,0,131,0,132,0,199,0,23,0,245,0,52,0,0,0,234,0,104,0,80,0,210,0,137,0,190,0,181,0,140,0,144,0,114,0,12,0,167,0,0,0,144,0,105,0,0,0,62,0,152,0,0,0,202,0,240,0,184,0,111,0,163,0,42,0,0,0,83,0,44,0,2,0,44,0,53,0,24,0,198,0,224,0,185,0,0,0,124,0,9,0,54,0,228,0,113,0,135,0,91,0,253,0,0,0,110,0,156,0,8,0,0,0,0,0,18,0,202,0,0,0,40,0,119,0,88,0,218,0,0,0,0,0,0,0,0,0,124,0,0,0,0,0,145,0,0,0,121,0,24,0,174,0,0,0,16,0,182,0,115,0,255,0,94,0,0,0,120,0,0,0,197,0,16,0,128,0,232,0,78,0,133,0,43,0,113,0,0,0,194,0,7,0,117,0,233,0,100,0,0,0,112,0,151,0,0,0,232,0,0,0,66,0,129,0,102,0,230,0,81,0,210,0,249,0,0,0,110,0,0,0,68,0,0,0,231,0,93,0,252,0,0,0,0,0,244,0,210,0,0,0,100,0,181,0,172,0,11,0,144,0,1,0,235,0,0,0,247,0,172,0,205,0,213,0,130,0,65,0,26,0,0,0,216,0,116,0,100,0,158,0,0,0,0,0,214,0,0,0,0,0,0,0,0,0,0,0,138,0,0,0,67,0,166,0,158,0,74,0,252,0,0,0,188,0,109,0,0,0,50,0,45,0,226,0,0,0,0,0,199,0,170,0,138,0,243,0,246,0,150,0,201,0,86,0,27,0,85,0,135,0,56,0,112,0,109,0,181,0,40,0,0,0,131,0,162,0,237,0,174,0,121,0,100,0,186,0,97,0,0,0,102,0,0,0,102,0,45,0,122,0,11,0,224,0,0,0,62,0,195,0,153,0,228,0,77,0,0,0,0,0,0,0,72,0,0,0,210,0,206,0,55,0,0,0,102,0,149,0,28,0,94,0,157,0,224,0,0,0,234,0,0,0,93,0,113,0,201,0,60,0,212,0,0,0,137,0,6,0,111,0,0,0,53,0,250,0,87,0,77,0,149,0,243,0,120,0,125,0,230,0,0,0,23,0,217,0,0,0,226,0,149,0,103,0,0,0,49,0,45,0,69,0,246,0,175,0,0,0,0,0,190,0,236,0,91,0,118,0,0,0,0,0,111,0,118,0,128,0,244,0,127,0,91,0,90,0,0,0,125,0,114,0,165,0,243,0,0,0,31,0,80,0,122,0,33,0,42,0,108,0,54,0,83,0,235,0,46,0,127,0,219,0,0,0,0,0,2,0,45,0,0,0,13,0,234,0,0,0,59,0,0,0,54,0,114,0,119,0,0,0,0,0,58,0,188,0,88,0,9,0,223,0,48,0,114,0,181,0,184,0,195,0,182,0,134,0,48,0,144,0,206,0,188,0,211,0,227,0,245,0,144,0,208,0,108,0,148,0,158,0,226,0,18,0,116,0,0,0,128,0,203,0,0,0,175,0,157,0,0,0,235,0,160,0,20,0,218,0,168,0,249,0,138,0,0,0,227,0,0,0,133,0,172,0,168,0,48,0,240,0,79,0,0,0,255,0,226,0,209,0,165,0,145,0,51,0,191,0,216,0,10,0,44,0,44,0,52,0,130,0,137,0,7,0,191,0,114,0,0,0,172,0,192,0,240,0,96,0,187,0,60,0,0,0,0,0,115,0,228,0,176,0,154,0,86,0,133,0,185,0,41,0,80,0,0,0,104,0,0,0,104,0,28,0,224,0,48,0,0,0,187,0,88,0,56,0,162,0,88,0,207,0,69,0,16,0,130,0,0,0,254,0,228,0,0,0,206,0,142,0,94,0,120,0,218,0,0,0,248,0,151,0,234,0,209,0,80,0,213,0,0,0,213,0,79,0,118,0,162,0,124,0,179,0,244,0,79,0,83,0,127,0,161,0,155,0,3,0,0,0,0,0,79,0,76,0,0,0,190,0,154,0,161,0,159,0,0,0,211,0,106,0,38,0,118,0,0,0,162,0,22,0,0,0,251,0,45,0,0,0,254,0,5,0,0,0,9,0,0,0,0,0,10,0,27,0,205,0,146,0,124,0,131,0,246,0,105,0,82,0,89,0,121,0,2,0,157,0,200,0,91,0,186,0,232,0,0,0,49,0,246,0,104,0,81,0,66,0,245,0,198,0,0,0,224,0,245,0,0,0,182,0,2,0,82,0,9,0,10,0,142,0,201,0,131,0,112,0,0,0,255,0,202,0,189,0,245,0,133,0,241,0,121,0,208,0,0,0,168,0,58,0,17,0,83,0,151,0,113,0,100,0,19,0,236,0,231,0,166,0,8,0,115,0,233,0,99,0,92,0,0,0,0,0,0,0,168,0,0,0,0,0,245,0,224,0,5,0,195,0,254,0,185,0,77,0,174,0,29,0,16,0,143,0,189,0,42,0,52,0,19,0,57,0,198,0,86,0,181,0,172,0,22,0,0,0,61,0,106,0,154,0,0,0,0,0,43,0,105,0,162,0,170,0,58,0,0,0,94,0,232,0,129,0,64,0,57,0,242,0,35,0,224,0,0,0,219,0,0,0,161,0,57,0,250,0,238,0,198,0,0,0,28,0,0,0,0,0,237,0,206,0,0,0,56,0,0,0,71,0,0,0,0,0,11,0,165,0,230,0,90,0,16,0,174,0,25,0,0,0,34,0,245,0,0,0,77,0,184,0,138,0,0,0,45,0,227,0,238,0,41,0,0,0,248,0,3,0,117,0,226,0,3,0,144,0,0,0,74,0,172,0,194,0,0,0,22,0,214,0,86,0,10,0,35,0,89,0,160,0,83,0,229,0,49,0,26,0,97,0,19,0,0,0,61,0,163,0,41,0,191,0,102,0,235,0,27,0,173,0,173,0,180,0,0,0,63,0,149,0,106,0,109,0,164,0,32,0,167,0,165,0,113,0,92,0,230,0,75,0,83,0,241,0,0,0,173,0,148,0,0,0,0,0,145,0,43,0,114,0,108,0,0,0,37,0,33,0,137,0,143,0,0,0,230,0,179,0,209,0,232,0,209,0,5,0,12,0,0,0,26,0,146,0,237,0,0,0,56,0,243,0,58,0,157,0,59,0,185,0,235,0,162,0,29,0,181,0,212,0,0,0,90,0,108,0,90,0,235,0,0,0,0,0,197,0,0,0,78,0,217,0,116,0,133,0,0,0,219,0,111,0,189,0,0,0,76,0,38,0,64,0,0,0,143,0,214,0,219,0,104,0,0,0,180,0,58,0,0,0,251,0,142,0,180,0,0,0,21,0,154,0,189,0,242,0,106,0,47,0,0,0,0,0,131,0,61,0,0,0,0,0,140,0,243,0,0,0,139,0,50,0,111,0,237,0,112,0,200,0,166,0,229,0,138,0,0,0,226,0,200,0,187,0,164,0,0,0,34,0,203,0,18,0,252,0,0,0,115,0,12,0,124,0,0,0,209,0,40,0,0,0,150,0,25,0,206,0,176,0,49,0,143,0,186,0,0,0,42,0,138,0,0,0,255,0,94,0,216,0,112,0,213,0,163,0,171,0,253,0,166,0,202,0,56,0,0,0,127,0,11,0,165,0,101,0,132,0,201,0,0,0,86,0,0,0,90,0,138,0,54,0,23,0,132,0,167,0,209,0,8,0,65,0,162,0,199,0,0,0,97,0,0,0,0,0,114,0,119,0,0,0,0,0,85,0,153,0,141,0,25,0,224,0,0,0,150,0,127,0,247,0,202,0,1,0,0,0,224,0,141,0,227,0,0,0);
signal scenario_full  : scenario_type := (26,31,81,31,160,31,169,31,176,31,176,30,44,31,254,31,254,30,87,31,19,31,16,31,131,31,10,31,53,31,96,31,96,30,146,31,150,31,163,31,43,31,43,30,209,31,133,31,73,31,116,31,211,31,209,31,189,31,189,30,241,31,218,31,115,31,134,31,12,31,31,31,31,30,39,31,31,31,31,30,94,31,119,31,14,31,104,31,107,31,251,31,152,31,255,31,163,31,97,31,131,31,132,31,199,31,23,31,245,31,52,31,52,30,234,31,104,31,80,31,210,31,137,31,190,31,181,31,140,31,144,31,114,31,12,31,167,31,167,30,144,31,105,31,105,30,62,31,152,31,152,30,202,31,240,31,184,31,111,31,163,31,42,31,42,30,83,31,44,31,2,31,44,31,53,31,24,31,198,31,224,31,185,31,185,30,124,31,9,31,54,31,228,31,113,31,135,31,91,31,253,31,253,30,110,31,156,31,8,31,8,30,8,29,18,31,202,31,202,30,40,31,119,31,88,31,218,31,218,30,218,29,218,28,218,27,124,31,124,30,124,29,145,31,145,30,121,31,24,31,174,31,174,30,16,31,182,31,115,31,255,31,94,31,94,30,120,31,120,30,197,31,16,31,128,31,232,31,78,31,133,31,43,31,113,31,113,30,194,31,7,31,117,31,233,31,100,31,100,30,112,31,151,31,151,30,232,31,232,30,66,31,129,31,102,31,230,31,81,31,210,31,249,31,249,30,110,31,110,30,68,31,68,30,231,31,93,31,252,31,252,30,252,29,244,31,210,31,210,30,100,31,181,31,172,31,11,31,144,31,1,31,235,31,235,30,247,31,172,31,205,31,213,31,130,31,65,31,26,31,26,30,216,31,116,31,100,31,158,31,158,30,158,29,214,31,214,30,214,29,214,28,214,27,214,26,138,31,138,30,67,31,166,31,158,31,74,31,252,31,252,30,188,31,109,31,109,30,50,31,45,31,226,31,226,30,226,29,199,31,170,31,138,31,243,31,246,31,150,31,201,31,86,31,27,31,85,31,135,31,56,31,112,31,109,31,181,31,40,31,40,30,131,31,162,31,237,31,174,31,121,31,100,31,186,31,97,31,97,30,102,31,102,30,102,31,45,31,122,31,11,31,224,31,224,30,62,31,195,31,153,31,228,31,77,31,77,30,77,29,77,28,72,31,72,30,210,31,206,31,55,31,55,30,102,31,149,31,28,31,94,31,157,31,224,31,224,30,234,31,234,30,93,31,113,31,201,31,60,31,212,31,212,30,137,31,6,31,111,31,111,30,53,31,250,31,87,31,77,31,149,31,243,31,120,31,125,31,230,31,230,30,23,31,217,31,217,30,226,31,149,31,103,31,103,30,49,31,45,31,69,31,246,31,175,31,175,30,175,29,190,31,236,31,91,31,118,31,118,30,118,29,111,31,118,31,128,31,244,31,127,31,91,31,90,31,90,30,125,31,114,31,165,31,243,31,243,30,31,31,80,31,122,31,33,31,42,31,108,31,54,31,83,31,235,31,46,31,127,31,219,31,219,30,219,29,2,31,45,31,45,30,13,31,234,31,234,30,59,31,59,30,54,31,114,31,119,31,119,30,119,29,58,31,188,31,88,31,9,31,223,31,48,31,114,31,181,31,184,31,195,31,182,31,134,31,48,31,144,31,206,31,188,31,211,31,227,31,245,31,144,31,208,31,108,31,148,31,158,31,226,31,18,31,116,31,116,30,128,31,203,31,203,30,175,31,157,31,157,30,235,31,160,31,20,31,218,31,168,31,249,31,138,31,138,30,227,31,227,30,133,31,172,31,168,31,48,31,240,31,79,31,79,30,255,31,226,31,209,31,165,31,145,31,51,31,191,31,216,31,10,31,44,31,44,31,52,31,130,31,137,31,7,31,191,31,114,31,114,30,172,31,192,31,240,31,96,31,187,31,60,31,60,30,60,29,115,31,228,31,176,31,154,31,86,31,133,31,185,31,41,31,80,31,80,30,104,31,104,30,104,31,28,31,224,31,48,31,48,30,187,31,88,31,56,31,162,31,88,31,207,31,69,31,16,31,130,31,130,30,254,31,228,31,228,30,206,31,142,31,94,31,120,31,218,31,218,30,248,31,151,31,234,31,209,31,80,31,213,31,213,30,213,31,79,31,118,31,162,31,124,31,179,31,244,31,79,31,83,31,127,31,161,31,155,31,3,31,3,30,3,29,79,31,76,31,76,30,190,31,154,31,161,31,159,31,159,30,211,31,106,31,38,31,118,31,118,30,162,31,22,31,22,30,251,31,45,31,45,30,254,31,5,31,5,30,9,31,9,30,9,29,10,31,27,31,205,31,146,31,124,31,131,31,246,31,105,31,82,31,89,31,121,31,2,31,157,31,200,31,91,31,186,31,232,31,232,30,49,31,246,31,104,31,81,31,66,31,245,31,198,31,198,30,224,31,245,31,245,30,182,31,2,31,82,31,9,31,10,31,142,31,201,31,131,31,112,31,112,30,255,31,202,31,189,31,245,31,133,31,241,31,121,31,208,31,208,30,168,31,58,31,17,31,83,31,151,31,113,31,100,31,19,31,236,31,231,31,166,31,8,31,115,31,233,31,99,31,92,31,92,30,92,29,92,28,168,31,168,30,168,29,245,31,224,31,5,31,195,31,254,31,185,31,77,31,174,31,29,31,16,31,143,31,189,31,42,31,52,31,19,31,57,31,198,31,86,31,181,31,172,31,22,31,22,30,61,31,106,31,154,31,154,30,154,29,43,31,105,31,162,31,170,31,58,31,58,30,94,31,232,31,129,31,64,31,57,31,242,31,35,31,224,31,224,30,219,31,219,30,161,31,57,31,250,31,238,31,198,31,198,30,28,31,28,30,28,29,237,31,206,31,206,30,56,31,56,30,71,31,71,30,71,29,11,31,165,31,230,31,90,31,16,31,174,31,25,31,25,30,34,31,245,31,245,30,77,31,184,31,138,31,138,30,45,31,227,31,238,31,41,31,41,30,248,31,3,31,117,31,226,31,3,31,144,31,144,30,74,31,172,31,194,31,194,30,22,31,214,31,86,31,10,31,35,31,89,31,160,31,83,31,229,31,49,31,26,31,97,31,19,31,19,30,61,31,163,31,41,31,191,31,102,31,235,31,27,31,173,31,173,31,180,31,180,30,63,31,149,31,106,31,109,31,164,31,32,31,167,31,165,31,113,31,92,31,230,31,75,31,83,31,241,31,241,30,173,31,148,31,148,30,148,29,145,31,43,31,114,31,108,31,108,30,37,31,33,31,137,31,143,31,143,30,230,31,179,31,209,31,232,31,209,31,5,31,12,31,12,30,26,31,146,31,237,31,237,30,56,31,243,31,58,31,157,31,59,31,185,31,235,31,162,31,29,31,181,31,212,31,212,30,90,31,108,31,90,31,235,31,235,30,235,29,197,31,197,30,78,31,217,31,116,31,133,31,133,30,219,31,111,31,189,31,189,30,76,31,38,31,64,31,64,30,143,31,214,31,219,31,104,31,104,30,180,31,58,31,58,30,251,31,142,31,180,31,180,30,21,31,154,31,189,31,242,31,106,31,47,31,47,30,47,29,131,31,61,31,61,30,61,29,140,31,243,31,243,30,139,31,50,31,111,31,237,31,112,31,200,31,166,31,229,31,138,31,138,30,226,31,200,31,187,31,164,31,164,30,34,31,203,31,18,31,252,31,252,30,115,31,12,31,124,31,124,30,209,31,40,31,40,30,150,31,25,31,206,31,176,31,49,31,143,31,186,31,186,30,42,31,138,31,138,30,255,31,94,31,216,31,112,31,213,31,163,31,171,31,253,31,166,31,202,31,56,31,56,30,127,31,11,31,165,31,101,31,132,31,201,31,201,30,86,31,86,30,90,31,138,31,54,31,23,31,132,31,167,31,209,31,8,31,65,31,162,31,199,31,199,30,97,31,97,30,97,29,114,31,119,31,119,30,119,29,85,31,153,31,141,31,25,31,224,31,224,30,150,31,127,31,247,31,202,31,1,31,1,30,224,31,141,31,227,31,227,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
