-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 248;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (254,0,75,0,183,0,34,0,58,0,61,0,226,0,0,0,240,0,0,0,162,0,0,0,144,0,217,0,157,0,35,0,218,0,145,0,158,0,140,0,0,0,210,0,56,0,0,0,244,0,91,0,0,0,254,0,45,0,150,0,18,0,19,0,99,0,14,0,131,0,105,0,6,0,250,0,0,0,216,0,93,0,229,0,55,0,181,0,144,0,0,0,0,0,114,0,219,0,205,0,18,0,192,0,192,0,205,0,225,0,17,0,0,0,204,0,242,0,17,0,113,0,200,0,0,0,165,0,49,0,241,0,61,0,71,0,63,0,5,0,140,0,167,0,186,0,121,0,140,0,242,0,98,0,0,0,14,0,187,0,37,0,219,0,0,0,216,0,242,0,18,0,138,0,0,0,44,0,98,0,79,0,78,0,21,0,121,0,90,0,79,0,139,0,0,0,29,0,140,0,0,0,58,0,117,0,98,0,220,0,174,0,210,0,0,0,95,0,30,0,0,0,195,0,6,0,228,0,70,0,235,0,138,0,14,0,221,0,0,0,141,0,236,0,0,0,0,0,24,0,3,0,0,0,231,0,0,0,99,0,167,0,0,0,126,0,147,0,8,0,0,0,135,0,57,0,62,0,136,0,150,0,108,0,108,0,83,0,129,0,0,0,65,0,22,0,232,0,56,0,146,0,76,0,0,0,0,0,0,0,87,0,174,0,143,0,47,0,18,0,0,0,82,0,56,0,250,0,63,0,132,0,145,0,196,0,15,0,244,0,171,0,242,0,157,0,219,0,107,0,148,0,202,0,179,0,25,0,0,0,0,0,144,0,53,0,15,0,41,0,107,0,202,0,117,0,125,0,199,0,81,0,16,0,229,0,0,0,0,0,164,0,101,0,167,0,125,0,12,0,0,0,2,0,0,0,27,0,133,0,223,0,0,0,219,0,251,0,13,0,182,0,195,0,6,0,217,0,147,0,95,0,138,0,0,0,0,0,0,0,130,0,192,0,32,0,103,0,174,0,139,0,194,0,118,0,0,0,0,0,0,0,198,0,220,0,243,0,0,0,82,0,193,0,58,0,0,0,209,0,29,0,27,0,171,0,224,0,100,0,90,0,158,0,117,0);
signal scenario_full  : scenario_type := (254,31,75,31,183,31,34,31,58,31,61,31,226,31,226,30,240,31,240,30,162,31,162,30,144,31,217,31,157,31,35,31,218,31,145,31,158,31,140,31,140,30,210,31,56,31,56,30,244,31,91,31,91,30,254,31,45,31,150,31,18,31,19,31,99,31,14,31,131,31,105,31,6,31,250,31,250,30,216,31,93,31,229,31,55,31,181,31,144,31,144,30,144,29,114,31,219,31,205,31,18,31,192,31,192,31,205,31,225,31,17,31,17,30,204,31,242,31,17,31,113,31,200,31,200,30,165,31,49,31,241,31,61,31,71,31,63,31,5,31,140,31,167,31,186,31,121,31,140,31,242,31,98,31,98,30,14,31,187,31,37,31,219,31,219,30,216,31,242,31,18,31,138,31,138,30,44,31,98,31,79,31,78,31,21,31,121,31,90,31,79,31,139,31,139,30,29,31,140,31,140,30,58,31,117,31,98,31,220,31,174,31,210,31,210,30,95,31,30,31,30,30,195,31,6,31,228,31,70,31,235,31,138,31,14,31,221,31,221,30,141,31,236,31,236,30,236,29,24,31,3,31,3,30,231,31,231,30,99,31,167,31,167,30,126,31,147,31,8,31,8,30,135,31,57,31,62,31,136,31,150,31,108,31,108,31,83,31,129,31,129,30,65,31,22,31,232,31,56,31,146,31,76,31,76,30,76,29,76,28,87,31,174,31,143,31,47,31,18,31,18,30,82,31,56,31,250,31,63,31,132,31,145,31,196,31,15,31,244,31,171,31,242,31,157,31,219,31,107,31,148,31,202,31,179,31,25,31,25,30,25,29,144,31,53,31,15,31,41,31,107,31,202,31,117,31,125,31,199,31,81,31,16,31,229,31,229,30,229,29,164,31,101,31,167,31,125,31,12,31,12,30,2,31,2,30,27,31,133,31,223,31,223,30,219,31,251,31,13,31,182,31,195,31,6,31,217,31,147,31,95,31,138,31,138,30,138,29,138,28,130,31,192,31,32,31,103,31,174,31,139,31,194,31,118,31,118,30,118,29,118,28,198,31,220,31,243,31,243,30,82,31,193,31,58,31,58,30,209,31,29,31,27,31,171,31,224,31,100,31,90,31,158,31,117,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
