-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 980;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (83,0,0,0,0,0,154,0,97,0,0,0,0,0,233,0,0,0,43,0,14,0,44,0,153,0,96,0,61,0,0,0,0,0,109,0,9,0,191,0,56,0,39,0,72,0,235,0,176,0,251,0,22,0,9,0,130,0,5,0,0,0,133,0,215,0,247,0,104,0,211,0,240,0,243,0,247,0,50,0,103,0,251,0,0,0,0,0,0,0,44,0,255,0,0,0,0,0,66,0,208,0,40,0,168,0,86,0,78,0,204,0,182,0,40,0,0,0,0,0,30,0,0,0,145,0,70,0,141,0,170,0,0,0,73,0,126,0,170,0,0,0,0,0,249,0,169,0,0,0,191,0,88,0,145,0,229,0,17,0,249,0,0,0,235,0,233,0,0,0,20,0,0,0,98,0,37,0,165,0,7,0,45,0,205,0,129,0,56,0,106,0,196,0,168,0,0,0,121,0,92,0,0,0,0,0,7,0,0,0,84,0,88,0,169,0,16,0,114,0,230,0,128,0,11,0,50,0,0,0,229,0,0,0,1,0,129,0,157,0,25,0,38,0,0,0,165,0,200,0,45,0,23,0,50,0,0,0,0,0,14,0,218,0,0,0,43,0,0,0,247,0,15,0,0,0,0,0,198,0,26,0,0,0,182,0,230,0,0,0,201,0,0,0,0,0,0,0,229,0,39,0,234,0,206,0,0,0,0,0,193,0,45,0,0,0,232,0,216,0,26,0,247,0,52,0,11,0,1,0,0,0,77,0,242,0,106,0,9,0,140,0,0,0,244,0,74,0,77,0,11,0,249,0,126,0,156,0,121,0,104,0,140,0,19,0,90,0,130,0,239,0,63,0,218,0,190,0,223,0,0,0,151,0,237,0,0,0,253,0,90,0,7,0,237,0,72,0,121,0,118,0,251,0,141,0,173,0,76,0,201,0,93,0,193,0,207,0,154,0,239,0,80,0,0,0,0,0,209,0,39,0,231,0,231,0,0,0,238,0,189,0,111,0,25,0,200,0,0,0,98,0,0,0,68,0,187,0,4,0,245,0,20,0,205,0,28,0,90,0,112,0,61,0,212,0,75,0,132,0,252,0,83,0,97,0,6,0,0,0,220,0,241,0,26,0,17,0,148,0,40,0,49,0,0,0,67,0,89,0,209,0,150,0,182,0,210,0,126,0,75,0,215,0,194,0,93,0,93,0,66,0,0,0,133,0,132,0,189,0,0,0,230,0,230,0,198,0,250,0,0,0,0,0,0,0,184,0,65,0,0,0,168,0,175,0,0,0,254,0,0,0,195,0,6,0,253,0,26,0,155,0,0,0,239,0,229,0,0,0,197,0,0,0,75,0,27,0,0,0,235,0,101,0,0,0,18,0,141,0,89,0,0,0,239,0,0,0,96,0,0,0,243,0,0,0,128,0,94,0,118,0,53,0,3,0,0,0,45,0,157,0,207,0,162,0,0,0,129,0,180,0,178,0,0,0,0,0,214,0,41,0,43,0,208,0,201,0,127,0,26,0,134,0,202,0,21,0,0,0,225,0,187,0,99,0,20,0,244,0,226,0,0,0,253,0,60,0,202,0,148,0,0,0,0,0,103,0,238,0,58,0,138,0,111,0,52,0,181,0,39,0,109,0,250,0,49,0,86,0,0,0,104,0,248,0,62,0,203,0,214,0,91,0,252,0,177,0,223,0,151,0,224,0,108,0,96,0,172,0,137,0,0,0,45,0,186,0,71,0,0,0,252,0,44,0,3,0,231,0,203,0,229,0,223,0,0,0,125,0,0,0,135,0,102,0,0,0,37,0,239,0,54,0,176,0,0,0,212,0,46,0,216,0,0,0,168,0,0,0,0,0,0,0,17,0,31,0,113,0,48,0,0,0,87,0,217,0,182,0,29,0,184,0,20,0,180,0,88,0,24,0,112,0,97,0,187,0,209,0,109,0,0,0,0,0,0,0,195,0,202,0,70,0,57,0,156,0,0,0,153,0,135,0,0,0,171,0,94,0,232,0,146,0,48,0,89,0,228,0,72,0,0,0,61,0,70,0,8,0,178,0,56,0,206,0,10,0,91,0,147,0,0,0,40,0,78,0,23,0,33,0,0,0,0,0,5,0,67,0,63,0,48,0,80,0,25,0,149,0,112,0,109,0,155,0,75,0,95,0,94,0,94,0,51,0,7,0,68,0,56,0,0,0,0,0,0,0,0,0,118,0,247,0,168,0,15,0,117,0,208,0,24,0,211,0,195,0,0,0,24,0,0,0,222,0,0,0,0,0,222,0,57,0,207,0,0,0,183,0,84,0,0,0,177,0,61,0,76,0,101,0,184,0,42,0,55,0,0,0,20,0,134,0,0,0,243,0,2,0,103,0,87,0,161,0,0,0,134,0,188,0,12,0,42,0,203,0,251,0,51,0,53,0,0,0,0,0,0,0,178,0,0,0,249,0,124,0,0,0,80,0,40,0,41,0,206,0,90,0,0,0,0,0,32,0,0,0,131,0,154,0,58,0,69,0,144,0,117,0,161,0,0,0,0,0,122,0,6,0,52,0,199,0,0,0,20,0,225,0,0,0,117,0,16,0,97,0,0,0,190,0,133,0,198,0,11,0,0,0,93,0,68,0,149,0,21,0,92,0,212,0,0,0,0,0,185,0,227,0,45,0,0,0,144,0,218,0,80,0,147,0,8,0,125,0,44,0,206,0,179,0,112,0,32,0,81,0,101,0,240,0,0,0,76,0,14,0,160,0,164,0,0,0,25,0,58,0,22,0,0,0,0,0,177,0,70,0,130,0,0,0,12,0,46,0,211,0,0,0,56,0,0,0,81,0,159,0,148,0,0,0,173,0,90,0,202,0,160,0,146,0,0,0,83,0,186,0,135,0,169,0,161,0,105,0,88,0,9,0,199,0,89,0,172,0,236,0,231,0,247,0,102,0,171,0,78,0,202,0,15,0,220,0,108,0,53,0,0,0,42,0,223,0,0,0,104,0,57,0,216,0,0,0,94,0,93,0,35,0,10,0,5,0,242,0,44,0,151,0,17,0,41,0,0,0,13,0,0,0,89,0,233,0,87,0,0,0,90,0,0,0,132,0,129,0,231,0,144,0,36,0,255,0,0,0,129,0,125,0,122,0,0,0,23,0,101,0,25,0,0,0,87,0,250,0,151,0,205,0,147,0,184,0,152,0,0,0,37,0,67,0,190,0,109,0,140,0,48,0,38,0,228,0,251,0,0,0,204,0,41,0,0,0,198,0,48,0,50,0,47,0,145,0,0,0,27,0,246,0,97,0,197,0,0,0,43,0,211,0,81,0,245,0,0,0,26,0,248,0,176,0,73,0,193,0,62,0,150,0,125,0,196,0,227,0,4,0,86,0,238,0,175,0,44,0,210,0,122,0,0,0,68,0,0,0,39,0,60,0,0,0,151,0,181,0,142,0,8,0,35,0,120,0,195,0,190,0,0,0,66,0,51,0,46,0,182,0,223,0,188,0,82,0,34,0,29,0,115,0,169,0,0,0,0,0,143,0,174,0,131,0,21,0,111,0,0,0,108,0,230,0,0,0,23,0,79,0,86,0,0,0,7,0,9,0,1,0,60,0,209,0,148,0,0,0,62,0,73,0,65,0,0,0,53,0,0,0,44,0,203,0,129,0,22,0,213,0,50,0,40,0,51,0,67,0,0,0,236,0,196,0,37,0,150,0,1,0,254,0,219,0,0,0,0,0,69,0,173,0,43,0,236,0,74,0,0,0,20,0,113,0,0,0,0,0,47,0,131,0,110,0,113,0,67,0,0,0,0,0,186,0,26,0,87,0,213,0,0,0,61,0,84,0,78,0,172,0,240,0,202,0,79,0,0,0,72,0,69,0,107,0,0,0,202,0,0,0,0,0,124,0,0,0,247,0,0,0,143,0,27,0,205,0,198,0,78,0,0,0,241,0,245,0,245,0,0,0,83,0,0,0,41,0,89,0,0,0,21,0,153,0,130,0,0,0,210,0,57,0,152,0,226,0,70,0,214,0,0,0,0,0,217,0,169,0,9,0,147,0,80,0,170,0,56,0,64,0,3,0,187,0,16,0,21,0,8,0,80,0,0,0,11,0,0,0,215,0,107,0,194,0,162,0,0,0,1,0,139,0,23,0,0,0,0,0,30,0,197,0,18,0,28,0,60,0,21,0,90,0,155,0,79,0,104,0,202,0,0,0,200,0,254,0,97,0,6,0,0,0,114,0,183,0,162,0,0,0,234,0,23,0,212,0,96,0,90,0,0,0,100,0,194,0,82,0,138,0,94,0,2,0,143,0,251,0,32,0,34,0,0,0,108,0,12,0,8,0,8,0,109,0,97,0,44,0,18,0,214,0,217,0,38,0,116,0,0,0,0,0,0,0,0,0,33,0,133,0,48,0);
signal scenario_full  : scenario_type := (83,31,83,30,83,29,154,31,97,31,97,30,97,29,233,31,233,30,43,31,14,31,44,31,153,31,96,31,61,31,61,30,61,29,109,31,9,31,191,31,56,31,39,31,72,31,235,31,176,31,251,31,22,31,9,31,130,31,5,31,5,30,133,31,215,31,247,31,104,31,211,31,240,31,243,31,247,31,50,31,103,31,251,31,251,30,251,29,251,28,44,31,255,31,255,30,255,29,66,31,208,31,40,31,168,31,86,31,78,31,204,31,182,31,40,31,40,30,40,29,30,31,30,30,145,31,70,31,141,31,170,31,170,30,73,31,126,31,170,31,170,30,170,29,249,31,169,31,169,30,191,31,88,31,145,31,229,31,17,31,249,31,249,30,235,31,233,31,233,30,20,31,20,30,98,31,37,31,165,31,7,31,45,31,205,31,129,31,56,31,106,31,196,31,168,31,168,30,121,31,92,31,92,30,92,29,7,31,7,30,84,31,88,31,169,31,16,31,114,31,230,31,128,31,11,31,50,31,50,30,229,31,229,30,1,31,129,31,157,31,25,31,38,31,38,30,165,31,200,31,45,31,23,31,50,31,50,30,50,29,14,31,218,31,218,30,43,31,43,30,247,31,15,31,15,30,15,29,198,31,26,31,26,30,182,31,230,31,230,30,201,31,201,30,201,29,201,28,229,31,39,31,234,31,206,31,206,30,206,29,193,31,45,31,45,30,232,31,216,31,26,31,247,31,52,31,11,31,1,31,1,30,77,31,242,31,106,31,9,31,140,31,140,30,244,31,74,31,77,31,11,31,249,31,126,31,156,31,121,31,104,31,140,31,19,31,90,31,130,31,239,31,63,31,218,31,190,31,223,31,223,30,151,31,237,31,237,30,253,31,90,31,7,31,237,31,72,31,121,31,118,31,251,31,141,31,173,31,76,31,201,31,93,31,193,31,207,31,154,31,239,31,80,31,80,30,80,29,209,31,39,31,231,31,231,31,231,30,238,31,189,31,111,31,25,31,200,31,200,30,98,31,98,30,68,31,187,31,4,31,245,31,20,31,205,31,28,31,90,31,112,31,61,31,212,31,75,31,132,31,252,31,83,31,97,31,6,31,6,30,220,31,241,31,26,31,17,31,148,31,40,31,49,31,49,30,67,31,89,31,209,31,150,31,182,31,210,31,126,31,75,31,215,31,194,31,93,31,93,31,66,31,66,30,133,31,132,31,189,31,189,30,230,31,230,31,198,31,250,31,250,30,250,29,250,28,184,31,65,31,65,30,168,31,175,31,175,30,254,31,254,30,195,31,6,31,253,31,26,31,155,31,155,30,239,31,229,31,229,30,197,31,197,30,75,31,27,31,27,30,235,31,101,31,101,30,18,31,141,31,89,31,89,30,239,31,239,30,96,31,96,30,243,31,243,30,128,31,94,31,118,31,53,31,3,31,3,30,45,31,157,31,207,31,162,31,162,30,129,31,180,31,178,31,178,30,178,29,214,31,41,31,43,31,208,31,201,31,127,31,26,31,134,31,202,31,21,31,21,30,225,31,187,31,99,31,20,31,244,31,226,31,226,30,253,31,60,31,202,31,148,31,148,30,148,29,103,31,238,31,58,31,138,31,111,31,52,31,181,31,39,31,109,31,250,31,49,31,86,31,86,30,104,31,248,31,62,31,203,31,214,31,91,31,252,31,177,31,223,31,151,31,224,31,108,31,96,31,172,31,137,31,137,30,45,31,186,31,71,31,71,30,252,31,44,31,3,31,231,31,203,31,229,31,223,31,223,30,125,31,125,30,135,31,102,31,102,30,37,31,239,31,54,31,176,31,176,30,212,31,46,31,216,31,216,30,168,31,168,30,168,29,168,28,17,31,31,31,113,31,48,31,48,30,87,31,217,31,182,31,29,31,184,31,20,31,180,31,88,31,24,31,112,31,97,31,187,31,209,31,109,31,109,30,109,29,109,28,195,31,202,31,70,31,57,31,156,31,156,30,153,31,135,31,135,30,171,31,94,31,232,31,146,31,48,31,89,31,228,31,72,31,72,30,61,31,70,31,8,31,178,31,56,31,206,31,10,31,91,31,147,31,147,30,40,31,78,31,23,31,33,31,33,30,33,29,5,31,67,31,63,31,48,31,80,31,25,31,149,31,112,31,109,31,155,31,75,31,95,31,94,31,94,31,51,31,7,31,68,31,56,31,56,30,56,29,56,28,56,27,118,31,247,31,168,31,15,31,117,31,208,31,24,31,211,31,195,31,195,30,24,31,24,30,222,31,222,30,222,29,222,31,57,31,207,31,207,30,183,31,84,31,84,30,177,31,61,31,76,31,101,31,184,31,42,31,55,31,55,30,20,31,134,31,134,30,243,31,2,31,103,31,87,31,161,31,161,30,134,31,188,31,12,31,42,31,203,31,251,31,51,31,53,31,53,30,53,29,53,28,178,31,178,30,249,31,124,31,124,30,80,31,40,31,41,31,206,31,90,31,90,30,90,29,32,31,32,30,131,31,154,31,58,31,69,31,144,31,117,31,161,31,161,30,161,29,122,31,6,31,52,31,199,31,199,30,20,31,225,31,225,30,117,31,16,31,97,31,97,30,190,31,133,31,198,31,11,31,11,30,93,31,68,31,149,31,21,31,92,31,212,31,212,30,212,29,185,31,227,31,45,31,45,30,144,31,218,31,80,31,147,31,8,31,125,31,44,31,206,31,179,31,112,31,32,31,81,31,101,31,240,31,240,30,76,31,14,31,160,31,164,31,164,30,25,31,58,31,22,31,22,30,22,29,177,31,70,31,130,31,130,30,12,31,46,31,211,31,211,30,56,31,56,30,81,31,159,31,148,31,148,30,173,31,90,31,202,31,160,31,146,31,146,30,83,31,186,31,135,31,169,31,161,31,105,31,88,31,9,31,199,31,89,31,172,31,236,31,231,31,247,31,102,31,171,31,78,31,202,31,15,31,220,31,108,31,53,31,53,30,42,31,223,31,223,30,104,31,57,31,216,31,216,30,94,31,93,31,35,31,10,31,5,31,242,31,44,31,151,31,17,31,41,31,41,30,13,31,13,30,89,31,233,31,87,31,87,30,90,31,90,30,132,31,129,31,231,31,144,31,36,31,255,31,255,30,129,31,125,31,122,31,122,30,23,31,101,31,25,31,25,30,87,31,250,31,151,31,205,31,147,31,184,31,152,31,152,30,37,31,67,31,190,31,109,31,140,31,48,31,38,31,228,31,251,31,251,30,204,31,41,31,41,30,198,31,48,31,50,31,47,31,145,31,145,30,27,31,246,31,97,31,197,31,197,30,43,31,211,31,81,31,245,31,245,30,26,31,248,31,176,31,73,31,193,31,62,31,150,31,125,31,196,31,227,31,4,31,86,31,238,31,175,31,44,31,210,31,122,31,122,30,68,31,68,30,39,31,60,31,60,30,151,31,181,31,142,31,8,31,35,31,120,31,195,31,190,31,190,30,66,31,51,31,46,31,182,31,223,31,188,31,82,31,34,31,29,31,115,31,169,31,169,30,169,29,143,31,174,31,131,31,21,31,111,31,111,30,108,31,230,31,230,30,23,31,79,31,86,31,86,30,7,31,9,31,1,31,60,31,209,31,148,31,148,30,62,31,73,31,65,31,65,30,53,31,53,30,44,31,203,31,129,31,22,31,213,31,50,31,40,31,51,31,67,31,67,30,236,31,196,31,37,31,150,31,1,31,254,31,219,31,219,30,219,29,69,31,173,31,43,31,236,31,74,31,74,30,20,31,113,31,113,30,113,29,47,31,131,31,110,31,113,31,67,31,67,30,67,29,186,31,26,31,87,31,213,31,213,30,61,31,84,31,78,31,172,31,240,31,202,31,79,31,79,30,72,31,69,31,107,31,107,30,202,31,202,30,202,29,124,31,124,30,247,31,247,30,143,31,27,31,205,31,198,31,78,31,78,30,241,31,245,31,245,31,245,30,83,31,83,30,41,31,89,31,89,30,21,31,153,31,130,31,130,30,210,31,57,31,152,31,226,31,70,31,214,31,214,30,214,29,217,31,169,31,9,31,147,31,80,31,170,31,56,31,64,31,3,31,187,31,16,31,21,31,8,31,80,31,80,30,11,31,11,30,215,31,107,31,194,31,162,31,162,30,1,31,139,31,23,31,23,30,23,29,30,31,197,31,18,31,28,31,60,31,21,31,90,31,155,31,79,31,104,31,202,31,202,30,200,31,254,31,97,31,6,31,6,30,114,31,183,31,162,31,162,30,234,31,23,31,212,31,96,31,90,31,90,30,100,31,194,31,82,31,138,31,94,31,2,31,143,31,251,31,32,31,34,31,34,30,108,31,12,31,8,31,8,31,109,31,97,31,44,31,18,31,214,31,217,31,38,31,116,31,116,30,116,29,116,28,116,27,33,31,133,31,48,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
