-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 660;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (145,0,172,0,0,0,233,0,174,0,74,0,61,0,0,0,159,0,119,0,168,0,45,0,0,0,11,0,0,0,122,0,73,0,0,0,195,0,0,0,29,0,0,0,31,0,247,0,3,0,121,0,60,0,0,0,82,0,125,0,234,0,202,0,155,0,147,0,59,0,191,0,125,0,44,0,204,0,89,0,101,0,0,0,0,0,80,0,70,0,158,0,238,0,137,0,0,0,242,0,250,0,22,0,23,0,129,0,248,0,138,0,118,0,13,0,132,0,178,0,175,0,0,0,0,0,172,0,22,0,177,0,172,0,63,0,120,0,138,0,30,0,235,0,75,0,180,0,0,0,223,0,0,0,140,0,42,0,0,0,131,0,130,0,0,0,46,0,195,0,95,0,231,0,142,0,160,0,57,0,159,0,35,0,0,0,135,0,208,0,0,0,86,0,194,0,0,0,127,0,105,0,176,0,5,0,0,0,42,0,201,0,224,0,96,0,169,0,104,0,24,0,0,0,0,0,86,0,0,0,0,0,0,0,201,0,122,0,40,0,0,0,170,0,107,0,56,0,82,0,141,0,25,0,0,0,74,0,0,0,101,0,14,0,1,0,9,0,154,0,25,0,211,0,101,0,0,0,229,0,190,0,85,0,200,0,236,0,15,0,80,0,0,0,0,0,0,0,0,0,122,0,0,0,195,0,0,0,0,0,81,0,104,0,0,0,101,0,255,0,126,0,0,0,232,0,0,0,66,0,0,0,25,0,253,0,78,0,0,0,244,0,235,0,0,0,0,0,44,0,0,0,68,0,62,0,15,0,179,0,181,0,51,0,112,0,0,0,44,0,89,0,84,0,121,0,244,0,243,0,224,0,196,0,137,0,7,0,177,0,28,0,223,0,0,0,217,0,249,0,125,0,195,0,115,0,164,0,87,0,175,0,74,0,161,0,146,0,158,0,0,0,0,0,43,0,149,0,198,0,116,0,214,0,180,0,33,0,222,0,206,0,250,0,0,0,0,0,250,0,235,0,253,0,152,0,228,0,202,0,107,0,147,0,22,0,182,0,220,0,38,0,115,0,155,0,35,0,179,0,0,0,76,0,0,0,136,0,29,0,0,0,68,0,240,0,208,0,29,0,0,0,208,0,0,0,211,0,173,0,0,0,241,0,221,0,7,0,206,0,123,0,0,0,75,0,0,0,237,0,134,0,126,0,44,0,128,0,211,0,251,0,116,0,172,0,40,0,107,0,105,0,254,0,154,0,154,0,0,0,8,0,32,0,77,0,248,0,241,0,0,0,4,0,119,0,0,0,69,0,145,0,22,0,94,0,0,0,0,0,83,0,13,0,138,0,0,0,182,0,92,0,108,0,172,0,203,0,22,0,0,0,244,0,97,0,165,0,24,0,255,0,7,0,242,0,209,0,0,0,98,0,0,0,28,0,74,0,225,0,103,0,18,0,253,0,197,0,123,0,54,0,18,0,0,0,7,0,205,0,8,0,159,0,236,0,94,0,83,0,0,0,228,0,160,0,181,0,197,0,241,0,106,0,184,0,0,0,195,0,0,0,0,0,198,0,0,0,141,0,0,0,99,0,77,0,38,0,48,0,94,0,0,0,51,0,128,0,126,0,151,0,39,0,33,0,0,0,200,0,78,0,205,0,147,0,115,0,176,0,213,0,118,0,192,0,236,0,60,0,102,0,63,0,0,0,229,0,0,0,225,0,128,0,184,0,242,0,101,0,124,0,107,0,104,0,0,0,163,0,0,0,77,0,0,0,0,0,71,0,58,0,43,0,133,0,0,0,79,0,247,0,127,0,3,0,211,0,126,0,0,0,196,0,55,0,208,0,138,0,166,0,88,0,52,0,209,0,0,0,56,0,74,0,35,0,216,0,123,0,167,0,0,0,0,0,220,0,72,0,192,0,77,0,245,0,190,0,51,0,242,0,22,0,159,0,120,0,82,0,0,0,65,0,0,0,0,0,160,0,244,0,242,0,15,0,194,0,14,0,0,0,11,0,170,0,223,0,0,0,110,0,212,0,104,0,160,0,111,0,119,0,0,0,34,0,92,0,169,0,131,0,193,0,247,0,85,0,95,0,201,0,131,0,129,0,150,0,0,0,113,0,0,0,50,0,166,0,104,0,35,0,89,0,0,0,19,0,55,0,136,0,134,0,0,0,197,0,0,0,147,0,241,0,0,0,254,0,0,0,205,0,36,0,142,0,71,0,164,0,8,0,0,0,78,0,250,0,127,0,125,0,92,0,0,0,0,0,0,0,22,0,83,0,184,0,0,0,178,0,55,0,205,0,54,0,0,0,51,0,127,0,44,0,0,0,99,0,218,0,111,0,0,0,233,0,223,0,5,0,108,0,0,0,6,0,237,0,0,0,173,0,0,0,49,0,0,0,205,0,0,0,241,0,148,0,0,0,34,0,0,0,84,0,120,0,158,0,21,0,0,0,184,0,211,0,85,0,46,0,217,0,141,0,0,0,0,0,156,0,66,0,0,0,73,0,30,0,153,0,112,0,242,0,223,0,43,0,57,0,215,0,197,0,250,0,204,0,86,0,8,0,198,0,189,0,148,0,6,0,64,0,0,0,12,0,235,0,121,0,165,0,0,0,142,0,180,0,230,0,0,0,0,0,157,0,187,0,14,0,156,0,210,0,135,0,0,0,232,0,102,0,75,0,237,0,234,0,247,0,241,0,251,0,0,0,0,0,213,0,0,0,165,0,96,0,253,0,0,0,220,0,0,0,177,0,89,0,209,0,52,0,143,0,227,0,138,0,0,0,23,0,139,0,0,0,250,0,18,0,20,0,1,0,0,0,167,0,68,0,243,0,112,0,197,0,2,0,165,0,94,0,19,0,195,0,130,0,0,0,0,0,124,0,137,0,207,0,232,0,199,0,0,0,131,0,102,0,69,0,57,0,206,0,0,0,138,0,0,0,134,0,65,0,0,0,252,0,133,0);
signal scenario_full  : scenario_type := (145,31,172,31,172,30,233,31,174,31,74,31,61,31,61,30,159,31,119,31,168,31,45,31,45,30,11,31,11,30,122,31,73,31,73,30,195,31,195,30,29,31,29,30,31,31,247,31,3,31,121,31,60,31,60,30,82,31,125,31,234,31,202,31,155,31,147,31,59,31,191,31,125,31,44,31,204,31,89,31,101,31,101,30,101,29,80,31,70,31,158,31,238,31,137,31,137,30,242,31,250,31,22,31,23,31,129,31,248,31,138,31,118,31,13,31,132,31,178,31,175,31,175,30,175,29,172,31,22,31,177,31,172,31,63,31,120,31,138,31,30,31,235,31,75,31,180,31,180,30,223,31,223,30,140,31,42,31,42,30,131,31,130,31,130,30,46,31,195,31,95,31,231,31,142,31,160,31,57,31,159,31,35,31,35,30,135,31,208,31,208,30,86,31,194,31,194,30,127,31,105,31,176,31,5,31,5,30,42,31,201,31,224,31,96,31,169,31,104,31,24,31,24,30,24,29,86,31,86,30,86,29,86,28,201,31,122,31,40,31,40,30,170,31,107,31,56,31,82,31,141,31,25,31,25,30,74,31,74,30,101,31,14,31,1,31,9,31,154,31,25,31,211,31,101,31,101,30,229,31,190,31,85,31,200,31,236,31,15,31,80,31,80,30,80,29,80,28,80,27,122,31,122,30,195,31,195,30,195,29,81,31,104,31,104,30,101,31,255,31,126,31,126,30,232,31,232,30,66,31,66,30,25,31,253,31,78,31,78,30,244,31,235,31,235,30,235,29,44,31,44,30,68,31,62,31,15,31,179,31,181,31,51,31,112,31,112,30,44,31,89,31,84,31,121,31,244,31,243,31,224,31,196,31,137,31,7,31,177,31,28,31,223,31,223,30,217,31,249,31,125,31,195,31,115,31,164,31,87,31,175,31,74,31,161,31,146,31,158,31,158,30,158,29,43,31,149,31,198,31,116,31,214,31,180,31,33,31,222,31,206,31,250,31,250,30,250,29,250,31,235,31,253,31,152,31,228,31,202,31,107,31,147,31,22,31,182,31,220,31,38,31,115,31,155,31,35,31,179,31,179,30,76,31,76,30,136,31,29,31,29,30,68,31,240,31,208,31,29,31,29,30,208,31,208,30,211,31,173,31,173,30,241,31,221,31,7,31,206,31,123,31,123,30,75,31,75,30,237,31,134,31,126,31,44,31,128,31,211,31,251,31,116,31,172,31,40,31,107,31,105,31,254,31,154,31,154,31,154,30,8,31,32,31,77,31,248,31,241,31,241,30,4,31,119,31,119,30,69,31,145,31,22,31,94,31,94,30,94,29,83,31,13,31,138,31,138,30,182,31,92,31,108,31,172,31,203,31,22,31,22,30,244,31,97,31,165,31,24,31,255,31,7,31,242,31,209,31,209,30,98,31,98,30,28,31,74,31,225,31,103,31,18,31,253,31,197,31,123,31,54,31,18,31,18,30,7,31,205,31,8,31,159,31,236,31,94,31,83,31,83,30,228,31,160,31,181,31,197,31,241,31,106,31,184,31,184,30,195,31,195,30,195,29,198,31,198,30,141,31,141,30,99,31,77,31,38,31,48,31,94,31,94,30,51,31,128,31,126,31,151,31,39,31,33,31,33,30,200,31,78,31,205,31,147,31,115,31,176,31,213,31,118,31,192,31,236,31,60,31,102,31,63,31,63,30,229,31,229,30,225,31,128,31,184,31,242,31,101,31,124,31,107,31,104,31,104,30,163,31,163,30,77,31,77,30,77,29,71,31,58,31,43,31,133,31,133,30,79,31,247,31,127,31,3,31,211,31,126,31,126,30,196,31,55,31,208,31,138,31,166,31,88,31,52,31,209,31,209,30,56,31,74,31,35,31,216,31,123,31,167,31,167,30,167,29,220,31,72,31,192,31,77,31,245,31,190,31,51,31,242,31,22,31,159,31,120,31,82,31,82,30,65,31,65,30,65,29,160,31,244,31,242,31,15,31,194,31,14,31,14,30,11,31,170,31,223,31,223,30,110,31,212,31,104,31,160,31,111,31,119,31,119,30,34,31,92,31,169,31,131,31,193,31,247,31,85,31,95,31,201,31,131,31,129,31,150,31,150,30,113,31,113,30,50,31,166,31,104,31,35,31,89,31,89,30,19,31,55,31,136,31,134,31,134,30,197,31,197,30,147,31,241,31,241,30,254,31,254,30,205,31,36,31,142,31,71,31,164,31,8,31,8,30,78,31,250,31,127,31,125,31,92,31,92,30,92,29,92,28,22,31,83,31,184,31,184,30,178,31,55,31,205,31,54,31,54,30,51,31,127,31,44,31,44,30,99,31,218,31,111,31,111,30,233,31,223,31,5,31,108,31,108,30,6,31,237,31,237,30,173,31,173,30,49,31,49,30,205,31,205,30,241,31,148,31,148,30,34,31,34,30,84,31,120,31,158,31,21,31,21,30,184,31,211,31,85,31,46,31,217,31,141,31,141,30,141,29,156,31,66,31,66,30,73,31,30,31,153,31,112,31,242,31,223,31,43,31,57,31,215,31,197,31,250,31,204,31,86,31,8,31,198,31,189,31,148,31,6,31,64,31,64,30,12,31,235,31,121,31,165,31,165,30,142,31,180,31,230,31,230,30,230,29,157,31,187,31,14,31,156,31,210,31,135,31,135,30,232,31,102,31,75,31,237,31,234,31,247,31,241,31,251,31,251,30,251,29,213,31,213,30,165,31,96,31,253,31,253,30,220,31,220,30,177,31,89,31,209,31,52,31,143,31,227,31,138,31,138,30,23,31,139,31,139,30,250,31,18,31,20,31,1,31,1,30,167,31,68,31,243,31,112,31,197,31,2,31,165,31,94,31,19,31,195,31,130,31,130,30,130,29,124,31,137,31,207,31,232,31,199,31,199,30,131,31,102,31,69,31,57,31,206,31,206,30,138,31,138,30,134,31,65,31,65,30,252,31,133,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
