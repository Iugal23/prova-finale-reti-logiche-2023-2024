-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 821;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (56,0,0,0,124,0,238,0,199,0,0,0,102,0,0,0,224,0,67,0,194,0,217,0,126,0,214,0,137,0,69,0,145,0,43,0,182,0,173,0,0,0,185,0,212,0,0,0,174,0,73,0,0,0,92,0,39,0,191,0,212,0,153,0,183,0,0,0,130,0,28,0,0,0,149,0,105,0,170,0,0,0,122,0,61,0,42,0,177,0,178,0,77,0,24,0,217,0,15,0,197,0,0,0,175,0,52,0,90,0,147,0,0,0,246,0,92,0,0,0,20,0,232,0,230,0,167,0,0,0,134,0,30,0,229,0,195,0,52,0,98,0,241,0,0,0,164,0,206,0,102,0,191,0,129,0,77,0,0,0,15,0,24,0,134,0,0,0,233,0,142,0,25,0,0,0,0,0,48,0,144,0,0,0,80,0,195,0,107,0,167,0,0,0,75,0,0,0,223,0,0,0,30,0,242,0,34,0,196,0,230,0,220,0,219,0,8,0,0,0,114,0,104,0,0,0,21,0,54,0,156,0,0,0,57,0,19,0,96,0,221,0,142,0,130,0,241,0,173,0,51,0,199,0,0,0,120,0,61,0,124,0,177,0,36,0,246,0,88,0,0,0,191,0,84,0,10,0,12,0,176,0,135,0,85,0,0,0,244,0,13,0,194,0,0,0,128,0,66,0,160,0,218,0,98,0,118,0,0,0,0,0,135,0,86,0,174,0,16,0,41,0,216,0,123,0,209,0,46,0,0,0,101,0,82,0,134,0,159,0,157,0,104,0,74,0,73,0,0,0,41,0,0,0,0,0,236,0,47,0,207,0,195,0,128,0,169,0,226,0,77,0,170,0,89,0,123,0,220,0,0,0,0,0,90,0,194,0,147,0,0,0,242,0,208,0,9,0,203,0,20,0,0,0,33,0,181,0,66,0,34,0,57,0,159,0,201,0,182,0,0,0,250,0,0,0,41,0,253,0,46,0,121,0,37,0,0,0,139,0,72,0,153,0,188,0,135,0,37,0,207,0,227,0,116,0,194,0,161,0,255,0,24,0,160,0,40,0,79,0,26,0,226,0,0,0,208,0,0,0,230,0,44,0,224,0,135,0,51,0,252,0,0,0,254,0,21,0,251,0,25,0,100,0,125,0,223,0,0,0,96,0,55,0,156,0,243,0,227,0,0,0,124,0,1,0,6,0,100,0,150,0,178,0,91,0,116,0,143,0,244,0,161,0,60,0,97,0,234,0,3,0,0,0,0,0,0,0,147,0,99,0,185,0,231,0,4,0,0,0,208,0,0,0,137,0,212,0,40,0,138,0,0,0,16,0,33,0,0,0,172,0,41,0,213,0,192,0,148,0,170,0,34,0,106,0,62,0,101,0,252,0,195,0,16,0,217,0,77,0,39,0,184,0,137,0,200,0,174,0,227,0,178,0,0,0,0,0,38,0,0,0,116,0,241,0,122,0,5,0,40,0,66,0,136,0,11,0,0,0,0,0,237,0,199,0,42,0,68,0,199,0,167,0,137,0,238,0,83,0,0,0,197,0,112,0,0,0,6,0,0,0,32,0,0,0,125,0,222,0,160,0,98,0,65,0,0,0,0,0,0,0,163,0,6,0,227,0,0,0,94,0,128,0,90,0,134,0,103,0,0,0,130,0,141,0,160,0,225,0,68,0,29,0,0,0,90,0,0,0,230,0,126,0,237,0,233,0,66,0,172,0,0,0,67,0,0,0,53,0,0,0,0,0,127,0,63,0,71,0,90,0,0,0,219,0,60,0,4,0,0,0,196,0,0,0,52,0,240,0,0,0,36,0,205,0,0,0,184,0,15,0,113,0,113,0,145,0,154,0,4,0,0,0,0,0,143,0,0,0,0,0,0,0,65,0,162,0,20,0,164,0,223,0,135,0,105,0,1,0,169,0,145,0,44,0,133,0,199,0,59,0,117,0,229,0,0,0,163,0,144,0,54,0,174,0,96,0,204,0,0,0,56,0,145,0,121,0,0,0,105,0,81,0,198,0,152,0,0,0,0,0,47,0,124,0,121,0,171,0,66,0,99,0,52,0,137,0,160,0,93,0,0,0,199,0,44,0,191,0,140,0,9,0,0,0,79,0,122,0,0,0,0,0,47,0,0,0,124,0,78,0,0,0,242,0,184,0,0,0,155,0,85,0,0,0,227,0,66,0,168,0,106,0,254,0,0,0,23,0,219,0,248,0,152,0,194,0,20,0,127,0,51,0,39,0,110,0,56,0,140,0,214,0,193,0,148,0,0,0,221,0,0,0,19,0,220,0,0,0,250,0,133,0,0,0,52,0,113,0,239,0,142,0,241,0,0,0,0,0,203,0,56,0,0,0,245,0,75,0,69,0,0,0,0,0,18,0,112,0,150,0,191,0,21,0,0,0,15,0,0,0,152,0,15,0,0,0,0,0,170,0,64,0,37,0,23,0,125,0,87,0,152,0,60,0,219,0,126,0,239,0,0,0,229,0,61,0,250,0,207,0,101,0,0,0,104,0,0,0,0,0,172,0,143,0,0,0,44,0,117,0,151,0,42,0,0,0,95,0,51,0,0,0,33,0,57,0,0,0,230,0,70,0,174,0,140,0,80,0,0,0,210,0,235,0,0,0,0,0,0,0,70,0,84,0,241,0,0,0,113,0,165,0,60,0,71,0,178,0,0,0,0,0,46,0,0,0,157,0,0,0,200,0,76,0,250,0,107,0,117,0,183,0,136,0,58,0,2,0,210,0,0,0,235,0,135,0,0,0,176,0,0,0,44,0,133,0,108,0,0,0,103,0,0,0,223,0,90,0,77,0,253,0,54,0,216,0,206,0,0,0,118,0,89,0,33,0,234,0,2,0,50,0,0,0,243,0,42,0,0,0,215,0,154,0,0,0,97,0,188,0,36,0,123,0,162,0,68,0,0,0,0,0,100,0,152,0,11,0,206,0,0,0,125,0,20,0,219,0,120,0,1,0,119,0,122,0,196,0,34,0,0,0,125,0,19,0,161,0,123,0,151,0,0,0,180,0,188,0,238,0,50,0,252,0,0,0,76,0,0,0,249,0,238,0,168,0,0,0,164,0,140,0,21,0,0,0,0,0,227,0,11,0,98,0,22,0,119,0,1,0,0,0,147,0,143,0,122,0,43,0,0,0,220,0,141,0,103,0,11,0,87,0,190,0,121,0,214,0,91,0,37,0,184,0,0,0,0,0,242,0,123,0,216,0,9,0,0,0,196,0,82,0,193,0,225,0,8,0,182,0,148,0,157,0,189,0,102,0,232,0,89,0,42,0,224,0,0,0,147,0,73,0,0,0,51,0,83,0,0,0,0,0,182,0,251,0,0,0,242,0,124,0,0,0,33,0,0,0,0,0,0,0,204,0,0,0,208,0,144,0,0,0,96,0,224,0,0,0,0,0,117,0,0,0,0,0,44,0,48,0,250,0,33,0,51,0,137,0,85,0,140,0,64,0,80,0,178,0,18,0,155,0,239,0,251,0,65,0,71,0,213,0,25,0,203,0,204,0,0,0,0,0,79,0,151,0,217,0,0,0,139,0,86,0,83,0,89,0,186,0,123,0,221,0,155,0,188,0,6,0,138,0,211,0,218,0,170,0,0,0,238,0,37,0,0,0,65,0,0,0,0,0,205,0,35,0,248,0,213,0,61,0,211,0,142,0,0,0,216,0);
signal scenario_full  : scenario_type := (56,31,56,30,124,31,238,31,199,31,199,30,102,31,102,30,224,31,67,31,194,31,217,31,126,31,214,31,137,31,69,31,145,31,43,31,182,31,173,31,173,30,185,31,212,31,212,30,174,31,73,31,73,30,92,31,39,31,191,31,212,31,153,31,183,31,183,30,130,31,28,31,28,30,149,31,105,31,170,31,170,30,122,31,61,31,42,31,177,31,178,31,77,31,24,31,217,31,15,31,197,31,197,30,175,31,52,31,90,31,147,31,147,30,246,31,92,31,92,30,20,31,232,31,230,31,167,31,167,30,134,31,30,31,229,31,195,31,52,31,98,31,241,31,241,30,164,31,206,31,102,31,191,31,129,31,77,31,77,30,15,31,24,31,134,31,134,30,233,31,142,31,25,31,25,30,25,29,48,31,144,31,144,30,80,31,195,31,107,31,167,31,167,30,75,31,75,30,223,31,223,30,30,31,242,31,34,31,196,31,230,31,220,31,219,31,8,31,8,30,114,31,104,31,104,30,21,31,54,31,156,31,156,30,57,31,19,31,96,31,221,31,142,31,130,31,241,31,173,31,51,31,199,31,199,30,120,31,61,31,124,31,177,31,36,31,246,31,88,31,88,30,191,31,84,31,10,31,12,31,176,31,135,31,85,31,85,30,244,31,13,31,194,31,194,30,128,31,66,31,160,31,218,31,98,31,118,31,118,30,118,29,135,31,86,31,174,31,16,31,41,31,216,31,123,31,209,31,46,31,46,30,101,31,82,31,134,31,159,31,157,31,104,31,74,31,73,31,73,30,41,31,41,30,41,29,236,31,47,31,207,31,195,31,128,31,169,31,226,31,77,31,170,31,89,31,123,31,220,31,220,30,220,29,90,31,194,31,147,31,147,30,242,31,208,31,9,31,203,31,20,31,20,30,33,31,181,31,66,31,34,31,57,31,159,31,201,31,182,31,182,30,250,31,250,30,41,31,253,31,46,31,121,31,37,31,37,30,139,31,72,31,153,31,188,31,135,31,37,31,207,31,227,31,116,31,194,31,161,31,255,31,24,31,160,31,40,31,79,31,26,31,226,31,226,30,208,31,208,30,230,31,44,31,224,31,135,31,51,31,252,31,252,30,254,31,21,31,251,31,25,31,100,31,125,31,223,31,223,30,96,31,55,31,156,31,243,31,227,31,227,30,124,31,1,31,6,31,100,31,150,31,178,31,91,31,116,31,143,31,244,31,161,31,60,31,97,31,234,31,3,31,3,30,3,29,3,28,147,31,99,31,185,31,231,31,4,31,4,30,208,31,208,30,137,31,212,31,40,31,138,31,138,30,16,31,33,31,33,30,172,31,41,31,213,31,192,31,148,31,170,31,34,31,106,31,62,31,101,31,252,31,195,31,16,31,217,31,77,31,39,31,184,31,137,31,200,31,174,31,227,31,178,31,178,30,178,29,38,31,38,30,116,31,241,31,122,31,5,31,40,31,66,31,136,31,11,31,11,30,11,29,237,31,199,31,42,31,68,31,199,31,167,31,137,31,238,31,83,31,83,30,197,31,112,31,112,30,6,31,6,30,32,31,32,30,125,31,222,31,160,31,98,31,65,31,65,30,65,29,65,28,163,31,6,31,227,31,227,30,94,31,128,31,90,31,134,31,103,31,103,30,130,31,141,31,160,31,225,31,68,31,29,31,29,30,90,31,90,30,230,31,126,31,237,31,233,31,66,31,172,31,172,30,67,31,67,30,53,31,53,30,53,29,127,31,63,31,71,31,90,31,90,30,219,31,60,31,4,31,4,30,196,31,196,30,52,31,240,31,240,30,36,31,205,31,205,30,184,31,15,31,113,31,113,31,145,31,154,31,4,31,4,30,4,29,143,31,143,30,143,29,143,28,65,31,162,31,20,31,164,31,223,31,135,31,105,31,1,31,169,31,145,31,44,31,133,31,199,31,59,31,117,31,229,31,229,30,163,31,144,31,54,31,174,31,96,31,204,31,204,30,56,31,145,31,121,31,121,30,105,31,81,31,198,31,152,31,152,30,152,29,47,31,124,31,121,31,171,31,66,31,99,31,52,31,137,31,160,31,93,31,93,30,199,31,44,31,191,31,140,31,9,31,9,30,79,31,122,31,122,30,122,29,47,31,47,30,124,31,78,31,78,30,242,31,184,31,184,30,155,31,85,31,85,30,227,31,66,31,168,31,106,31,254,31,254,30,23,31,219,31,248,31,152,31,194,31,20,31,127,31,51,31,39,31,110,31,56,31,140,31,214,31,193,31,148,31,148,30,221,31,221,30,19,31,220,31,220,30,250,31,133,31,133,30,52,31,113,31,239,31,142,31,241,31,241,30,241,29,203,31,56,31,56,30,245,31,75,31,69,31,69,30,69,29,18,31,112,31,150,31,191,31,21,31,21,30,15,31,15,30,152,31,15,31,15,30,15,29,170,31,64,31,37,31,23,31,125,31,87,31,152,31,60,31,219,31,126,31,239,31,239,30,229,31,61,31,250,31,207,31,101,31,101,30,104,31,104,30,104,29,172,31,143,31,143,30,44,31,117,31,151,31,42,31,42,30,95,31,51,31,51,30,33,31,57,31,57,30,230,31,70,31,174,31,140,31,80,31,80,30,210,31,235,31,235,30,235,29,235,28,70,31,84,31,241,31,241,30,113,31,165,31,60,31,71,31,178,31,178,30,178,29,46,31,46,30,157,31,157,30,200,31,76,31,250,31,107,31,117,31,183,31,136,31,58,31,2,31,210,31,210,30,235,31,135,31,135,30,176,31,176,30,44,31,133,31,108,31,108,30,103,31,103,30,223,31,90,31,77,31,253,31,54,31,216,31,206,31,206,30,118,31,89,31,33,31,234,31,2,31,50,31,50,30,243,31,42,31,42,30,215,31,154,31,154,30,97,31,188,31,36,31,123,31,162,31,68,31,68,30,68,29,100,31,152,31,11,31,206,31,206,30,125,31,20,31,219,31,120,31,1,31,119,31,122,31,196,31,34,31,34,30,125,31,19,31,161,31,123,31,151,31,151,30,180,31,188,31,238,31,50,31,252,31,252,30,76,31,76,30,249,31,238,31,168,31,168,30,164,31,140,31,21,31,21,30,21,29,227,31,11,31,98,31,22,31,119,31,1,31,1,30,147,31,143,31,122,31,43,31,43,30,220,31,141,31,103,31,11,31,87,31,190,31,121,31,214,31,91,31,37,31,184,31,184,30,184,29,242,31,123,31,216,31,9,31,9,30,196,31,82,31,193,31,225,31,8,31,182,31,148,31,157,31,189,31,102,31,232,31,89,31,42,31,224,31,224,30,147,31,73,31,73,30,51,31,83,31,83,30,83,29,182,31,251,31,251,30,242,31,124,31,124,30,33,31,33,30,33,29,33,28,204,31,204,30,208,31,144,31,144,30,96,31,224,31,224,30,224,29,117,31,117,30,117,29,44,31,48,31,250,31,33,31,51,31,137,31,85,31,140,31,64,31,80,31,178,31,18,31,155,31,239,31,251,31,65,31,71,31,213,31,25,31,203,31,204,31,204,30,204,29,79,31,151,31,217,31,217,30,139,31,86,31,83,31,89,31,186,31,123,31,221,31,155,31,188,31,6,31,138,31,211,31,218,31,170,31,170,30,238,31,37,31,37,30,65,31,65,30,65,29,205,31,35,31,248,31,213,31,61,31,211,31,142,31,142,30,216,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
