-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_657 is
end project_tb_657;

architecture project_tb_arch_657 of project_tb_657 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 630;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,247,0,65,0,124,0,68,0,141,0,188,0,111,0,128,0,134,0,134,0,93,0,222,0,122,0,70,0,214,0,95,0,230,0,18,0,0,0,90,0,123,0,0,0,220,0,70,0,0,0,136,0,0,0,172,0,156,0,126,0,0,0,0,0,47,0,254,0,130,0,11,0,44,0,162,0,0,0,70,0,190,0,164,0,57,0,198,0,9,0,247,0,184,0,211,0,62,0,0,0,0,0,138,0,14,0,23,0,89,0,98,0,143,0,0,0,253,0,111,0,215,0,200,0,197,0,0,0,240,0,0,0,23,0,113,0,81,0,0,0,249,0,66,0,0,0,253,0,0,0,76,0,209,0,232,0,0,0,187,0,226,0,150,0,195,0,0,0,214,0,0,0,139,0,223,0,0,0,163,0,95,0,248,0,193,0,239,0,141,0,0,0,126,0,0,0,96,0,0,0,107,0,0,0,0,0,239,0,51,0,45,0,0,0,0,0,0,0,0,0,220,0,12,0,64,0,126,0,232,0,189,0,0,0,0,0,0,0,180,0,243,0,126,0,238,0,184,0,0,0,153,0,242,0,0,0,57,0,43,0,104,0,220,0,140,0,0,0,86,0,101,0,0,0,209,0,0,0,188,0,0,0,83,0,229,0,240,0,69,0,94,0,55,0,22,0,78,0,153,0,102,0,0,0,93,0,245,0,0,0,8,0,199,0,192,0,226,0,0,0,0,0,100,0,96,0,19,0,236,0,0,0,116,0,57,0,199,0,33,0,0,0,0,0,39,0,0,0,0,0,160,0,223,0,0,0,251,0,84,0,69,0,141,0,226,0,0,0,22,0,234,0,168,0,163,0,191,0,12,0,244,0,246,0,143,0,172,0,220,0,90,0,86,0,0,0,28,0,0,0,15,0,251,0,15,0,207,0,219,0,0,0,73,0,100,0,113,0,24,0,0,0,27,0,0,0,51,0,111,0,0,0,167,0,0,0,184,0,0,0,242,0,193,0,52,0,243,0,249,0,123,0,58,0,237,0,73,0,223,0,81,0,11,0,226,0,0,0,23,0,110,0,0,0,0,0,132,0,246,0,128,0,90,0,239,0,176,0,103,0,30,0,0,0,233,0,31,0,57,0,37,0,205,0,62,0,202,0,0,0,0,0,97,0,93,0,67,0,0,0,147,0,0,0,39,0,252,0,0,0,0,0,0,0,129,0,148,0,69,0,141,0,64,0,108,0,246,0,45,0,38,0,198,0,153,0,146,0,0,0,9,0,82,0,0,0,136,0,50,0,170,0,108,0,75,0,0,0,254,0,149,0,0,0,202,0,230,0,205,0,0,0,253,0,70,0,153,0,68,0,245,0,226,0,212,0,56,0,41,0,0,0,15,0,63,0,63,0,149,0,0,0,157,0,124,0,148,0,70,0,238,0,40,0,26,0,121,0,50,0,103,0,72,0,160,0,122,0,0,0,40,0,147,0,136,0,116,0,0,0,0,0,0,0,172,0,0,0,181,0,0,0,2,0,130,0,139,0,0,0,116,0,0,0,212,0,7,0,0,0,40,0,12,0,197,0,23,0,0,0,126,0,0,0,216,0,0,0,182,0,167,0,0,0,85,0,0,0,0,0,0,0,16,0,97,0,162,0,139,0,0,0,190,0,73,0,116,0,231,0,14,0,114,0,230,0,0,0,0,0,249,0,0,0,13,0,221,0,231,0,22,0,215,0,0,0,179,0,0,0,0,0,140,0,0,0,157,0,0,0,0,0,96,0,0,0,184,0,58,0,202,0,0,0,126,0,237,0,0,0,0,0,21,0,81,0,66,0,72,0,254,0,237,0,0,0,229,0,51,0,29,0,138,0,226,0,0,0,24,0,253,0,189,0,166,0,0,0,0,0,4,0,67,0,207,0,201,0,113,0,0,0,236,0,0,0,211,0,144,0,127,0,146,0,146,0,0,0,216,0,0,0,227,0,19,0,29,0,228,0,23,0,88,0,197,0,0,0,0,0,0,0,178,0,191,0,143,0,0,0,158,0,46,0,162,0,161,0,189,0,118,0,19,0,0,0,86,0,42,0,169,0,163,0,0,0,20,0,49,0,14,0,47,0,8,0,0,0,61,0,155,0,230,0,162,0,49,0,255,0,64,0,49,0,147,0,80,0,125,0,176,0,203,0,105,0,47,0,71,0,0,0,27,0,36,0,0,0,13,0,0,0,0,0,140,0,0,0,205,0,146,0,221,0,0,0,253,0,175,0,0,0,124,0,0,0,211,0,249,0,91,0,202,0,166,0,0,0,146,0,121,0,0,0,217,0,225,0,0,0,0,0,0,0,30,0,188,0,235,0,219,0,139,0,15,0,253,0,0,0,0,0,159,0,37,0,100,0,45,0,210,0,251,0,154,0,0,0,16,0,44,0,170,0,185,0,170,0,93,0,0,0,21,0,0,0,195,0,142,0,135,0,208,0,244,0,231,0,62,0,172,0,172,0,252,0,139,0,16,0,5,0,0,0,192,0,143,0,243,0,7,0,0,0,39,0,0,0,155,0,0,0,223,0,0,0,242,0,115,0,78,0,172,0,0,0,93,0,0,0,237,0,72,0,191,0,0,0,105,0,42,0,155,0,202,0,74,0,5,0,3,0,197,0,151,0,21,0,86,0,120,0,79,0,35,0,6,0,97,0,0,0,149,0,0,0,20,0,171,0,92,0,117,0,114,0,118,0,120,0,105,0,60,0,92,0,0,0,177,0,190,0,184,0,72,0,16,0,149,0,2,0,252,0,29,0,71,0,92,0,210,0,74,0,238,0,0,0,79,0,109,0,126,0,219,0,38,0);
signal scenario_full  : scenario_type := (0,0,247,31,65,31,124,31,68,31,141,31,188,31,111,31,128,31,134,31,134,31,93,31,222,31,122,31,70,31,214,31,95,31,230,31,18,31,18,30,90,31,123,31,123,30,220,31,70,31,70,30,136,31,136,30,172,31,156,31,126,31,126,30,126,29,47,31,254,31,130,31,11,31,44,31,162,31,162,30,70,31,190,31,164,31,57,31,198,31,9,31,247,31,184,31,211,31,62,31,62,30,62,29,138,31,14,31,23,31,89,31,98,31,143,31,143,30,253,31,111,31,215,31,200,31,197,31,197,30,240,31,240,30,23,31,113,31,81,31,81,30,249,31,66,31,66,30,253,31,253,30,76,31,209,31,232,31,232,30,187,31,226,31,150,31,195,31,195,30,214,31,214,30,139,31,223,31,223,30,163,31,95,31,248,31,193,31,239,31,141,31,141,30,126,31,126,30,96,31,96,30,107,31,107,30,107,29,239,31,51,31,45,31,45,30,45,29,45,28,45,27,220,31,12,31,64,31,126,31,232,31,189,31,189,30,189,29,189,28,180,31,243,31,126,31,238,31,184,31,184,30,153,31,242,31,242,30,57,31,43,31,104,31,220,31,140,31,140,30,86,31,101,31,101,30,209,31,209,30,188,31,188,30,83,31,229,31,240,31,69,31,94,31,55,31,22,31,78,31,153,31,102,31,102,30,93,31,245,31,245,30,8,31,199,31,192,31,226,31,226,30,226,29,100,31,96,31,19,31,236,31,236,30,116,31,57,31,199,31,33,31,33,30,33,29,39,31,39,30,39,29,160,31,223,31,223,30,251,31,84,31,69,31,141,31,226,31,226,30,22,31,234,31,168,31,163,31,191,31,12,31,244,31,246,31,143,31,172,31,220,31,90,31,86,31,86,30,28,31,28,30,15,31,251,31,15,31,207,31,219,31,219,30,73,31,100,31,113,31,24,31,24,30,27,31,27,30,51,31,111,31,111,30,167,31,167,30,184,31,184,30,242,31,193,31,52,31,243,31,249,31,123,31,58,31,237,31,73,31,223,31,81,31,11,31,226,31,226,30,23,31,110,31,110,30,110,29,132,31,246,31,128,31,90,31,239,31,176,31,103,31,30,31,30,30,233,31,31,31,57,31,37,31,205,31,62,31,202,31,202,30,202,29,97,31,93,31,67,31,67,30,147,31,147,30,39,31,252,31,252,30,252,29,252,28,129,31,148,31,69,31,141,31,64,31,108,31,246,31,45,31,38,31,198,31,153,31,146,31,146,30,9,31,82,31,82,30,136,31,50,31,170,31,108,31,75,31,75,30,254,31,149,31,149,30,202,31,230,31,205,31,205,30,253,31,70,31,153,31,68,31,245,31,226,31,212,31,56,31,41,31,41,30,15,31,63,31,63,31,149,31,149,30,157,31,124,31,148,31,70,31,238,31,40,31,26,31,121,31,50,31,103,31,72,31,160,31,122,31,122,30,40,31,147,31,136,31,116,31,116,30,116,29,116,28,172,31,172,30,181,31,181,30,2,31,130,31,139,31,139,30,116,31,116,30,212,31,7,31,7,30,40,31,12,31,197,31,23,31,23,30,126,31,126,30,216,31,216,30,182,31,167,31,167,30,85,31,85,30,85,29,85,28,16,31,97,31,162,31,139,31,139,30,190,31,73,31,116,31,231,31,14,31,114,31,230,31,230,30,230,29,249,31,249,30,13,31,221,31,231,31,22,31,215,31,215,30,179,31,179,30,179,29,140,31,140,30,157,31,157,30,157,29,96,31,96,30,184,31,58,31,202,31,202,30,126,31,237,31,237,30,237,29,21,31,81,31,66,31,72,31,254,31,237,31,237,30,229,31,51,31,29,31,138,31,226,31,226,30,24,31,253,31,189,31,166,31,166,30,166,29,4,31,67,31,207,31,201,31,113,31,113,30,236,31,236,30,211,31,144,31,127,31,146,31,146,31,146,30,216,31,216,30,227,31,19,31,29,31,228,31,23,31,88,31,197,31,197,30,197,29,197,28,178,31,191,31,143,31,143,30,158,31,46,31,162,31,161,31,189,31,118,31,19,31,19,30,86,31,42,31,169,31,163,31,163,30,20,31,49,31,14,31,47,31,8,31,8,30,61,31,155,31,230,31,162,31,49,31,255,31,64,31,49,31,147,31,80,31,125,31,176,31,203,31,105,31,47,31,71,31,71,30,27,31,36,31,36,30,13,31,13,30,13,29,140,31,140,30,205,31,146,31,221,31,221,30,253,31,175,31,175,30,124,31,124,30,211,31,249,31,91,31,202,31,166,31,166,30,146,31,121,31,121,30,217,31,225,31,225,30,225,29,225,28,30,31,188,31,235,31,219,31,139,31,15,31,253,31,253,30,253,29,159,31,37,31,100,31,45,31,210,31,251,31,154,31,154,30,16,31,44,31,170,31,185,31,170,31,93,31,93,30,21,31,21,30,195,31,142,31,135,31,208,31,244,31,231,31,62,31,172,31,172,31,252,31,139,31,16,31,5,31,5,30,192,31,143,31,243,31,7,31,7,30,39,31,39,30,155,31,155,30,223,31,223,30,242,31,115,31,78,31,172,31,172,30,93,31,93,30,237,31,72,31,191,31,191,30,105,31,42,31,155,31,202,31,74,31,5,31,3,31,197,31,151,31,21,31,86,31,120,31,79,31,35,31,6,31,97,31,97,30,149,31,149,30,20,31,171,31,92,31,117,31,114,31,118,31,120,31,105,31,60,31,92,31,92,30,177,31,190,31,184,31,72,31,16,31,149,31,2,31,252,31,29,31,71,31,92,31,210,31,74,31,238,31,238,30,79,31,109,31,126,31,219,31,38,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
