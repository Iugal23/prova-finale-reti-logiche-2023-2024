-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 621;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (53,0,33,0,194,0,36,0,42,0,121,0,253,0,186,0,190,0,74,0,141,0,222,0,3,0,81,0,0,0,227,0,0,0,181,0,225,0,205,0,160,0,172,0,72,0,28,0,0,0,210,0,97,0,236,0,0,0,0,0,52,0,157,0,52,0,0,0,0,0,170,0,43,0,159,0,213,0,225,0,219,0,145,0,95,0,58,0,31,0,0,0,0,0,121,0,0,0,207,0,155,0,52,0,0,0,45,0,82,0,151,0,0,0,182,0,248,0,235,0,22,0,0,0,0,0,13,0,10,0,55,0,36,0,200,0,32,0,50,0,0,0,15,0,187,0,179,0,24,0,0,0,36,0,213,0,0,0,157,0,0,0,99,0,233,0,149,0,131,0,0,0,0,0,101,0,0,0,0,0,211,0,250,0,235,0,227,0,164,0,0,0,65,0,0,0,0,0,86,0,39,0,90,0,0,0,34,0,0,0,60,0,194,0,238,0,202,0,145,0,174,0,153,0,122,0,144,0,176,0,171,0,0,0,210,0,202,0,0,0,121,0,87,0,43,0,119,0,239,0,45,0,211,0,48,0,40,0,25,0,48,0,233,0,169,0,156,0,23,0,49,0,72,0,171,0,0,0,32,0,184,0,0,0,0,0,230,0,0,0,0,0,107,0,0,0,14,0,249,0,109,0,20,0,207,0,204,0,0,0,165,0,184,0,68,0,114,0,141,0,179,0,234,0,26,0,194,0,120,0,35,0,0,0,6,0,77,0,24,0,65,0,0,0,114,0,34,0,82,0,45,0,16,0,86,0,93,0,11,0,0,0,116,0,128,0,0,0,0,0,22,0,0,0,162,0,89,0,0,0,0,0,186,0,88,0,173,0,0,0,34,0,0,0,242,0,0,0,0,0,251,0,213,0,196,0,0,0,2,0,0,0,190,0,51,0,59,0,0,0,232,0,0,0,22,0,18,0,57,0,159,0,189,0,95,0,132,0,82,0,0,0,17,0,0,0,88,0,22,0,28,0,132,0,175,0,187,0,226,0,196,0,109,0,100,0,0,0,126,0,186,0,189,0,190,0,0,0,11,0,34,0,138,0,97,0,0,0,196,0,91,0,82,0,105,0,105,0,18,0,120,0,0,0,140,0,19,0,82,0,234,0,30,0,103,0,113,0,76,0,0,0,147,0,0,0,0,0,12,0,204,0,189,0,137,0,0,0,114,0,52,0,0,0,34,0,195,0,10,0,91,0,124,0,0,0,88,0,140,0,0,0,133,0,230,0,115,0,0,0,137,0,0,0,27,0,0,0,5,0,158,0,178,0,214,0,75,0,157,0,45,0,111,0,26,0,34,0,50,0,3,0,132,0,0,0,133,0,122,0,128,0,89,0,181,0,41,0,0,0,0,0,0,0,164,0,191,0,0,0,213,0,55,0,40,0,185,0,254,0,64,0,155,0,91,0,52,0,111,0,251,0,180,0,155,0,99,0,84,0,84,0,127,0,25,0,196,0,0,0,183,0,109,0,171,0,0,0,246,0,73,0,109,0,16,0,38,0,245,0,169,0,0,0,87,0,130,0,206,0,231,0,0,0,80,0,145,0,124,0,0,0,116,0,28,0,168,0,0,0,228,0,0,0,74,0,220,0,29,0,255,0,146,0,117,0,17,0,3,0,120,0,175,0,235,0,123,0,0,0,174,0,184,0,214,0,180,0,145,0,105,0,249,0,146,0,205,0,246,0,51,0,204,0,31,0,22,0,86,0,158,0,231,0,0,0,81,0,129,0,200,0,20,0,162,0,73,0,255,0,76,0,150,0,36,0,0,0,0,0,116,0,189,0,75,0,0,0,179,0,160,0,194,0,224,0,179,0,228,0,0,0,177,0,6,0,217,0,163,0,71,0,119,0,54,0,228,0,0,0,52,0,173,0,61,0,164,0,96,0,0,0,182,0,233,0,101,0,94,0,166,0,0,0,194,0,0,0,0,0,254,0,161,0,225,0,127,0,0,0,157,0,0,0,103,0,0,0,121,0,105,0,207,0,0,0,94,0,0,0,80,0,0,0,252,0,98,0,226,0,48,0,16,0,243,0,89,0,92,0,232,0,117,0,251,0,0,0,210,0,227,0,95,0,0,0,203,0,102,0,250,0,146,0,148,0,141,0,184,0,0,0,123,0,126,0,0,0,203,0,0,0,49,0,165,0,142,0,27,0,234,0,117,0,156,0,85,0,14,0,167,0,6,0,23,0,114,0,98,0,179,0,79,0,134,0,49,0,171,0,97,0,0,0,122,0,160,0,237,0,155,0,43,0,135,0,111,0,69,0,196,0,0,0,157,0,116,0,145,0,0,0,61,0,214,0,65,0,156,0,107,0,124,0,0,0,82,0,236,0,0,0,94,0,237,0,0,0,0,0,17,0,161,0,0,0,0,0,0,0,92,0,59,0,124,0,211,0,0,0,49,0,220,0,48,0,139,0,17,0,102,0,204,0,184,0,212,0,71,0,0,0,0,0,221,0,142,0,110,0,229,0,0,0,62,0,165,0,65,0,0,0,203,0,20,0,0,0,167,0,106,0,0,0,0,0,0,0,50,0,137,0,80,0,121,0,130,0,219,0,185,0,252,0,248,0,95,0,248,0,0,0,210,0,61,0,85,0,204,0,0,0,211,0,0,0,0,0,200,0,116,0,0,0,112,0,154,0,140,0,137,0,133,0,216,0,0,0,0,0,38,0,243,0,42,0,76,0,117,0,48,0,196,0,170,0,234,0,0,0,250,0,250,0,243,0,212,0,103,0,145,0);
signal scenario_full  : scenario_type := (53,31,33,31,194,31,36,31,42,31,121,31,253,31,186,31,190,31,74,31,141,31,222,31,3,31,81,31,81,30,227,31,227,30,181,31,225,31,205,31,160,31,172,31,72,31,28,31,28,30,210,31,97,31,236,31,236,30,236,29,52,31,157,31,52,31,52,30,52,29,170,31,43,31,159,31,213,31,225,31,219,31,145,31,95,31,58,31,31,31,31,30,31,29,121,31,121,30,207,31,155,31,52,31,52,30,45,31,82,31,151,31,151,30,182,31,248,31,235,31,22,31,22,30,22,29,13,31,10,31,55,31,36,31,200,31,32,31,50,31,50,30,15,31,187,31,179,31,24,31,24,30,36,31,213,31,213,30,157,31,157,30,99,31,233,31,149,31,131,31,131,30,131,29,101,31,101,30,101,29,211,31,250,31,235,31,227,31,164,31,164,30,65,31,65,30,65,29,86,31,39,31,90,31,90,30,34,31,34,30,60,31,194,31,238,31,202,31,145,31,174,31,153,31,122,31,144,31,176,31,171,31,171,30,210,31,202,31,202,30,121,31,87,31,43,31,119,31,239,31,45,31,211,31,48,31,40,31,25,31,48,31,233,31,169,31,156,31,23,31,49,31,72,31,171,31,171,30,32,31,184,31,184,30,184,29,230,31,230,30,230,29,107,31,107,30,14,31,249,31,109,31,20,31,207,31,204,31,204,30,165,31,184,31,68,31,114,31,141,31,179,31,234,31,26,31,194,31,120,31,35,31,35,30,6,31,77,31,24,31,65,31,65,30,114,31,34,31,82,31,45,31,16,31,86,31,93,31,11,31,11,30,116,31,128,31,128,30,128,29,22,31,22,30,162,31,89,31,89,30,89,29,186,31,88,31,173,31,173,30,34,31,34,30,242,31,242,30,242,29,251,31,213,31,196,31,196,30,2,31,2,30,190,31,51,31,59,31,59,30,232,31,232,30,22,31,18,31,57,31,159,31,189,31,95,31,132,31,82,31,82,30,17,31,17,30,88,31,22,31,28,31,132,31,175,31,187,31,226,31,196,31,109,31,100,31,100,30,126,31,186,31,189,31,190,31,190,30,11,31,34,31,138,31,97,31,97,30,196,31,91,31,82,31,105,31,105,31,18,31,120,31,120,30,140,31,19,31,82,31,234,31,30,31,103,31,113,31,76,31,76,30,147,31,147,30,147,29,12,31,204,31,189,31,137,31,137,30,114,31,52,31,52,30,34,31,195,31,10,31,91,31,124,31,124,30,88,31,140,31,140,30,133,31,230,31,115,31,115,30,137,31,137,30,27,31,27,30,5,31,158,31,178,31,214,31,75,31,157,31,45,31,111,31,26,31,34,31,50,31,3,31,132,31,132,30,133,31,122,31,128,31,89,31,181,31,41,31,41,30,41,29,41,28,164,31,191,31,191,30,213,31,55,31,40,31,185,31,254,31,64,31,155,31,91,31,52,31,111,31,251,31,180,31,155,31,99,31,84,31,84,31,127,31,25,31,196,31,196,30,183,31,109,31,171,31,171,30,246,31,73,31,109,31,16,31,38,31,245,31,169,31,169,30,87,31,130,31,206,31,231,31,231,30,80,31,145,31,124,31,124,30,116,31,28,31,168,31,168,30,228,31,228,30,74,31,220,31,29,31,255,31,146,31,117,31,17,31,3,31,120,31,175,31,235,31,123,31,123,30,174,31,184,31,214,31,180,31,145,31,105,31,249,31,146,31,205,31,246,31,51,31,204,31,31,31,22,31,86,31,158,31,231,31,231,30,81,31,129,31,200,31,20,31,162,31,73,31,255,31,76,31,150,31,36,31,36,30,36,29,116,31,189,31,75,31,75,30,179,31,160,31,194,31,224,31,179,31,228,31,228,30,177,31,6,31,217,31,163,31,71,31,119,31,54,31,228,31,228,30,52,31,173,31,61,31,164,31,96,31,96,30,182,31,233,31,101,31,94,31,166,31,166,30,194,31,194,30,194,29,254,31,161,31,225,31,127,31,127,30,157,31,157,30,103,31,103,30,121,31,105,31,207,31,207,30,94,31,94,30,80,31,80,30,252,31,98,31,226,31,48,31,16,31,243,31,89,31,92,31,232,31,117,31,251,31,251,30,210,31,227,31,95,31,95,30,203,31,102,31,250,31,146,31,148,31,141,31,184,31,184,30,123,31,126,31,126,30,203,31,203,30,49,31,165,31,142,31,27,31,234,31,117,31,156,31,85,31,14,31,167,31,6,31,23,31,114,31,98,31,179,31,79,31,134,31,49,31,171,31,97,31,97,30,122,31,160,31,237,31,155,31,43,31,135,31,111,31,69,31,196,31,196,30,157,31,116,31,145,31,145,30,61,31,214,31,65,31,156,31,107,31,124,31,124,30,82,31,236,31,236,30,94,31,237,31,237,30,237,29,17,31,161,31,161,30,161,29,161,28,92,31,59,31,124,31,211,31,211,30,49,31,220,31,48,31,139,31,17,31,102,31,204,31,184,31,212,31,71,31,71,30,71,29,221,31,142,31,110,31,229,31,229,30,62,31,165,31,65,31,65,30,203,31,20,31,20,30,167,31,106,31,106,30,106,29,106,28,50,31,137,31,80,31,121,31,130,31,219,31,185,31,252,31,248,31,95,31,248,31,248,30,210,31,61,31,85,31,204,31,204,30,211,31,211,30,211,29,200,31,116,31,116,30,112,31,154,31,140,31,137,31,133,31,216,31,216,30,216,29,38,31,243,31,42,31,76,31,117,31,48,31,196,31,170,31,234,31,234,30,250,31,250,31,243,31,212,31,103,31,145,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
