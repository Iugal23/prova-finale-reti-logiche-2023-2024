-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 187;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (229,0,0,0,194,0,203,0,182,0,0,0,240,0,0,0,9,0,0,0,28,0,2,0,172,0,176,0,0,0,0,0,0,0,118,0,137,0,188,0,96,0,161,0,122,0,208,0,59,0,0,0,92,0,153,0,0,0,78,0,105,0,98,0,40,0,3,0,164,0,186,0,96,0,218,0,186,0,171,0,0,0,0,0,0,0,39,0,166,0,63,0,25,0,63,0,0,0,231,0,0,0,129,0,203,0,158,0,0,0,0,0,250,0,56,0,189,0,145,0,187,0,97,0,150,0,87,0,0,0,61,0,48,0,0,0,191,0,128,0,255,0,145,0,46,0,226,0,201,0,8,0,16,0,169,0,77,0,54,0,74,0,33,0,153,0,132,0,48,0,53,0,227,0,16,0,176,0,0,0,179,0,66,0,0,0,0,0,98,0,0,0,0,0,169,0,104,0,128,0,66,0,38,0,0,0,52,0,205,0,136,0,115,0,74,0,221,0,73,0,0,0,0,0,167,0,183,0,160,0,0,0,38,0,212,0,105,0,0,0,184,0,48,0,89,0,126,0,36,0,39,0,148,0,48,0,175,0,159,0,251,0,192,0,84,0,255,0,21,0,137,0,235,0,215,0,198,0,49,0,65,0,0,0,180,0,0,0,197,0,0,0,143,0,0,0,106,0,42,0,9,0,164,0,19,0,177,0,0,0,24,0,0,0,110,0,0,0,117,0,62,0,18,0,12,0,31,0,181,0,140,0,25,0,50,0,72,0,201,0,186,0,45,0,156,0,111,0,119,0,115,0,0,0,42,0,228,0,152,0,37,0,0,0,0,0,120,0,0,0,77,0,216,0);
signal scenario_full  : scenario_type := (229,31,229,30,194,31,203,31,182,31,182,30,240,31,240,30,9,31,9,30,28,31,2,31,172,31,176,31,176,30,176,29,176,28,118,31,137,31,188,31,96,31,161,31,122,31,208,31,59,31,59,30,92,31,153,31,153,30,78,31,105,31,98,31,40,31,3,31,164,31,186,31,96,31,218,31,186,31,171,31,171,30,171,29,171,28,39,31,166,31,63,31,25,31,63,31,63,30,231,31,231,30,129,31,203,31,158,31,158,30,158,29,250,31,56,31,189,31,145,31,187,31,97,31,150,31,87,31,87,30,61,31,48,31,48,30,191,31,128,31,255,31,145,31,46,31,226,31,201,31,8,31,16,31,169,31,77,31,54,31,74,31,33,31,153,31,132,31,48,31,53,31,227,31,16,31,176,31,176,30,179,31,66,31,66,30,66,29,98,31,98,30,98,29,169,31,104,31,128,31,66,31,38,31,38,30,52,31,205,31,136,31,115,31,74,31,221,31,73,31,73,30,73,29,167,31,183,31,160,31,160,30,38,31,212,31,105,31,105,30,184,31,48,31,89,31,126,31,36,31,39,31,148,31,48,31,175,31,159,31,251,31,192,31,84,31,255,31,21,31,137,31,235,31,215,31,198,31,49,31,65,31,65,30,180,31,180,30,197,31,197,30,143,31,143,30,106,31,42,31,9,31,164,31,19,31,177,31,177,30,24,31,24,30,110,31,110,30,117,31,62,31,18,31,12,31,31,31,181,31,140,31,25,31,50,31,72,31,201,31,186,31,45,31,156,31,111,31,119,31,115,31,115,30,42,31,228,31,152,31,37,31,37,30,37,29,120,31,120,30,77,31,216,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
