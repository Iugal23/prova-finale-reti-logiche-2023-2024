-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 903;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (239,0,152,0,60,0,24,0,36,0,42,0,173,0,144,0,72,0,8,0,101,0,0,0,109,0,179,0,22,0,191,0,0,0,175,0,0,0,86,0,0,0,0,0,9,0,0,0,250,0,98,0,57,0,0,0,0,0,0,0,132,0,170,0,198,0,158,0,154,0,27,0,202,0,0,0,241,0,125,0,107,0,106,0,233,0,185,0,148,0,108,0,39,0,71,0,81,0,209,0,236,0,0,0,212,0,0,0,0,0,0,0,54,0,0,0,21,0,110,0,215,0,0,0,73,0,245,0,239,0,159,0,113,0,243,0,197,0,0,0,10,0,204,0,31,0,182,0,122,0,0,0,250,0,183,0,143,0,0,0,133,0,165,0,75,0,0,0,170,0,134,0,120,0,214,0,0,0,0,0,0,0,243,0,137,0,227,0,44,0,245,0,237,0,187,0,75,0,164,0,40,0,125,0,143,0,27,0,215,0,143,0,31,0,51,0,46,0,8,0,0,0,114,0,151,0,44,0,53,0,182,0,0,0,70,0,0,0,241,0,197,0,239,0,241,0,121,0,40,0,217,0,225,0,255,0,0,0,0,0,223,0,27,0,61,0,60,0,91,0,0,0,155,0,222,0,106,0,49,0,18,0,101,0,125,0,83,0,57,0,101,0,38,0,214,0,87,0,0,0,10,0,193,0,122,0,151,0,108,0,0,0,143,0,81,0,24,0,0,0,0,0,130,0,42,0,0,0,164,0,133,0,0,0,32,0,0,0,16,0,175,0,0,0,202,0,0,0,0,0,119,0,4,0,124,0,110,0,255,0,199,0,0,0,94,0,69,0,120,0,103,0,107,0,252,0,54,0,0,0,230,0,112,0,0,0,106,0,238,0,145,0,57,0,93,0,72,0,0,0,54,0,48,0,0,0,0,0,0,0,168,0,78,0,0,0,225,0,30,0,202,0,204,0,0,0,189,0,0,0,0,0,117,0,96,0,219,0,172,0,0,0,137,0,200,0,46,0,45,0,125,0,23,0,23,0,238,0,169,0,201,0,153,0,51,0,227,0,226,0,81,0,180,0,129,0,0,0,95,0,157,0,255,0,96,0,0,0,170,0,171,0,138,0,0,0,27,0,0,0,191,0,20,0,232,0,205,0,235,0,92,0,18,0,94,0,245,0,36,0,104,0,49,0,204,0,109,0,237,0,232,0,161,0,0,0,211,0,50,0,205,0,200,0,118,0,55,0,36,0,59,0,131,0,0,0,0,0,253,0,0,0,159,0,0,0,172,0,194,0,214,0,0,0,213,0,209,0,0,0,166,0,39,0,48,0,124,0,114,0,4,0,93,0,228,0,242,0,8,0,142,0,27,0,0,0,227,0,139,0,37,0,184,0,145,0,231,0,104,0,81,0,201,0,132,0,0,0,32,0,230,0,242,0,107,0,81,0,181,0,0,0,4,0,244,0,20,0,49,0,43,0,99,0,0,0,143,0,30,0,254,0,98,0,195,0,0,0,216,0,154,0,239,0,0,0,131,0,0,0,0,0,105,0,193,0,86,0,179,0,224,0,17,0,0,0,245,0,199,0,0,0,108,0,48,0,34,0,164,0,22,0,0,0,0,0,71,0,4,0,214,0,0,0,96,0,207,0,0,0,144,0,107,0,37,0,80,0,197,0,0,0,2,0,100,0,0,0,198,0,121,0,7,0,33,0,84,0,21,0,0,0,0,0,0,0,17,0,64,0,181,0,172,0,13,0,230,0,45,0,0,0,0,0,0,0,150,0,230,0,150,0,251,0,9,0,56,0,227,0,1,0,88,0,0,0,179,0,178,0,43,0,44,0,91,0,205,0,26,0,221,0,0,0,186,0,106,0,6,0,90,0,95,0,38,0,25,0,198,0,78,0,22,0,42,0,146,0,14,0,141,0,19,0,224,0,252,0,39,0,58,0,135,0,212,0,251,0,55,0,119,0,106,0,174,0,202,0,24,0,236,0,237,0,254,0,181,0,0,0,0,0,63,0,249,0,189,0,10,0,145,0,224,0,171,0,0,0,106,0,205,0,93,0,210,0,126,0,76,0,52,0,24,0,213,0,90,0,215,0,0,0,0,0,241,0,3,0,44,0,205,0,24,0,251,0,162,0,242,0,198,0,22,0,71,0,118,0,13,0,108,0,207,0,29,0,85,0,77,0,35,0,240,0,100,0,65,0,196,0,109,0,194,0,177,0,0,0,163,0,183,0,154,0,14,0,0,0,105,0,62,0,167,0,101,0,231,0,199,0,88,0,0,0,0,0,0,0,139,0,224,0,188,0,0,0,156,0,141,0,66,0,88,0,8,0,58,0,0,0,162,0,0,0,210,0,211,0,100,0,211,0,12,0,249,0,171,0,13,0,4,0,93,0,84,0,227,0,0,0,62,0,126,0,0,0,205,0,110,0,0,0,0,0,228,0,0,0,186,0,63,0,186,0,129,0,58,0,139,0,42,0,0,0,231,0,68,0,0,0,90,0,113,0,49,0,193,0,0,0,87,0,211,0,145,0,103,0,96,0,175,0,2,0,240,0,16,0,161,0,125,0,0,0,159,0,164,0,38,0,152,0,0,0,173,0,175,0,147,0,60,0,49,0,157,0,241,0,29,0,183,0,0,0,123,0,163,0,175,0,0,0,176,0,45,0,202,0,173,0,249,0,97,0,84,0,149,0,108,0,226,0,114,0,0,0,0,0,35,0,191,0,0,0,65,0,101,0,121,0,88,0,0,0,47,0,98,0,59,0,197,0,0,0,86,0,0,0,84,0,45,0,171,0,235,0,0,0,33,0,0,0,151,0,72,0,47,0,61,0,34,0,107,0,238,0,0,0,255,0,0,0,176,0,57,0,0,0,147,0,120,0,0,0,3,0,0,0,167,0,168,0,154,0,191,0,154,0,0,0,145,0,5,0,192,0,225,0,41,0,145,0,91,0,0,0,204,0,0,0,45,0,119,0,227,0,148,0,0,0,0,0,198,0,197,0,121,0,142,0,140,0,0,0,180,0,215,0,198,0,40,0,254,0,99,0,62,0,0,0,169,0,36,0,228,0,92,0,0,0,0,0,0,0,54,0,132,0,238,0,0,0,0,0,244,0,102,0,0,0,5,0,0,0,132,0,97,0,0,0,204,0,155,0,134,0,189,0,68,0,167,0,204,0,0,0,20,0,96,0,102,0,12,0,126,0,200,0,186,0,160,0,0,0,0,0,0,0,52,0,0,0,216,0,0,0,220,0,199,0,241,0,236,0,19,0,14,0,100,0,0,0,28,0,0,0,75,0,79,0,0,0,77,0,105,0,37,0,238,0,0,0,233,0,0,0,0,0,0,0,216,0,0,0,196,0,161,0,108,0,0,0,174,0,129,0,0,0,148,0,185,0,208,0,120,0,77,0,175,0,250,0,193,0,225,0,27,0,0,0,198,0,203,0,0,0,246,0,196,0,180,0,118,0,0,0,77,0,145,0,205,0,149,0,107,0,220,0,166,0,0,0,130,0,243,0,22,0,0,0,153,0,209,0,131,0,229,0,249,0,13,0,0,0,141,0,71,0,234,0,0,0,98,0,43,0,160,0,0,0,1,0,0,0,208,0,81,0,32,0,253,0,110,0,100,0,94,0,0,0,143,0,240,0,253,0,48,0,239,0,53,0,74,0,110,0,39,0,58,0,142,0,0,0,0,0,61,0,86,0,223,0,236,0,0,0,0,0,0,0,0,0,95,0,243,0,0,0,0,0,159,0,0,0,57,0,120,0,7,0,0,0,17,0,0,0,137,0,251,0,126,0,92,0,108,0,29,0,192,0,221,0,245,0,0,0,232,0,0,0,243,0,39,0,34,0,128,0,0,0,173,0,246,0,177,0,0,0,143,0,79,0,0,0,61,0,0,0,221,0,193,0,36,0,93,0,226,0,0,0,0,0,173,0,48,0,101,0,195,0,240,0,0,0,0,0,88,0,168,0,238,0,64,0,0,0,216,0,234,0,150,0,1,0,0,0,77,0,135,0,236,0,16,0,150,0,218,0,248,0,0,0,0,0,105,0);
signal scenario_full  : scenario_type := (239,31,152,31,60,31,24,31,36,31,42,31,173,31,144,31,72,31,8,31,101,31,101,30,109,31,179,31,22,31,191,31,191,30,175,31,175,30,86,31,86,30,86,29,9,31,9,30,250,31,98,31,57,31,57,30,57,29,57,28,132,31,170,31,198,31,158,31,154,31,27,31,202,31,202,30,241,31,125,31,107,31,106,31,233,31,185,31,148,31,108,31,39,31,71,31,81,31,209,31,236,31,236,30,212,31,212,30,212,29,212,28,54,31,54,30,21,31,110,31,215,31,215,30,73,31,245,31,239,31,159,31,113,31,243,31,197,31,197,30,10,31,204,31,31,31,182,31,122,31,122,30,250,31,183,31,143,31,143,30,133,31,165,31,75,31,75,30,170,31,134,31,120,31,214,31,214,30,214,29,214,28,243,31,137,31,227,31,44,31,245,31,237,31,187,31,75,31,164,31,40,31,125,31,143,31,27,31,215,31,143,31,31,31,51,31,46,31,8,31,8,30,114,31,151,31,44,31,53,31,182,31,182,30,70,31,70,30,241,31,197,31,239,31,241,31,121,31,40,31,217,31,225,31,255,31,255,30,255,29,223,31,27,31,61,31,60,31,91,31,91,30,155,31,222,31,106,31,49,31,18,31,101,31,125,31,83,31,57,31,101,31,38,31,214,31,87,31,87,30,10,31,193,31,122,31,151,31,108,31,108,30,143,31,81,31,24,31,24,30,24,29,130,31,42,31,42,30,164,31,133,31,133,30,32,31,32,30,16,31,175,31,175,30,202,31,202,30,202,29,119,31,4,31,124,31,110,31,255,31,199,31,199,30,94,31,69,31,120,31,103,31,107,31,252,31,54,31,54,30,230,31,112,31,112,30,106,31,238,31,145,31,57,31,93,31,72,31,72,30,54,31,48,31,48,30,48,29,48,28,168,31,78,31,78,30,225,31,30,31,202,31,204,31,204,30,189,31,189,30,189,29,117,31,96,31,219,31,172,31,172,30,137,31,200,31,46,31,45,31,125,31,23,31,23,31,238,31,169,31,201,31,153,31,51,31,227,31,226,31,81,31,180,31,129,31,129,30,95,31,157,31,255,31,96,31,96,30,170,31,171,31,138,31,138,30,27,31,27,30,191,31,20,31,232,31,205,31,235,31,92,31,18,31,94,31,245,31,36,31,104,31,49,31,204,31,109,31,237,31,232,31,161,31,161,30,211,31,50,31,205,31,200,31,118,31,55,31,36,31,59,31,131,31,131,30,131,29,253,31,253,30,159,31,159,30,172,31,194,31,214,31,214,30,213,31,209,31,209,30,166,31,39,31,48,31,124,31,114,31,4,31,93,31,228,31,242,31,8,31,142,31,27,31,27,30,227,31,139,31,37,31,184,31,145,31,231,31,104,31,81,31,201,31,132,31,132,30,32,31,230,31,242,31,107,31,81,31,181,31,181,30,4,31,244,31,20,31,49,31,43,31,99,31,99,30,143,31,30,31,254,31,98,31,195,31,195,30,216,31,154,31,239,31,239,30,131,31,131,30,131,29,105,31,193,31,86,31,179,31,224,31,17,31,17,30,245,31,199,31,199,30,108,31,48,31,34,31,164,31,22,31,22,30,22,29,71,31,4,31,214,31,214,30,96,31,207,31,207,30,144,31,107,31,37,31,80,31,197,31,197,30,2,31,100,31,100,30,198,31,121,31,7,31,33,31,84,31,21,31,21,30,21,29,21,28,17,31,64,31,181,31,172,31,13,31,230,31,45,31,45,30,45,29,45,28,150,31,230,31,150,31,251,31,9,31,56,31,227,31,1,31,88,31,88,30,179,31,178,31,43,31,44,31,91,31,205,31,26,31,221,31,221,30,186,31,106,31,6,31,90,31,95,31,38,31,25,31,198,31,78,31,22,31,42,31,146,31,14,31,141,31,19,31,224,31,252,31,39,31,58,31,135,31,212,31,251,31,55,31,119,31,106,31,174,31,202,31,24,31,236,31,237,31,254,31,181,31,181,30,181,29,63,31,249,31,189,31,10,31,145,31,224,31,171,31,171,30,106,31,205,31,93,31,210,31,126,31,76,31,52,31,24,31,213,31,90,31,215,31,215,30,215,29,241,31,3,31,44,31,205,31,24,31,251,31,162,31,242,31,198,31,22,31,71,31,118,31,13,31,108,31,207,31,29,31,85,31,77,31,35,31,240,31,100,31,65,31,196,31,109,31,194,31,177,31,177,30,163,31,183,31,154,31,14,31,14,30,105,31,62,31,167,31,101,31,231,31,199,31,88,31,88,30,88,29,88,28,139,31,224,31,188,31,188,30,156,31,141,31,66,31,88,31,8,31,58,31,58,30,162,31,162,30,210,31,211,31,100,31,211,31,12,31,249,31,171,31,13,31,4,31,93,31,84,31,227,31,227,30,62,31,126,31,126,30,205,31,110,31,110,30,110,29,228,31,228,30,186,31,63,31,186,31,129,31,58,31,139,31,42,31,42,30,231,31,68,31,68,30,90,31,113,31,49,31,193,31,193,30,87,31,211,31,145,31,103,31,96,31,175,31,2,31,240,31,16,31,161,31,125,31,125,30,159,31,164,31,38,31,152,31,152,30,173,31,175,31,147,31,60,31,49,31,157,31,241,31,29,31,183,31,183,30,123,31,163,31,175,31,175,30,176,31,45,31,202,31,173,31,249,31,97,31,84,31,149,31,108,31,226,31,114,31,114,30,114,29,35,31,191,31,191,30,65,31,101,31,121,31,88,31,88,30,47,31,98,31,59,31,197,31,197,30,86,31,86,30,84,31,45,31,171,31,235,31,235,30,33,31,33,30,151,31,72,31,47,31,61,31,34,31,107,31,238,31,238,30,255,31,255,30,176,31,57,31,57,30,147,31,120,31,120,30,3,31,3,30,167,31,168,31,154,31,191,31,154,31,154,30,145,31,5,31,192,31,225,31,41,31,145,31,91,31,91,30,204,31,204,30,45,31,119,31,227,31,148,31,148,30,148,29,198,31,197,31,121,31,142,31,140,31,140,30,180,31,215,31,198,31,40,31,254,31,99,31,62,31,62,30,169,31,36,31,228,31,92,31,92,30,92,29,92,28,54,31,132,31,238,31,238,30,238,29,244,31,102,31,102,30,5,31,5,30,132,31,97,31,97,30,204,31,155,31,134,31,189,31,68,31,167,31,204,31,204,30,20,31,96,31,102,31,12,31,126,31,200,31,186,31,160,31,160,30,160,29,160,28,52,31,52,30,216,31,216,30,220,31,199,31,241,31,236,31,19,31,14,31,100,31,100,30,28,31,28,30,75,31,79,31,79,30,77,31,105,31,37,31,238,31,238,30,233,31,233,30,233,29,233,28,216,31,216,30,196,31,161,31,108,31,108,30,174,31,129,31,129,30,148,31,185,31,208,31,120,31,77,31,175,31,250,31,193,31,225,31,27,31,27,30,198,31,203,31,203,30,246,31,196,31,180,31,118,31,118,30,77,31,145,31,205,31,149,31,107,31,220,31,166,31,166,30,130,31,243,31,22,31,22,30,153,31,209,31,131,31,229,31,249,31,13,31,13,30,141,31,71,31,234,31,234,30,98,31,43,31,160,31,160,30,1,31,1,30,208,31,81,31,32,31,253,31,110,31,100,31,94,31,94,30,143,31,240,31,253,31,48,31,239,31,53,31,74,31,110,31,39,31,58,31,142,31,142,30,142,29,61,31,86,31,223,31,236,31,236,30,236,29,236,28,236,27,95,31,243,31,243,30,243,29,159,31,159,30,57,31,120,31,7,31,7,30,17,31,17,30,137,31,251,31,126,31,92,31,108,31,29,31,192,31,221,31,245,31,245,30,232,31,232,30,243,31,39,31,34,31,128,31,128,30,173,31,246,31,177,31,177,30,143,31,79,31,79,30,61,31,61,30,221,31,193,31,36,31,93,31,226,31,226,30,226,29,173,31,48,31,101,31,195,31,240,31,240,30,240,29,88,31,168,31,238,31,64,31,64,30,216,31,234,31,150,31,1,31,1,30,77,31,135,31,236,31,16,31,150,31,218,31,248,31,248,30,248,29,105,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
