-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 971;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (52,0,0,0,0,0,242,0,0,0,0,0,227,0,115,0,219,0,51,0,0,0,89,0,126,0,210,0,146,0,23,0,0,0,182,0,96,0,79,0,124,0,0,0,0,0,0,0,0,0,11,0,55,0,0,0,0,0,200,0,24,0,249,0,0,0,243,0,84,0,144,0,0,0,0,0,108,0,85,0,120,0,74,0,227,0,0,0,164,0,59,0,254,0,127,0,123,0,197,0,223,0,23,0,213,0,171,0,77,0,181,0,87,0,19,0,192,0,0,0,0,0,0,0,67,0,188,0,2,0,29,0,0,0,28,0,131,0,109,0,96,0,172,0,227,0,156,0,248,0,58,0,0,0,0,0,192,0,197,0,96,0,166,0,233,0,119,0,200,0,0,0,0,0,2,0,0,0,94,0,240,0,0,0,35,0,41,0,10,0,173,0,242,0,0,0,207,0,0,0,109,0,230,0,0,0,187,0,148,0,92,0,47,0,71,0,125,0,77,0,75,0,0,0,198,0,12,0,121,0,0,0,62,0,107,0,194,0,246,0,0,0,255,0,0,0,195,0,147,0,74,0,221,0,209,0,101,0,247,0,0,0,97,0,236,0,39,0,254,0,239,0,8,0,193,0,212,0,3,0,0,0,12,0,0,0,137,0,49,0,228,0,174,0,2,0,0,0,98,0,154,0,148,0,85,0,38,0,0,0,110,0,147,0,0,0,252,0,133,0,183,0,217,0,53,0,81,0,247,0,0,0,41,0,133,0,246,0,249,0,0,0,0,0,255,0,53,0,0,0,0,0,137,0,0,0,0,0,17,0,42,0,0,0,49,0,58,0,226,0,251,0,26,0,226,0,28,0,1,0,165,0,253,0,0,0,188,0,232,0,203,0,219,0,147,0,191,0,135,0,108,0,10,0,0,0,178,0,109,0,88,0,0,0,130,0,37,0,0,0,102,0,226,0,153,0,0,0,126,0,42,0,0,0,0,0,34,0,20,0,0,0,0,0,68,0,110,0,85,0,0,0,152,0,52,0,151,0,0,0,201,0,190,0,25,0,239,0,224,0,34,0,0,0,0,0,172,0,197,0,56,0,227,0,217,0,0,0,155,0,151,0,127,0,188,0,0,0,0,0,240,0,181,0,33,0,154,0,0,0,16,0,17,0,176,0,127,0,0,0,183,0,123,0,170,0,36,0,151,0,0,0,241,0,63,0,38,0,230,0,0,0,0,0,0,0,69,0,123,0,7,0,1,0,242,0,24,0,17,0,60,0,101,0,90,0,145,0,254,0,200,0,39,0,126,0,163,0,192,0,50,0,10,0,200,0,89,0,67,0,180,0,218,0,245,0,114,0,142,0,22,0,44,0,0,0,0,0,81,0,173,0,4,0,43,0,36,0,0,0,158,0,0,0,0,0,233,0,218,0,253,0,190,0,220,0,214,0,148,0,120,0,149,0,208,0,19,0,17,0,0,0,43,0,74,0,240,0,103,0,41,0,218,0,230,0,196,0,155,0,209,0,212,0,100,0,0,0,138,0,105,0,0,0,0,0,0,0,4,0,137,0,115,0,176,0,63,0,80,0,2,0,132,0,0,0,245,0,169,0,143,0,219,0,233,0,149,0,17,0,0,0,119,0,158,0,215,0,163,0,94,0,134,0,157,0,108,0,20,0,27,0,254,0,207,0,71,0,0,0,255,0,110,0,35,0,226,0,0,0,53,0,31,0,137,0,217,0,197,0,250,0,0,0,87,0,243,0,0,0,26,0,137,0,215,0,169,0,137,0,24,0,0,0,72,0,106,0,86,0,240,0,224,0,141,0,212,0,36,0,48,0,0,0,46,0,141,0,251,0,151,0,0,0,127,0,179,0,147,0,0,0,4,0,178,0,134,0,71,0,140,0,0,0,0,0,61,0,168,0,0,0,82,0,27,0,0,0,199,0,23,0,197,0,196,0,119,0,173,0,102,0,87,0,83,0,215,0,175,0,135,0,142,0,191,0,165,0,0,0,0,0,175,0,220,0,0,0,89,0,222,0,67,0,100,0,0,0,0,0,16,0,8,0,43,0,40,0,0,0,122,0,5,0,87,0,67,0,187,0,255,0,37,0,119,0,8,0,183,0,10,0,126,0,157,0,0,0,225,0,8,0,0,0,176,0,73,0,0,0,180,0,218,0,0,0,43,0,148,0,78,0,3,0,131,0,37,0,194,0,0,0,22,0,0,0,166,0,120,0,1,0,0,0,107,0,214,0,136,0,84,0,75,0,0,0,245,0,194,0,55,0,0,0,170,0,217,0,201,0,0,0,237,0,133,0,81,0,0,0,0,0,77,0,0,0,106,0,77,0,0,0,216,0,107,0,135,0,38,0,113,0,196,0,112,0,0,0,40,0,0,0,203,0,190,0,214,0,212,0,20,0,32,0,0,0,63,0,0,0,0,0,236,0,0,0,99,0,148,0,8,0,0,0,99,0,249,0,138,0,241,0,60,0,113,0,0,0,250,0,54,0,14,0,55,0,0,0,174,0,1,0,239,0,0,0,0,0,141,0,120,0,238,0,112,0,109,0,96,0,186,0,12,0,84,0,241,0,244,0,64,0,37,0,98,0,0,0,149,0,214,0,108,0,0,0,109,0,94,0,165,0,13,0,0,0,101,0,136,0,72,0,0,0,184,0,148,0,127,0,176,0,0,0,59,0,38,0,0,0,11,0,213,0,174,0,127,0,39,0,0,0,70,0,200,0,62,0,70,0,82,0,127,0,6,0,0,0,130,0,241,0,0,0,121,0,219,0,0,0,170,0,0,0,0,0,129,0,92,0,171,0,0,0,126,0,124,0,151,0,0,0,0,0,152,0,186,0,161,0,81,0,0,0,231,0,82,0,20,0,15,0,165,0,237,0,0,0,171,0,0,0,123,0,35,0,149,0,247,0,235,0,255,0,202,0,182,0,239,0,0,0,71,0,0,0,119,0,217,0,21,0,159,0,17,0,0,0,68,0,0,0,60,0,145,0,146,0,148,0,33,0,0,0,22,0,6,0,0,0,111,0,114,0,138,0,101,0,194,0,73,0,0,0,60,0,122,0,0,0,205,0,198,0,31,0,63,0,213,0,91,0,163,0,74,0,228,0,111,0,72,0,0,0,0,0,0,0,74,0,45,0,104,0,191,0,85,0,161,0,102,0,137,0,198,0,116,0,0,0,195,0,167,0,144,0,241,0,212,0,0,0,145,0,152,0,219,0,158,0,95,0,23,0,220,0,211,0,0,0,111,0,0,0,207,0,200,0,224,0,112,0,41,0,157,0,196,0,2,0,77,0,178,0,248,0,0,0,0,0,255,0,46,0,114,0,0,0,180,0,61,0,176,0,106,0,249,0,225,0,72,0,84,0,0,0,0,0,166,0,43,0,0,0,160,0,233,0,22,0,140,0,102,0,122,0,0,0,97,0,10,0,216,0,148,0,27,0,86,0,66,0,103,0,115,0,41,0,0,0,0,0,167,0,67,0,33,0,20,0,0,0,0,0,77,0,0,0,213,0,137,0,239,0,42,0,100,0,50,0,0,0,142,0,59,0,57,0,102,0,208,0,121,0,103,0,144,0,140,0,0,0,128,0,188,0,12,0,76,0,39,0,76,0,215,0,156,0,168,0,197,0,231,0,44,0,0,0,182,0,0,0,9,0,0,0,92,0,170,0,202,0,159,0,223,0,85,0,0,0,0,0,229,0,151,0,14,0,103,0,129,0,99,0,73,0,74,0,199,0,109,0,42,0,191,0,133,0,0,0,55,0,156,0,0,0,0,0,79,0,135,0,52,0,70,0,0,0,134,0,79,0,207,0,111,0,186,0,0,0,9,0,128,0,0,0,26,0,205,0,12,0,114,0,124,0,132,0,0,0,0,0,117,0,124,0,22,0,236,0,135,0,22,0,242,0,0,0,0,0,146,0,0,0,0,0,0,0,13,0,64,0,219,0,0,0,87,0,145,0,223,0,167,0,126,0,108,0,252,0,46,0,168,0,112,0,0,0,0,0,124,0,70,0,191,0,103,0,249,0,88,0,38,0,80,0,24,0,237,0,149,0,20,0,163,0,62,0,13,0,252,0,165,0,0,0,113,0,176,0,20,0,107,0,128,0,0,0,22,0,75,0,230,0,120,0,164,0,0,0,105,0,122,0,0,0,203,0,153,0,0,0,0,0,175,0,152,0,195,0,68,0,135,0,237,0,0,0,100,0,90,0,69,0,145,0,0,0,221,0,251,0,243,0,37,0,17,0,0,0,1,0,0,0,200,0,0,0,206,0,51,0,226,0,59,0,132,0,167,0,122,0,0,0,104,0,59,0,195,0,183,0,58,0,0,0,217,0,166,0,69,0);
signal scenario_full  : scenario_type := (52,31,52,30,52,29,242,31,242,30,242,29,227,31,115,31,219,31,51,31,51,30,89,31,126,31,210,31,146,31,23,31,23,30,182,31,96,31,79,31,124,31,124,30,124,29,124,28,124,27,11,31,55,31,55,30,55,29,200,31,24,31,249,31,249,30,243,31,84,31,144,31,144,30,144,29,108,31,85,31,120,31,74,31,227,31,227,30,164,31,59,31,254,31,127,31,123,31,197,31,223,31,23,31,213,31,171,31,77,31,181,31,87,31,19,31,192,31,192,30,192,29,192,28,67,31,188,31,2,31,29,31,29,30,28,31,131,31,109,31,96,31,172,31,227,31,156,31,248,31,58,31,58,30,58,29,192,31,197,31,96,31,166,31,233,31,119,31,200,31,200,30,200,29,2,31,2,30,94,31,240,31,240,30,35,31,41,31,10,31,173,31,242,31,242,30,207,31,207,30,109,31,230,31,230,30,187,31,148,31,92,31,47,31,71,31,125,31,77,31,75,31,75,30,198,31,12,31,121,31,121,30,62,31,107,31,194,31,246,31,246,30,255,31,255,30,195,31,147,31,74,31,221,31,209,31,101,31,247,31,247,30,97,31,236,31,39,31,254,31,239,31,8,31,193,31,212,31,3,31,3,30,12,31,12,30,137,31,49,31,228,31,174,31,2,31,2,30,98,31,154,31,148,31,85,31,38,31,38,30,110,31,147,31,147,30,252,31,133,31,183,31,217,31,53,31,81,31,247,31,247,30,41,31,133,31,246,31,249,31,249,30,249,29,255,31,53,31,53,30,53,29,137,31,137,30,137,29,17,31,42,31,42,30,49,31,58,31,226,31,251,31,26,31,226,31,28,31,1,31,165,31,253,31,253,30,188,31,232,31,203,31,219,31,147,31,191,31,135,31,108,31,10,31,10,30,178,31,109,31,88,31,88,30,130,31,37,31,37,30,102,31,226,31,153,31,153,30,126,31,42,31,42,30,42,29,34,31,20,31,20,30,20,29,68,31,110,31,85,31,85,30,152,31,52,31,151,31,151,30,201,31,190,31,25,31,239,31,224,31,34,31,34,30,34,29,172,31,197,31,56,31,227,31,217,31,217,30,155,31,151,31,127,31,188,31,188,30,188,29,240,31,181,31,33,31,154,31,154,30,16,31,17,31,176,31,127,31,127,30,183,31,123,31,170,31,36,31,151,31,151,30,241,31,63,31,38,31,230,31,230,30,230,29,230,28,69,31,123,31,7,31,1,31,242,31,24,31,17,31,60,31,101,31,90,31,145,31,254,31,200,31,39,31,126,31,163,31,192,31,50,31,10,31,200,31,89,31,67,31,180,31,218,31,245,31,114,31,142,31,22,31,44,31,44,30,44,29,81,31,173,31,4,31,43,31,36,31,36,30,158,31,158,30,158,29,233,31,218,31,253,31,190,31,220,31,214,31,148,31,120,31,149,31,208,31,19,31,17,31,17,30,43,31,74,31,240,31,103,31,41,31,218,31,230,31,196,31,155,31,209,31,212,31,100,31,100,30,138,31,105,31,105,30,105,29,105,28,4,31,137,31,115,31,176,31,63,31,80,31,2,31,132,31,132,30,245,31,169,31,143,31,219,31,233,31,149,31,17,31,17,30,119,31,158,31,215,31,163,31,94,31,134,31,157,31,108,31,20,31,27,31,254,31,207,31,71,31,71,30,255,31,110,31,35,31,226,31,226,30,53,31,31,31,137,31,217,31,197,31,250,31,250,30,87,31,243,31,243,30,26,31,137,31,215,31,169,31,137,31,24,31,24,30,72,31,106,31,86,31,240,31,224,31,141,31,212,31,36,31,48,31,48,30,46,31,141,31,251,31,151,31,151,30,127,31,179,31,147,31,147,30,4,31,178,31,134,31,71,31,140,31,140,30,140,29,61,31,168,31,168,30,82,31,27,31,27,30,199,31,23,31,197,31,196,31,119,31,173,31,102,31,87,31,83,31,215,31,175,31,135,31,142,31,191,31,165,31,165,30,165,29,175,31,220,31,220,30,89,31,222,31,67,31,100,31,100,30,100,29,16,31,8,31,43,31,40,31,40,30,122,31,5,31,87,31,67,31,187,31,255,31,37,31,119,31,8,31,183,31,10,31,126,31,157,31,157,30,225,31,8,31,8,30,176,31,73,31,73,30,180,31,218,31,218,30,43,31,148,31,78,31,3,31,131,31,37,31,194,31,194,30,22,31,22,30,166,31,120,31,1,31,1,30,107,31,214,31,136,31,84,31,75,31,75,30,245,31,194,31,55,31,55,30,170,31,217,31,201,31,201,30,237,31,133,31,81,31,81,30,81,29,77,31,77,30,106,31,77,31,77,30,216,31,107,31,135,31,38,31,113,31,196,31,112,31,112,30,40,31,40,30,203,31,190,31,214,31,212,31,20,31,32,31,32,30,63,31,63,30,63,29,236,31,236,30,99,31,148,31,8,31,8,30,99,31,249,31,138,31,241,31,60,31,113,31,113,30,250,31,54,31,14,31,55,31,55,30,174,31,1,31,239,31,239,30,239,29,141,31,120,31,238,31,112,31,109,31,96,31,186,31,12,31,84,31,241,31,244,31,64,31,37,31,98,31,98,30,149,31,214,31,108,31,108,30,109,31,94,31,165,31,13,31,13,30,101,31,136,31,72,31,72,30,184,31,148,31,127,31,176,31,176,30,59,31,38,31,38,30,11,31,213,31,174,31,127,31,39,31,39,30,70,31,200,31,62,31,70,31,82,31,127,31,6,31,6,30,130,31,241,31,241,30,121,31,219,31,219,30,170,31,170,30,170,29,129,31,92,31,171,31,171,30,126,31,124,31,151,31,151,30,151,29,152,31,186,31,161,31,81,31,81,30,231,31,82,31,20,31,15,31,165,31,237,31,237,30,171,31,171,30,123,31,35,31,149,31,247,31,235,31,255,31,202,31,182,31,239,31,239,30,71,31,71,30,119,31,217,31,21,31,159,31,17,31,17,30,68,31,68,30,60,31,145,31,146,31,148,31,33,31,33,30,22,31,6,31,6,30,111,31,114,31,138,31,101,31,194,31,73,31,73,30,60,31,122,31,122,30,205,31,198,31,31,31,63,31,213,31,91,31,163,31,74,31,228,31,111,31,72,31,72,30,72,29,72,28,74,31,45,31,104,31,191,31,85,31,161,31,102,31,137,31,198,31,116,31,116,30,195,31,167,31,144,31,241,31,212,31,212,30,145,31,152,31,219,31,158,31,95,31,23,31,220,31,211,31,211,30,111,31,111,30,207,31,200,31,224,31,112,31,41,31,157,31,196,31,2,31,77,31,178,31,248,31,248,30,248,29,255,31,46,31,114,31,114,30,180,31,61,31,176,31,106,31,249,31,225,31,72,31,84,31,84,30,84,29,166,31,43,31,43,30,160,31,233,31,22,31,140,31,102,31,122,31,122,30,97,31,10,31,216,31,148,31,27,31,86,31,66,31,103,31,115,31,41,31,41,30,41,29,167,31,67,31,33,31,20,31,20,30,20,29,77,31,77,30,213,31,137,31,239,31,42,31,100,31,50,31,50,30,142,31,59,31,57,31,102,31,208,31,121,31,103,31,144,31,140,31,140,30,128,31,188,31,12,31,76,31,39,31,76,31,215,31,156,31,168,31,197,31,231,31,44,31,44,30,182,31,182,30,9,31,9,30,92,31,170,31,202,31,159,31,223,31,85,31,85,30,85,29,229,31,151,31,14,31,103,31,129,31,99,31,73,31,74,31,199,31,109,31,42,31,191,31,133,31,133,30,55,31,156,31,156,30,156,29,79,31,135,31,52,31,70,31,70,30,134,31,79,31,207,31,111,31,186,31,186,30,9,31,128,31,128,30,26,31,205,31,12,31,114,31,124,31,132,31,132,30,132,29,117,31,124,31,22,31,236,31,135,31,22,31,242,31,242,30,242,29,146,31,146,30,146,29,146,28,13,31,64,31,219,31,219,30,87,31,145,31,223,31,167,31,126,31,108,31,252,31,46,31,168,31,112,31,112,30,112,29,124,31,70,31,191,31,103,31,249,31,88,31,38,31,80,31,24,31,237,31,149,31,20,31,163,31,62,31,13,31,252,31,165,31,165,30,113,31,176,31,20,31,107,31,128,31,128,30,22,31,75,31,230,31,120,31,164,31,164,30,105,31,122,31,122,30,203,31,153,31,153,30,153,29,175,31,152,31,195,31,68,31,135,31,237,31,237,30,100,31,90,31,69,31,145,31,145,30,221,31,251,31,243,31,37,31,17,31,17,30,1,31,1,30,200,31,200,30,206,31,51,31,226,31,59,31,132,31,167,31,122,31,122,30,104,31,59,31,195,31,183,31,58,31,58,30,217,31,166,31,69,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
