-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 528;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (168,0,200,0,250,0,0,0,38,0,92,0,196,0,225,0,84,0,0,0,199,0,93,0,173,0,0,0,0,0,186,0,0,0,0,0,224,0,0,0,86,0,169,0,0,0,197,0,26,0,127,0,234,0,162,0,80,0,12,0,113,0,0,0,0,0,101,0,0,0,0,0,173,0,89,0,0,0,0,0,61,0,183,0,1,0,52,0,167,0,0,0,216,0,235,0,11,0,0,0,104,0,66,0,74,0,66,0,146,0,101,0,0,0,242,0,194,0,0,0,219,0,163,0,61,0,10,0,157,0,0,0,137,0,212,0,0,0,106,0,196,0,198,0,146,0,167,0,176,0,20,0,164,0,207,0,0,0,211,0,95,0,188,0,253,0,50,0,203,0,61,0,76,0,10,0,22,0,8,0,180,0,175,0,0,0,75,0,182,0,215,0,144,0,68,0,3,0,112,0,34,0,253,0,12,0,25,0,95,0,149,0,0,0,6,0,133,0,99,0,0,0,155,0,0,0,186,0,0,0,0,0,21,0,91,0,196,0,205,0,41,0,57,0,38,0,66,0,252,0,226,0,198,0,129,0,195,0,162,0,0,0,235,0,202,0,86,0,53,0,124,0,7,0,0,0,51,0,0,0,111,0,121,0,236,0,0,0,238,0,237,0,0,0,176,0,0,0,75,0,170,0,30,0,162,0,130,0,0,0,176,0,152,0,0,0,100,0,42,0,11,0,164,0,200,0,105,0,99,0,0,0,208,0,210,0,147,0,11,0,78,0,0,0,132,0,0,0,177,0,0,0,168,0,98,0,243,0,134,0,219,0,141,0,79,0,200,0,19,0,45,0,16,0,0,0,122,0,0,0,251,0,76,0,168,0,210,0,164,0,209,0,0,0,168,0,234,0,39,0,31,0,167,0,193,0,43,0,0,0,0,0,39,0,100,0,229,0,107,0,124,0,88,0,0,0,168,0,34,0,227,0,138,0,114,0,163,0,21,0,0,0,13,0,205,0,0,0,2,0,106,0,166,0,101,0,0,0,78,0,124,0,0,0,1,0,228,0,114,0,138,0,0,0,0,0,185,0,121,0,0,0,232,0,78,0,100,0,68,0,0,0,47,0,74,0,112,0,220,0,205,0,249,0,0,0,0,0,61,0,62,0,98,0,54,0,2,0,188,0,202,0,59,0,174,0,0,0,216,0,23,0,138,0,0,0,177,0,0,0,45,0,203,0,19,0,148,0,163,0,0,0,0,0,211,0,232,0,109,0,149,0,230,0,0,0,160,0,159,0,119,0,233,0,161,0,0,0,157,0,206,0,255,0,0,0,226,0,5,0,125,0,151,0,246,0,20,0,217,0,235,0,0,0,0,0,243,0,14,0,138,0,195,0,184,0,0,0,0,0,178,0,93,0,182,0,73,0,184,0,152,0,176,0,22,0,221,0,180,0,0,0,0,0,0,0,254,0,240,0,0,0,81,0,65,0,192,0,89,0,44,0,156,0,248,0,1,0,127,0,0,0,194,0,242,0,0,0,207,0,0,0,0,0,184,0,108,0,95,0,128,0,0,0,55,0,119,0,0,0,199,0,223,0,240,0,0,0,94,0,82,0,209,0,72,0,70,0,20,0,228,0,67,0,57,0,0,0,140,0,193,0,172,0,120,0,191,0,187,0,249,0,0,0,222,0,207,0,56,0,0,0,28,0,0,0,93,0,0,0,14,0,0,0,0,0,52,0,150,0,0,0,114,0,80,0,0,0,0,0,35,0,103,0,0,0,137,0,87,0,142,0,39,0,43,0,167,0,0,0,185,0,166,0,0,0,195,0,80,0,47,0,99,0,197,0,0,0,136,0,218,0,174,0,15,0,0,0,140,0,3,0,0,0,255,0,173,0,71,0,47,0,230,0,0,0,103,0,215,0,209,0,176,0,153,0,116,0,204,0,0,0,73,0,0,0,235,0,19,0,0,0,254,0,200,0,56,0,37,0,0,0,53,0,39,0,0,0,93,0,168,0,20,0,228,0,110,0,132,0,126,0,210,0,198,0,242,0,116,0,48,0,84,0,79,0,0,0,221,0,196,0,96,0,240,0,11,0,0,0,246,0,0,0,0,0,60,0,106,0,132,0,136,0,0,0,212,0,0,0,62,0,72,0,5,0,0,0,68,0,0,0,0,0,157,0,45,0,34,0,42,0,142,0,133,0,21,0,0,0,2,0,33,0,0,0,0,0,0,0,0,0,0,0,109,0,42,0,0,0,0,0,12,0,0,0,165,0,0,0,217,0,62,0,50,0,167,0,217,0,241,0,57,0,1,0,195,0,63,0,0,0,98,0,222,0,217,0,33,0,3,0,240,0,30,0,0,0,0,0,197,0,102,0,106,0);
signal scenario_full  : scenario_type := (168,31,200,31,250,31,250,30,38,31,92,31,196,31,225,31,84,31,84,30,199,31,93,31,173,31,173,30,173,29,186,31,186,30,186,29,224,31,224,30,86,31,169,31,169,30,197,31,26,31,127,31,234,31,162,31,80,31,12,31,113,31,113,30,113,29,101,31,101,30,101,29,173,31,89,31,89,30,89,29,61,31,183,31,1,31,52,31,167,31,167,30,216,31,235,31,11,31,11,30,104,31,66,31,74,31,66,31,146,31,101,31,101,30,242,31,194,31,194,30,219,31,163,31,61,31,10,31,157,31,157,30,137,31,212,31,212,30,106,31,196,31,198,31,146,31,167,31,176,31,20,31,164,31,207,31,207,30,211,31,95,31,188,31,253,31,50,31,203,31,61,31,76,31,10,31,22,31,8,31,180,31,175,31,175,30,75,31,182,31,215,31,144,31,68,31,3,31,112,31,34,31,253,31,12,31,25,31,95,31,149,31,149,30,6,31,133,31,99,31,99,30,155,31,155,30,186,31,186,30,186,29,21,31,91,31,196,31,205,31,41,31,57,31,38,31,66,31,252,31,226,31,198,31,129,31,195,31,162,31,162,30,235,31,202,31,86,31,53,31,124,31,7,31,7,30,51,31,51,30,111,31,121,31,236,31,236,30,238,31,237,31,237,30,176,31,176,30,75,31,170,31,30,31,162,31,130,31,130,30,176,31,152,31,152,30,100,31,42,31,11,31,164,31,200,31,105,31,99,31,99,30,208,31,210,31,147,31,11,31,78,31,78,30,132,31,132,30,177,31,177,30,168,31,98,31,243,31,134,31,219,31,141,31,79,31,200,31,19,31,45,31,16,31,16,30,122,31,122,30,251,31,76,31,168,31,210,31,164,31,209,31,209,30,168,31,234,31,39,31,31,31,167,31,193,31,43,31,43,30,43,29,39,31,100,31,229,31,107,31,124,31,88,31,88,30,168,31,34,31,227,31,138,31,114,31,163,31,21,31,21,30,13,31,205,31,205,30,2,31,106,31,166,31,101,31,101,30,78,31,124,31,124,30,1,31,228,31,114,31,138,31,138,30,138,29,185,31,121,31,121,30,232,31,78,31,100,31,68,31,68,30,47,31,74,31,112,31,220,31,205,31,249,31,249,30,249,29,61,31,62,31,98,31,54,31,2,31,188,31,202,31,59,31,174,31,174,30,216,31,23,31,138,31,138,30,177,31,177,30,45,31,203,31,19,31,148,31,163,31,163,30,163,29,211,31,232,31,109,31,149,31,230,31,230,30,160,31,159,31,119,31,233,31,161,31,161,30,157,31,206,31,255,31,255,30,226,31,5,31,125,31,151,31,246,31,20,31,217,31,235,31,235,30,235,29,243,31,14,31,138,31,195,31,184,31,184,30,184,29,178,31,93,31,182,31,73,31,184,31,152,31,176,31,22,31,221,31,180,31,180,30,180,29,180,28,254,31,240,31,240,30,81,31,65,31,192,31,89,31,44,31,156,31,248,31,1,31,127,31,127,30,194,31,242,31,242,30,207,31,207,30,207,29,184,31,108,31,95,31,128,31,128,30,55,31,119,31,119,30,199,31,223,31,240,31,240,30,94,31,82,31,209,31,72,31,70,31,20,31,228,31,67,31,57,31,57,30,140,31,193,31,172,31,120,31,191,31,187,31,249,31,249,30,222,31,207,31,56,31,56,30,28,31,28,30,93,31,93,30,14,31,14,30,14,29,52,31,150,31,150,30,114,31,80,31,80,30,80,29,35,31,103,31,103,30,137,31,87,31,142,31,39,31,43,31,167,31,167,30,185,31,166,31,166,30,195,31,80,31,47,31,99,31,197,31,197,30,136,31,218,31,174,31,15,31,15,30,140,31,3,31,3,30,255,31,173,31,71,31,47,31,230,31,230,30,103,31,215,31,209,31,176,31,153,31,116,31,204,31,204,30,73,31,73,30,235,31,19,31,19,30,254,31,200,31,56,31,37,31,37,30,53,31,39,31,39,30,93,31,168,31,20,31,228,31,110,31,132,31,126,31,210,31,198,31,242,31,116,31,48,31,84,31,79,31,79,30,221,31,196,31,96,31,240,31,11,31,11,30,246,31,246,30,246,29,60,31,106,31,132,31,136,31,136,30,212,31,212,30,62,31,72,31,5,31,5,30,68,31,68,30,68,29,157,31,45,31,34,31,42,31,142,31,133,31,21,31,21,30,2,31,33,31,33,30,33,29,33,28,33,27,33,26,109,31,42,31,42,30,42,29,12,31,12,30,165,31,165,30,217,31,62,31,50,31,167,31,217,31,241,31,57,31,1,31,195,31,63,31,63,30,98,31,222,31,217,31,33,31,3,31,240,31,30,31,30,30,30,29,197,31,102,31,106,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
