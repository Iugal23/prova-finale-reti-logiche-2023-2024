-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 352;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (143,0,40,0,41,0,217,0,179,0,46,0,78,0,92,0,129,0,147,0,58,0,123,0,240,0,201,0,0,0,230,0,0,0,0,0,42,0,0,0,230,0,166,0,144,0,19,0,93,0,0,0,135,0,18,0,191,0,146,0,0,0,250,0,51,0,115,0,189,0,165,0,164,0,0,0,179,0,227,0,15,0,157,0,89,0,0,0,0,0,167,0,183,0,0,0,194,0,0,0,22,0,150,0,0,0,58,0,140,0,145,0,44,0,62,0,187,0,239,0,38,0,0,0,184,0,44,0,0,0,0,0,105,0,239,0,0,0,20,0,27,0,237,0,0,0,212,0,0,0,0,0,201,0,37,0,97,0,22,0,221,0,102,0,42,0,47,0,250,0,188,0,57,0,188,0,51,0,213,0,152,0,106,0,151,0,67,0,242,0,0,0,16,0,15,0,0,0,57,0,0,0,222,0,100,0,169,0,142,0,247,0,209,0,159,0,166,0,0,0,121,0,103,0,0,0,0,0,54,0,0,0,205,0,29,0,0,0,114,0,0,0,0,0,101,0,132,0,32,0,243,0,246,0,0,0,243,0,27,0,75,0,34,0,141,0,17,0,0,0,0,0,70,0,105,0,66,0,189,0,43,0,238,0,124,0,0,0,182,0,157,0,225,0,6,0,110,0,0,0,38,0,122,0,0,0,0,0,0,0,48,0,0,0,185,0,181,0,88,0,75,0,219,0,213,0,96,0,127,0,170,0,110,0,3,0,95,0,27,0,0,0,239,0,223,0,192,0,251,0,119,0,0,0,129,0,250,0,187,0,94,0,0,0,0,0,118,0,0,0,45,0,10,0,0,0,0,0,128,0,64,0,41,0,61,0,106,0,153,0,150,0,223,0,101,0,166,0,243,0,0,0,88,0,111,0,198,0,1,0,158,0,37,0,169,0,191,0,0,0,0,0,190,0,95,0,194,0,38,0,167,0,243,0,71,0,174,0,0,0,2,0,195,0,93,0,141,0,113,0,229,0,219,0,197,0,214,0,0,0,230,0,229,0,144,0,101,0,221,0,248,0,80,0,12,0,144,0,137,0,176,0,177,0,179,0,88,0,98,0,32,0,231,0,248,0,0,0,0,0,0,0,154,0,0,0,150,0,0,0,116,0,18,0,245,0,0,0,232,0,119,0,76,0,183,0,67,0,156,0,230,0,251,0,0,0,16,0,0,0,143,0,220,0,220,0,157,0,150,0,23,0,0,0,93,0,109,0,0,0,5,0,178,0,252,0,40,0,228,0,141,0,107,0,35,0,252,0,141,0,34,0,102,0,163,0,76,0,33,0,0,0,71,0,126,0,0,0,0,0,214,0,0,0,212,0,176,0,10,0,150,0,6,0,47,0,141,0,12,0,52,0,92,0,214,0,85,0,232,0,133,0,163,0,192,0,239,0,201,0,181,0,0,0,80,0,78,0,0,0,61,0,38,0,0,0,10,0,51,0,232,0,32,0,91,0,109,0,205,0,0,0,24,0,163,0,144,0,239,0,215,0,136,0,21,0,11,0,30,0,152,0,96,0,54,0,200,0,46,0,45,0,10,0);
signal scenario_full  : scenario_type := (143,31,40,31,41,31,217,31,179,31,46,31,78,31,92,31,129,31,147,31,58,31,123,31,240,31,201,31,201,30,230,31,230,30,230,29,42,31,42,30,230,31,166,31,144,31,19,31,93,31,93,30,135,31,18,31,191,31,146,31,146,30,250,31,51,31,115,31,189,31,165,31,164,31,164,30,179,31,227,31,15,31,157,31,89,31,89,30,89,29,167,31,183,31,183,30,194,31,194,30,22,31,150,31,150,30,58,31,140,31,145,31,44,31,62,31,187,31,239,31,38,31,38,30,184,31,44,31,44,30,44,29,105,31,239,31,239,30,20,31,27,31,237,31,237,30,212,31,212,30,212,29,201,31,37,31,97,31,22,31,221,31,102,31,42,31,47,31,250,31,188,31,57,31,188,31,51,31,213,31,152,31,106,31,151,31,67,31,242,31,242,30,16,31,15,31,15,30,57,31,57,30,222,31,100,31,169,31,142,31,247,31,209,31,159,31,166,31,166,30,121,31,103,31,103,30,103,29,54,31,54,30,205,31,29,31,29,30,114,31,114,30,114,29,101,31,132,31,32,31,243,31,246,31,246,30,243,31,27,31,75,31,34,31,141,31,17,31,17,30,17,29,70,31,105,31,66,31,189,31,43,31,238,31,124,31,124,30,182,31,157,31,225,31,6,31,110,31,110,30,38,31,122,31,122,30,122,29,122,28,48,31,48,30,185,31,181,31,88,31,75,31,219,31,213,31,96,31,127,31,170,31,110,31,3,31,95,31,27,31,27,30,239,31,223,31,192,31,251,31,119,31,119,30,129,31,250,31,187,31,94,31,94,30,94,29,118,31,118,30,45,31,10,31,10,30,10,29,128,31,64,31,41,31,61,31,106,31,153,31,150,31,223,31,101,31,166,31,243,31,243,30,88,31,111,31,198,31,1,31,158,31,37,31,169,31,191,31,191,30,191,29,190,31,95,31,194,31,38,31,167,31,243,31,71,31,174,31,174,30,2,31,195,31,93,31,141,31,113,31,229,31,219,31,197,31,214,31,214,30,230,31,229,31,144,31,101,31,221,31,248,31,80,31,12,31,144,31,137,31,176,31,177,31,179,31,88,31,98,31,32,31,231,31,248,31,248,30,248,29,248,28,154,31,154,30,150,31,150,30,116,31,18,31,245,31,245,30,232,31,119,31,76,31,183,31,67,31,156,31,230,31,251,31,251,30,16,31,16,30,143,31,220,31,220,31,157,31,150,31,23,31,23,30,93,31,109,31,109,30,5,31,178,31,252,31,40,31,228,31,141,31,107,31,35,31,252,31,141,31,34,31,102,31,163,31,76,31,33,31,33,30,71,31,126,31,126,30,126,29,214,31,214,30,212,31,176,31,10,31,150,31,6,31,47,31,141,31,12,31,52,31,92,31,214,31,85,31,232,31,133,31,163,31,192,31,239,31,201,31,181,31,181,30,80,31,78,31,78,30,61,31,38,31,38,30,10,31,51,31,232,31,32,31,91,31,109,31,205,31,205,30,24,31,163,31,144,31,239,31,215,31,136,31,21,31,11,31,30,31,152,31,96,31,54,31,200,31,46,31,45,31,10,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
