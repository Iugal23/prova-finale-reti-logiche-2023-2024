-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_945 is
end project_tb_945;

architecture project_tb_arch_945 of project_tb_945 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 905;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (113,0,0,0,131,0,185,0,104,0,230,0,157,0,149,0,191,0,205,0,223,0,61,0,22,0,224,0,180,0,44,0,118,0,228,0,71,0,40,0,0,0,27,0,19,0,0,0,15,0,0,0,3,0,226,0,0,0,144,0,183,0,135,0,120,0,187,0,42,0,210,0,206,0,70,0,111,0,27,0,13,0,0,0,197,0,0,0,0,0,112,0,255,0,91,0,225,0,0,0,217,0,34,0,34,0,244,0,0,0,79,0,0,0,0,0,111,0,93,0,227,0,153,0,38,0,224,0,0,0,0,0,220,0,130,0,130,0,58,0,15,0,0,0,61,0,35,0,143,0,0,0,175,0,154,0,0,0,0,0,207,0,250,0,209,0,0,0,72,0,189,0,177,0,252,0,65,0,244,0,48,0,112,0,0,0,175,0,173,0,156,0,249,0,106,0,202,0,137,0,118,0,2,0,30,0,64,0,234,0,114,0,0,0,0,0,254,0,171,0,3,0,47,0,199,0,141,0,98,0,0,0,121,0,217,0,218,0,20,0,0,0,118,0,69,0,241,0,178,0,191,0,0,0,46,0,0,0,0,0,157,0,130,0,6,0,0,0,86,0,115,0,0,0,77,0,98,0,31,0,0,0,128,0,63,0,99,0,72,0,253,0,163,0,147,0,105,0,82,0,255,0,0,0,73,0,140,0,0,0,150,0,62,0,203,0,161,0,122,0,0,0,252,0,61,0,172,0,67,0,0,0,200,0,222,0,0,0,245,0,0,0,78,0,0,0,239,0,0,0,111,0,0,0,198,0,0,0,144,0,136,0,159,0,139,0,162,0,8,0,207,0,17,0,13,0,32,0,139,0,158,0,211,0,160,0,88,0,0,0,0,0,115,0,207,0,53,0,0,0,221,0,229,0,255,0,0,0,69,0,64,0,136,0,16,0,8,0,78,0,3,0,128,0,211,0,221,0,191,0,0,0,89,0,149,0,99,0,158,0,220,0,30,0,118,0,109,0,0,0,247,0,103,0,185,0,56,0,23,0,152,0,105,0,125,0,0,0,171,0,36,0,113,0,201,0,195,0,253,0,84,0,148,0,192,0,0,0,82,0,92,0,189,0,144,0,0,0,0,0,164,0,50,0,190,0,0,0,189,0,0,0,115,0,59,0,163,0,182,0,43,0,154,0,0,0,122,0,0,0,105,0,185,0,168,0,0,0,0,0,187,0,40,0,0,0,189,0,22,0,227,0,58,0,242,0,101,0,80,0,207,0,238,0,29,0,238,0,90,0,0,0,166,0,79,0,55,0,0,0,133,0,68,0,164,0,99,0,0,0,0,0,46,0,31,0,104,0,176,0,5,0,145,0,150,0,52,0,231,0,162,0,38,0,0,0,102,0,7,0,179,0,62,0,25,0,0,0,0,0,0,0,179,0,10,0,96,0,185,0,224,0,91,0,148,0,137,0,189,0,127,0,147,0,0,0,40,0,0,0,0,0,73,0,110,0,0,0,216,0,0,0,196,0,0,0,147,0,100,0,81,0,0,0,180,0,206,0,183,0,0,0,117,0,23,0,40,0,117,0,225,0,146,0,200,0,64,0,208,0,29,0,215,0,39,0,171,0,217,0,0,0,33,0,79,0,0,0,42,0,169,0,66,0,3,0,168,0,145,0,48,0,12,0,198,0,248,0,21,0,82,0,161,0,13,0,121,0,177,0,123,0,112,0,207,0,235,0,0,0,50,0,69,0,137,0,50,0,231,0,0,0,181,0,7,0,20,0,0,0,185,0,53,0,96,0,72,0,199,0,189,0,148,0,134,0,30,0,246,0,182,0,12,0,123,0,0,0,9,0,157,0,12,0,11,0,76,0,203,0,145,0,0,0,0,0,0,0,0,0,217,0,11,0,3,0,25,0,0,0,76,0,152,0,0,0,0,0,108,0,0,0,0,0,132,0,53,0,81,0,187,0,84,0,189,0,185,0,29,0,118,0,0,0,69,0,60,0,32,0,154,0,12,0,59,0,0,0,45,0,139,0,253,0,0,0,0,0,226,0,0,0,25,0,146,0,220,0,30,0,24,0,130,0,54,0,0,0,0,0,110,0,134,0,204,0,177,0,56,0,0,0,246,0,198,0,0,0,7,0,0,0,185,0,76,0,252,0,26,0,0,0,34,0,254,0,0,0,143,0,215,0,254,0,38,0,0,0,19,0,150,0,56,0,231,0,151,0,0,0,0,0,186,0,68,0,41,0,139,0,85,0,0,0,165,0,166,0,85,0,143,0,0,0,141,0,172,0,248,0,4,0,172,0,57,0,218,0,94,0,0,0,28,0,191,0,155,0,47,0,97,0,249,0,215,0,176,0,0,0,125,0,92,0,213,0,159,0,163,0,0,0,255,0,185,0,0,0,5,0,34,0,27,0,0,0,13,0,119,0,225,0,160,0,12,0,212,0,5,0,227,0,105,0,0,0,170,0,179,0,227,0,84,0,210,0,0,0,24,0,0,0,172,0,0,0,237,0,26,0,0,0,196,0,0,0,140,0,107,0,96,0,63,0,222,0,223,0,113,0,0,0,46,0,0,0,132,0,202,0,97,0,171,0,103,0,0,0,218,0,56,0,70,0,89,0,12,0,180,0,0,0,188,0,163,0,0,0,227,0,79,0,222,0,219,0,196,0,233,0,134,0,216,0,0,0,251,0,0,0,4,0,138,0,55,0,82,0,239,0,59,0,173,0,212,0,181,0,233,0,0,0,229,0,151,0,73,0,185,0,169,0,0,0,105,0,98,0,34,0,107,0,0,0,42,0,84,0,56,0,25,0,190,0,46,0,213,0,223,0,0,0,128,0,0,0,0,0,117,0,62,0,19,0,56,0,26,0,0,0,0,0,0,0,237,0,0,0,0,0,138,0,30,0,26,0,91,0,0,0,0,0,19,0,243,0,166,0,0,0,27,0,158,0,42,0,157,0,0,0,0,0,3,0,64,0,157,0,0,0,21,0,10,0,99,0,98,0,32,0,0,0,138,0,32,0,140,0,143,0,208,0,209,0,160,0,214,0,177,0,157,0,206,0,0,0,86,0,156,0,132,0,98,0,47,0,163,0,178,0,165,0,201,0,153,0,197,0,115,0,216,0,0,0,0,0,124,0,0,0,172,0,153,0,84,0,221,0,45,0,87,0,128,0,42,0,86,0,246,0,214,0,224,0,95,0,18,0,139,0,198,0,0,0,127,0,189,0,175,0,34,0,0,0,215,0,138,0,246,0,105,0,65,0,121,0,0,0,101,0,254,0,143,0,192,0,219,0,171,0,12,0,197,0,0,0,174,0,141,0,105,0,0,0,14,0,243,0,81,0,87,0,60,0,4,0,95,0,162,0,0,0,252,0,172,0,8,0,0,0,55,0,0,0,78,0,212,0,39,0,0,0,81,0,216,0,0,0,110,0,238,0,30,0,100,0,21,0,58,0,0,0,75,0,128,0,137,0,0,0,164,0,0,0,133,0,77,0,30,0,230,0,9,0,35,0,0,0,0,0,0,0,64,0,42,0,136,0,100,0,198,0,100,0,169,0,181,0,177,0,160,0,0,0,208,0,180,0,0,0,45,0,0,0,225,0,203,0,213,0,32,0,35,0,187,0,0,0,221,0,74,0,98,0,0,0,0,0,64,0,0,0,200,0,88,0,41,0,32,0,72,0,202,0,100,0,86,0,70,0,142,0,0,0,34,0,0,0,25,0,226,0,62,0,96,0,137,0,0,0,0,0,205,0,61,0,16,0,55,0,0,0,0,0,52,0,124,0,0,0,222,0,141,0,0,0,174,0,154,0,30,0,44,0,113,0,0,0,56,0,0,0,202,0,27,0,209,0,204,0,0,0,123,0,0,0,97,0,66,0,251,0,132,0,147,0,0,0,30,0,0,0,0,0,0,0,0,0,136,0,77,0,204,0,67,0,0,0,0,0,0,0,151,0,89,0,214,0,19,0,134,0,11,0,133,0,126,0,0,0,172,0,8,0,154,0,64,0,104,0,45,0,0,0,184,0,169,0,112,0,22,0,34,0,196,0,215,0,116,0);
signal scenario_full  : scenario_type := (113,31,113,30,131,31,185,31,104,31,230,31,157,31,149,31,191,31,205,31,223,31,61,31,22,31,224,31,180,31,44,31,118,31,228,31,71,31,40,31,40,30,27,31,19,31,19,30,15,31,15,30,3,31,226,31,226,30,144,31,183,31,135,31,120,31,187,31,42,31,210,31,206,31,70,31,111,31,27,31,13,31,13,30,197,31,197,30,197,29,112,31,255,31,91,31,225,31,225,30,217,31,34,31,34,31,244,31,244,30,79,31,79,30,79,29,111,31,93,31,227,31,153,31,38,31,224,31,224,30,224,29,220,31,130,31,130,31,58,31,15,31,15,30,61,31,35,31,143,31,143,30,175,31,154,31,154,30,154,29,207,31,250,31,209,31,209,30,72,31,189,31,177,31,252,31,65,31,244,31,48,31,112,31,112,30,175,31,173,31,156,31,249,31,106,31,202,31,137,31,118,31,2,31,30,31,64,31,234,31,114,31,114,30,114,29,254,31,171,31,3,31,47,31,199,31,141,31,98,31,98,30,121,31,217,31,218,31,20,31,20,30,118,31,69,31,241,31,178,31,191,31,191,30,46,31,46,30,46,29,157,31,130,31,6,31,6,30,86,31,115,31,115,30,77,31,98,31,31,31,31,30,128,31,63,31,99,31,72,31,253,31,163,31,147,31,105,31,82,31,255,31,255,30,73,31,140,31,140,30,150,31,62,31,203,31,161,31,122,31,122,30,252,31,61,31,172,31,67,31,67,30,200,31,222,31,222,30,245,31,245,30,78,31,78,30,239,31,239,30,111,31,111,30,198,31,198,30,144,31,136,31,159,31,139,31,162,31,8,31,207,31,17,31,13,31,32,31,139,31,158,31,211,31,160,31,88,31,88,30,88,29,115,31,207,31,53,31,53,30,221,31,229,31,255,31,255,30,69,31,64,31,136,31,16,31,8,31,78,31,3,31,128,31,211,31,221,31,191,31,191,30,89,31,149,31,99,31,158,31,220,31,30,31,118,31,109,31,109,30,247,31,103,31,185,31,56,31,23,31,152,31,105,31,125,31,125,30,171,31,36,31,113,31,201,31,195,31,253,31,84,31,148,31,192,31,192,30,82,31,92,31,189,31,144,31,144,30,144,29,164,31,50,31,190,31,190,30,189,31,189,30,115,31,59,31,163,31,182,31,43,31,154,31,154,30,122,31,122,30,105,31,185,31,168,31,168,30,168,29,187,31,40,31,40,30,189,31,22,31,227,31,58,31,242,31,101,31,80,31,207,31,238,31,29,31,238,31,90,31,90,30,166,31,79,31,55,31,55,30,133,31,68,31,164,31,99,31,99,30,99,29,46,31,31,31,104,31,176,31,5,31,145,31,150,31,52,31,231,31,162,31,38,31,38,30,102,31,7,31,179,31,62,31,25,31,25,30,25,29,25,28,179,31,10,31,96,31,185,31,224,31,91,31,148,31,137,31,189,31,127,31,147,31,147,30,40,31,40,30,40,29,73,31,110,31,110,30,216,31,216,30,196,31,196,30,147,31,100,31,81,31,81,30,180,31,206,31,183,31,183,30,117,31,23,31,40,31,117,31,225,31,146,31,200,31,64,31,208,31,29,31,215,31,39,31,171,31,217,31,217,30,33,31,79,31,79,30,42,31,169,31,66,31,3,31,168,31,145,31,48,31,12,31,198,31,248,31,21,31,82,31,161,31,13,31,121,31,177,31,123,31,112,31,207,31,235,31,235,30,50,31,69,31,137,31,50,31,231,31,231,30,181,31,7,31,20,31,20,30,185,31,53,31,96,31,72,31,199,31,189,31,148,31,134,31,30,31,246,31,182,31,12,31,123,31,123,30,9,31,157,31,12,31,11,31,76,31,203,31,145,31,145,30,145,29,145,28,145,27,217,31,11,31,3,31,25,31,25,30,76,31,152,31,152,30,152,29,108,31,108,30,108,29,132,31,53,31,81,31,187,31,84,31,189,31,185,31,29,31,118,31,118,30,69,31,60,31,32,31,154,31,12,31,59,31,59,30,45,31,139,31,253,31,253,30,253,29,226,31,226,30,25,31,146,31,220,31,30,31,24,31,130,31,54,31,54,30,54,29,110,31,134,31,204,31,177,31,56,31,56,30,246,31,198,31,198,30,7,31,7,30,185,31,76,31,252,31,26,31,26,30,34,31,254,31,254,30,143,31,215,31,254,31,38,31,38,30,19,31,150,31,56,31,231,31,151,31,151,30,151,29,186,31,68,31,41,31,139,31,85,31,85,30,165,31,166,31,85,31,143,31,143,30,141,31,172,31,248,31,4,31,172,31,57,31,218,31,94,31,94,30,28,31,191,31,155,31,47,31,97,31,249,31,215,31,176,31,176,30,125,31,92,31,213,31,159,31,163,31,163,30,255,31,185,31,185,30,5,31,34,31,27,31,27,30,13,31,119,31,225,31,160,31,12,31,212,31,5,31,227,31,105,31,105,30,170,31,179,31,227,31,84,31,210,31,210,30,24,31,24,30,172,31,172,30,237,31,26,31,26,30,196,31,196,30,140,31,107,31,96,31,63,31,222,31,223,31,113,31,113,30,46,31,46,30,132,31,202,31,97,31,171,31,103,31,103,30,218,31,56,31,70,31,89,31,12,31,180,31,180,30,188,31,163,31,163,30,227,31,79,31,222,31,219,31,196,31,233,31,134,31,216,31,216,30,251,31,251,30,4,31,138,31,55,31,82,31,239,31,59,31,173,31,212,31,181,31,233,31,233,30,229,31,151,31,73,31,185,31,169,31,169,30,105,31,98,31,34,31,107,31,107,30,42,31,84,31,56,31,25,31,190,31,46,31,213,31,223,31,223,30,128,31,128,30,128,29,117,31,62,31,19,31,56,31,26,31,26,30,26,29,26,28,237,31,237,30,237,29,138,31,30,31,26,31,91,31,91,30,91,29,19,31,243,31,166,31,166,30,27,31,158,31,42,31,157,31,157,30,157,29,3,31,64,31,157,31,157,30,21,31,10,31,99,31,98,31,32,31,32,30,138,31,32,31,140,31,143,31,208,31,209,31,160,31,214,31,177,31,157,31,206,31,206,30,86,31,156,31,132,31,98,31,47,31,163,31,178,31,165,31,201,31,153,31,197,31,115,31,216,31,216,30,216,29,124,31,124,30,172,31,153,31,84,31,221,31,45,31,87,31,128,31,42,31,86,31,246,31,214,31,224,31,95,31,18,31,139,31,198,31,198,30,127,31,189,31,175,31,34,31,34,30,215,31,138,31,246,31,105,31,65,31,121,31,121,30,101,31,254,31,143,31,192,31,219,31,171,31,12,31,197,31,197,30,174,31,141,31,105,31,105,30,14,31,243,31,81,31,87,31,60,31,4,31,95,31,162,31,162,30,252,31,172,31,8,31,8,30,55,31,55,30,78,31,212,31,39,31,39,30,81,31,216,31,216,30,110,31,238,31,30,31,100,31,21,31,58,31,58,30,75,31,128,31,137,31,137,30,164,31,164,30,133,31,77,31,30,31,230,31,9,31,35,31,35,30,35,29,35,28,64,31,42,31,136,31,100,31,198,31,100,31,169,31,181,31,177,31,160,31,160,30,208,31,180,31,180,30,45,31,45,30,225,31,203,31,213,31,32,31,35,31,187,31,187,30,221,31,74,31,98,31,98,30,98,29,64,31,64,30,200,31,88,31,41,31,32,31,72,31,202,31,100,31,86,31,70,31,142,31,142,30,34,31,34,30,25,31,226,31,62,31,96,31,137,31,137,30,137,29,205,31,61,31,16,31,55,31,55,30,55,29,52,31,124,31,124,30,222,31,141,31,141,30,174,31,154,31,30,31,44,31,113,31,113,30,56,31,56,30,202,31,27,31,209,31,204,31,204,30,123,31,123,30,97,31,66,31,251,31,132,31,147,31,147,30,30,31,30,30,30,29,30,28,30,27,136,31,77,31,204,31,67,31,67,30,67,29,67,28,151,31,89,31,214,31,19,31,134,31,11,31,133,31,126,31,126,30,172,31,8,31,154,31,64,31,104,31,45,31,45,30,184,31,169,31,112,31,22,31,34,31,196,31,215,31,116,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
