-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_219 is
end project_tb_219;

architecture project_tb_arch_219 of project_tb_219 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 924;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (90,0,172,0,168,0,57,0,198,0,151,0,29,0,197,0,43,0,81,0,3,0,7,0,59,0,95,0,108,0,107,0,172,0,141,0,0,0,138,0,112,0,34,0,0,0,146,0,43,0,0,0,178,0,0,0,19,0,0,0,246,0,20,0,0,0,158,0,0,0,4,0,225,0,24,0,103,0,254,0,0,0,115,0,6,0,191,0,125,0,45,0,0,0,139,0,249,0,222,0,45,0,73,0,162,0,146,0,75,0,229,0,44,0,0,0,239,0,0,0,135,0,0,0,0,0,155,0,44,0,196,0,231,0,133,0,156,0,17,0,34,0,0,0,240,0,0,0,5,0,61,0,36,0,197,0,30,0,143,0,164,0,249,0,19,0,55,0,26,0,0,0,248,0,146,0,113,0,97,0,221,0,227,0,87,0,0,0,0,0,166,0,143,0,216,0,161,0,149,0,128,0,0,0,0,0,65,0,0,0,0,0,111,0,133,0,214,0,130,0,108,0,32,0,13,0,202,0,0,0,243,0,11,0,192,0,197,0,221,0,127,0,71,0,20,0,169,0,0,0,65,0,78,0,117,0,41,0,0,0,108,0,115,0,0,0,222,0,250,0,146,0,59,0,84,0,78,0,109,0,44,0,137,0,146,0,0,0,0,0,0,0,39,0,203,0,0,0,111,0,100,0,121,0,133,0,212,0,100,0,51,0,161,0,192,0,34,0,249,0,57,0,53,0,112,0,98,0,0,0,228,0,22,0,68,0,255,0,194,0,190,0,23,0,30,0,174,0,27,0,75,0,72,0,183,0,74,0,111,0,0,0,215,0,185,0,214,0,114,0,119,0,0,0,0,0,123,0,176,0,104,0,68,0,91,0,78,0,96,0,175,0,64,0,0,0,232,0,167,0,63,0,0,0,27,0,126,0,123,0,188,0,86,0,211,0,132,0,132,0,31,0,84,0,14,0,65,0,88,0,165,0,71,0,93,0,234,0,132,0,82,0,0,0,115,0,211,0,0,0,90,0,0,0,84,0,173,0,185,0,119,0,202,0,125,0,40,0,249,0,0,0,173,0,135,0,192,0,0,0,240,0,122,0,92,0,217,0,115,0,113,0,0,0,188,0,147,0,0,0,126,0,89,0,81,0,0,0,128,0,0,0,72,0,133,0,0,0,131,0,203,0,0,0,216,0,183,0,198,0,0,0,0,0,20,0,78,0,210,0,0,0,89,0,32,0,0,0,204,0,113,0,23,0,95,0,143,0,0,0,115,0,0,0,154,0,168,0,15,0,66,0,35,0,0,0,72,0,88,0,156,0,247,0,74,0,182,0,225,0,155,0,173,0,0,0,0,0,123,0,137,0,89,0,192,0,126,0,91,0,235,0,152,0,36,0,165,0,10,0,245,0,126,0,0,0,0,0,0,0,30,0,136,0,1,0,158,0,0,0,110,0,52,0,132,0,56,0,108,0,41,0,27,0,131,0,192,0,229,0,58,0,31,0,0,0,146,0,17,0,170,0,21,0,211,0,68,0,76,0,43,0,0,0,195,0,193,0,193,0,88,0,12,0,213,0,49,0,0,0,52,0,34,0,0,0,7,0,75,0,229,0,131,0,113,0,91,0,63,0,165,0,182,0,228,0,111,0,73,0,164,0,205,0,14,0,0,0,36,0,185,0,54,0,104,0,45,0,198,0,222,0,38,0,35,0,123,0,214,0,134,0,185,0,74,0,174,0,30,0,191,0,178,0,127,0,178,0,0,0,71,0,28,0,0,0,174,0,3,0,123,0,0,0,65,0,68,0,0,0,53,0,0,0,110,0,179,0,0,0,0,0,134,0,110,0,240,0,232,0,189,0,207,0,80,0,244,0,21,0,107,0,30,0,215,0,218,0,145,0,1,0,0,0,0,0,51,0,0,0,0,0,35,0,49,0,170,0,202,0,0,0,0,0,178,0,0,0,215,0,58,0,222,0,185,0,64,0,0,0,0,0,0,0,0,0,186,0,38,0,251,0,222,0,0,0,202,0,85,0,5,0,18,0,212,0,98,0,0,0,238,0,93,0,239,0,137,0,0,0,223,0,254,0,192,0,0,0,116,0,96,0,101,0,144,0,130,0,217,0,206,0,53,0,103,0,166,0,112,0,233,0,31,0,75,0,234,0,0,0,73,0,210,0,0,0,13,0,65,0,234,0,111,0,211,0,67,0,130,0,43,0,9,0,0,0,0,0,2,0,187,0,249,0,22,0,0,0,215,0,201,0,0,0,132,0,28,0,0,0,0,0,38,0,0,0,214,0,65,0,0,0,166,0,0,0,205,0,67,0,66,0,19,0,195,0,134,0,229,0,114,0,199,0,0,0,167,0,147,0,0,0,15,0,0,0,0,0,84,0,45,0,113,0,32,0,110,0,105,0,188,0,254,0,236,0,175,0,117,0,214,0,3,0,0,0,162,0,141,0,205,0,0,0,0,0,184,0,186,0,167,0,236,0,151,0,0,0,63,0,222,0,95,0,0,0,206,0,124,0,247,0,28,0,182,0,145,0,65,0,192,0,180,0,46,0,109,0,57,0,13,0,176,0,50,0,139,0,0,0,21,0,240,0,182,0,0,0,191,0,209,0,115,0,0,0,35,0,39,0,0,0,0,0,70,0,191,0,0,0,58,0,0,0,117,0,139,0,26,0,0,0,180,0,150,0,122,0,0,0,1,0,105,0,0,0,113,0,51,0,0,0,170,0,183,0,0,0,46,0,232,0,226,0,176,0,143,0,52,0,146,0,231,0,61,0,165,0,0,0,74,0,0,0,86,0,151,0,190,0,88,0,31,0,54,0,199,0,0,0,0,0,114,0,53,0,95,0,78,0,9,0,245,0,27,0,0,0,73,0,79,0,162,0,211,0,105,0,0,0,245,0,46,0,2,0,5,0,54,0,27,0,191,0,34,0,207,0,0,0,224,0,86,0,224,0,0,0,4,0,12,0,0,0,94,0,169,0,122,0,72,0,7,0,12,0,192,0,0,0,13,0,238,0,108,0,127,0,0,0,64,0,184,0,0,0,175,0,68,0,0,0,62,0,197,0,105,0,138,0,0,0,168,0,80,0,126,0,240,0,115,0,133,0,8,0,234,0,73,0,127,0,11,0,192,0,210,0,251,0,122,0,106,0,0,0,24,0,218,0,83,0,46,0,44,0,137,0,210,0,185,0,175,0,148,0,191,0,0,0,198,0,75,0,158,0,89,0,70,0,173,0,110,0,228,0,0,0,84,0,148,0,181,0,94,0,128,0,48,0,90,0,19,0,1,0,249,0,223,0,18,0,33,0,244,0,246,0,0,0,72,0,135,0,0,0,0,0,57,0,0,0,0,0,18,0,103,0,0,0,0,0,0,0,0,0,215,0,213,0,0,0,113,0,247,0,136,0,48,0,0,0,100,0,2,0,0,0,52,0,135,0,110,0,54,0,110,0,0,0,254,0,51,0,214,0,245,0,0,0,121,0,164,0,137,0,215,0,112,0,87,0,53,0,49,0,73,0,243,0,73,0,18,0,0,0,187,0,35,0,136,0,243,0,0,0,10,0,221,0,68,0,216,0,13,0,178,0,0,0,0,0,45,0,0,0,181,0,0,0,62,0,7,0,193,0,0,0,122,0,49,0,91,0,50,0,133,0,0,0,211,0,10,0,8,0,233,0,0,0,183,0,99,0,236,0,230,0,144,0,72,0,233,0,0,0,0,0,0,0,216,0,100,0,26,0,193,0,43,0,227,0,150,0,37,0,193,0,61,0,118,0,0,0,0,0,99,0,237,0,241,0,118,0,0,0,168,0,4,0,34,0,218,0,0,0,68,0,242,0,229,0,157,0,0,0,41,0,47,0,59,0,1,0,163,0,219,0,189,0,229,0,96,0,24,0,0,0,164,0,119,0,182,0,3,0,100,0,0,0,46,0,26,0,152,0,63,0,140,0,154,0,4,0,108,0,0,0,236,0,186,0,155,0,21,0,71,0,234,0,122,0,228,0,140,0,248,0,0,0,100,0,37,0,4,0,0,0,74,0,147,0,217,0,169,0,56,0,130,0,0,0,22,0,72,0,176,0,191,0,59,0,40,0,80,0,109,0,0,0,124,0,17,0,136,0,0,0,154,0,110,0,197,0,72,0,128,0);
signal scenario_full  : scenario_type := (90,31,172,31,168,31,57,31,198,31,151,31,29,31,197,31,43,31,81,31,3,31,7,31,59,31,95,31,108,31,107,31,172,31,141,31,141,30,138,31,112,31,34,31,34,30,146,31,43,31,43,30,178,31,178,30,19,31,19,30,246,31,20,31,20,30,158,31,158,30,4,31,225,31,24,31,103,31,254,31,254,30,115,31,6,31,191,31,125,31,45,31,45,30,139,31,249,31,222,31,45,31,73,31,162,31,146,31,75,31,229,31,44,31,44,30,239,31,239,30,135,31,135,30,135,29,155,31,44,31,196,31,231,31,133,31,156,31,17,31,34,31,34,30,240,31,240,30,5,31,61,31,36,31,197,31,30,31,143,31,164,31,249,31,19,31,55,31,26,31,26,30,248,31,146,31,113,31,97,31,221,31,227,31,87,31,87,30,87,29,166,31,143,31,216,31,161,31,149,31,128,31,128,30,128,29,65,31,65,30,65,29,111,31,133,31,214,31,130,31,108,31,32,31,13,31,202,31,202,30,243,31,11,31,192,31,197,31,221,31,127,31,71,31,20,31,169,31,169,30,65,31,78,31,117,31,41,31,41,30,108,31,115,31,115,30,222,31,250,31,146,31,59,31,84,31,78,31,109,31,44,31,137,31,146,31,146,30,146,29,146,28,39,31,203,31,203,30,111,31,100,31,121,31,133,31,212,31,100,31,51,31,161,31,192,31,34,31,249,31,57,31,53,31,112,31,98,31,98,30,228,31,22,31,68,31,255,31,194,31,190,31,23,31,30,31,174,31,27,31,75,31,72,31,183,31,74,31,111,31,111,30,215,31,185,31,214,31,114,31,119,31,119,30,119,29,123,31,176,31,104,31,68,31,91,31,78,31,96,31,175,31,64,31,64,30,232,31,167,31,63,31,63,30,27,31,126,31,123,31,188,31,86,31,211,31,132,31,132,31,31,31,84,31,14,31,65,31,88,31,165,31,71,31,93,31,234,31,132,31,82,31,82,30,115,31,211,31,211,30,90,31,90,30,84,31,173,31,185,31,119,31,202,31,125,31,40,31,249,31,249,30,173,31,135,31,192,31,192,30,240,31,122,31,92,31,217,31,115,31,113,31,113,30,188,31,147,31,147,30,126,31,89,31,81,31,81,30,128,31,128,30,72,31,133,31,133,30,131,31,203,31,203,30,216,31,183,31,198,31,198,30,198,29,20,31,78,31,210,31,210,30,89,31,32,31,32,30,204,31,113,31,23,31,95,31,143,31,143,30,115,31,115,30,154,31,168,31,15,31,66,31,35,31,35,30,72,31,88,31,156,31,247,31,74,31,182,31,225,31,155,31,173,31,173,30,173,29,123,31,137,31,89,31,192,31,126,31,91,31,235,31,152,31,36,31,165,31,10,31,245,31,126,31,126,30,126,29,126,28,30,31,136,31,1,31,158,31,158,30,110,31,52,31,132,31,56,31,108,31,41,31,27,31,131,31,192,31,229,31,58,31,31,31,31,30,146,31,17,31,170,31,21,31,211,31,68,31,76,31,43,31,43,30,195,31,193,31,193,31,88,31,12,31,213,31,49,31,49,30,52,31,34,31,34,30,7,31,75,31,229,31,131,31,113,31,91,31,63,31,165,31,182,31,228,31,111,31,73,31,164,31,205,31,14,31,14,30,36,31,185,31,54,31,104,31,45,31,198,31,222,31,38,31,35,31,123,31,214,31,134,31,185,31,74,31,174,31,30,31,191,31,178,31,127,31,178,31,178,30,71,31,28,31,28,30,174,31,3,31,123,31,123,30,65,31,68,31,68,30,53,31,53,30,110,31,179,31,179,30,179,29,134,31,110,31,240,31,232,31,189,31,207,31,80,31,244,31,21,31,107,31,30,31,215,31,218,31,145,31,1,31,1,30,1,29,51,31,51,30,51,29,35,31,49,31,170,31,202,31,202,30,202,29,178,31,178,30,215,31,58,31,222,31,185,31,64,31,64,30,64,29,64,28,64,27,186,31,38,31,251,31,222,31,222,30,202,31,85,31,5,31,18,31,212,31,98,31,98,30,238,31,93,31,239,31,137,31,137,30,223,31,254,31,192,31,192,30,116,31,96,31,101,31,144,31,130,31,217,31,206,31,53,31,103,31,166,31,112,31,233,31,31,31,75,31,234,31,234,30,73,31,210,31,210,30,13,31,65,31,234,31,111,31,211,31,67,31,130,31,43,31,9,31,9,30,9,29,2,31,187,31,249,31,22,31,22,30,215,31,201,31,201,30,132,31,28,31,28,30,28,29,38,31,38,30,214,31,65,31,65,30,166,31,166,30,205,31,67,31,66,31,19,31,195,31,134,31,229,31,114,31,199,31,199,30,167,31,147,31,147,30,15,31,15,30,15,29,84,31,45,31,113,31,32,31,110,31,105,31,188,31,254,31,236,31,175,31,117,31,214,31,3,31,3,30,162,31,141,31,205,31,205,30,205,29,184,31,186,31,167,31,236,31,151,31,151,30,63,31,222,31,95,31,95,30,206,31,124,31,247,31,28,31,182,31,145,31,65,31,192,31,180,31,46,31,109,31,57,31,13,31,176,31,50,31,139,31,139,30,21,31,240,31,182,31,182,30,191,31,209,31,115,31,115,30,35,31,39,31,39,30,39,29,70,31,191,31,191,30,58,31,58,30,117,31,139,31,26,31,26,30,180,31,150,31,122,31,122,30,1,31,105,31,105,30,113,31,51,31,51,30,170,31,183,31,183,30,46,31,232,31,226,31,176,31,143,31,52,31,146,31,231,31,61,31,165,31,165,30,74,31,74,30,86,31,151,31,190,31,88,31,31,31,54,31,199,31,199,30,199,29,114,31,53,31,95,31,78,31,9,31,245,31,27,31,27,30,73,31,79,31,162,31,211,31,105,31,105,30,245,31,46,31,2,31,5,31,54,31,27,31,191,31,34,31,207,31,207,30,224,31,86,31,224,31,224,30,4,31,12,31,12,30,94,31,169,31,122,31,72,31,7,31,12,31,192,31,192,30,13,31,238,31,108,31,127,31,127,30,64,31,184,31,184,30,175,31,68,31,68,30,62,31,197,31,105,31,138,31,138,30,168,31,80,31,126,31,240,31,115,31,133,31,8,31,234,31,73,31,127,31,11,31,192,31,210,31,251,31,122,31,106,31,106,30,24,31,218,31,83,31,46,31,44,31,137,31,210,31,185,31,175,31,148,31,191,31,191,30,198,31,75,31,158,31,89,31,70,31,173,31,110,31,228,31,228,30,84,31,148,31,181,31,94,31,128,31,48,31,90,31,19,31,1,31,249,31,223,31,18,31,33,31,244,31,246,31,246,30,72,31,135,31,135,30,135,29,57,31,57,30,57,29,18,31,103,31,103,30,103,29,103,28,103,27,215,31,213,31,213,30,113,31,247,31,136,31,48,31,48,30,100,31,2,31,2,30,52,31,135,31,110,31,54,31,110,31,110,30,254,31,51,31,214,31,245,31,245,30,121,31,164,31,137,31,215,31,112,31,87,31,53,31,49,31,73,31,243,31,73,31,18,31,18,30,187,31,35,31,136,31,243,31,243,30,10,31,221,31,68,31,216,31,13,31,178,31,178,30,178,29,45,31,45,30,181,31,181,30,62,31,7,31,193,31,193,30,122,31,49,31,91,31,50,31,133,31,133,30,211,31,10,31,8,31,233,31,233,30,183,31,99,31,236,31,230,31,144,31,72,31,233,31,233,30,233,29,233,28,216,31,100,31,26,31,193,31,43,31,227,31,150,31,37,31,193,31,61,31,118,31,118,30,118,29,99,31,237,31,241,31,118,31,118,30,168,31,4,31,34,31,218,31,218,30,68,31,242,31,229,31,157,31,157,30,41,31,47,31,59,31,1,31,163,31,219,31,189,31,229,31,96,31,24,31,24,30,164,31,119,31,182,31,3,31,100,31,100,30,46,31,26,31,152,31,63,31,140,31,154,31,4,31,108,31,108,30,236,31,186,31,155,31,21,31,71,31,234,31,122,31,228,31,140,31,248,31,248,30,100,31,37,31,4,31,4,30,74,31,147,31,217,31,169,31,56,31,130,31,130,30,22,31,72,31,176,31,191,31,59,31,40,31,80,31,109,31,109,30,124,31,17,31,136,31,136,30,154,31,110,31,197,31,72,31,128,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
