-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_94 is
end project_tb_94;

architecture project_tb_arch_94 of project_tb_94 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 745;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (39,0,0,0,126,0,0,0,193,0,100,0,182,0,183,0,234,0,77,0,60,0,70,0,0,0,243,0,229,0,61,0,119,0,25,0,214,0,0,0,231,0,239,0,147,0,93,0,241,0,94,0,0,0,188,0,6,0,100,0,0,0,212,0,251,0,0,0,174,0,212,0,205,0,196,0,81,0,130,0,84,0,12,0,0,0,111,0,15,0,0,0,135,0,17,0,91,0,69,0,68,0,161,0,189,0,106,0,0,0,181,0,73,0,40,0,5,0,0,0,0,0,205,0,227,0,0,0,163,0,0,0,235,0,0,0,104,0,145,0,137,0,60,0,139,0,107,0,41,0,184,0,223,0,0,0,77,0,158,0,0,0,231,0,44,0,24,0,0,0,71,0,237,0,138,0,36,0,46,0,141,0,82,0,159,0,72,0,240,0,152,0,76,0,21,0,73,0,89,0,0,0,116,0,0,0,103,0,0,0,20,0,224,0,137,0,0,0,151,0,152,0,0,0,25,0,56,0,52,0,93,0,239,0,11,0,240,0,0,0,0,0,183,0,191,0,165,0,252,0,18,0,0,0,164,0,129,0,0,0,216,0,0,0,0,0,8,0,240,0,0,0,40,0,56,0,197,0,138,0,208,0,71,0,95,0,214,0,16,0,129,0,150,0,197,0,132,0,174,0,179,0,204,0,194,0,167,0,147,0,75,0,152,0,86,0,104,0,196,0,180,0,0,0,52,0,193,0,114,0,0,0,194,0,117,0,212,0,238,0,29,0,151,0,48,0,210,0,127,0,45,0,17,0,176,0,0,0,78,0,83,0,0,0,42,0,203,0,158,0,177,0,235,0,170,0,204,0,126,0,231,0,4,0,87,0,36,0,77,0,16,0,27,0,183,0,5,0,38,0,189,0,0,0,53,0,176,0,13,0,64,0,64,0,181,0,0,0,68,0,107,0,81,0,184,0,222,0,154,0,65,0,185,0,29,0,8,0,101,0,76,0,91,0,90,0,250,0,114,0,146,0,230,0,25,0,0,0,0,0,64,0,0,0,140,0,188,0,134,0,163,0,215,0,195,0,0,0,96,0,93,0,52,0,53,0,254,0,6,0,99,0,67,0,85,0,0,0,238,0,146,0,87,0,0,0,211,0,229,0,0,0,145,0,233,0,135,0,169,0,252,0,172,0,73,0,0,0,173,0,0,0,125,0,215,0,0,0,220,0,178,0,131,0,95,0,3,0,32,0,41,0,32,0,0,0,197,0,0,0,81,0,151,0,30,0,24,0,254,0,24,0,227,0,115,0,79,0,0,0,113,0,126,0,16,0,194,0,6,0,139,0,87,0,117,0,210,0,225,0,247,0,143,0,0,0,33,0,0,0,104,0,32,0,46,0,227,0,28,0,248,0,62,0,0,0,174,0,83,0,245,0,43,0,175,0,250,0,0,0,0,0,223,0,154,0,28,0,220,0,0,0,40,0,59,0,15,0,245,0,212,0,0,0,164,0,241,0,129,0,0,0,168,0,114,0,119,0,142,0,231,0,228,0,198,0,105,0,80,0,49,0,1,0,219,0,63,0,219,0,137,0,227,0,62,0,230,0,135,0,0,0,106,0,78,0,76,0,0,0,0,0,120,0,63,0,56,0,94,0,0,0,208,0,0,0,120,0,60,0,71,0,199,0,0,0,156,0,58,0,122,0,124,0,206,0,8,0,151,0,180,0,0,0,0,0,39,0,61,0,25,0,0,0,0,0,19,0,0,0,132,0,85,0,238,0,253,0,165,0,54,0,154,0,0,0,101,0,126,0,159,0,195,0,97,0,206,0,235,0,161,0,214,0,113,0,217,0,83,0,167,0,237,0,246,0,11,0,135,0,0,0,199,0,0,0,50,0,3,0,222,0,100,0,105,0,79,0,0,0,30,0,209,0,227,0,0,0,218,0,144,0,151,0,95,0,173,0,27,0,245,0,172,0,28,0,114,0,124,0,0,0,100,0,0,0,174,0,66,0,178,0,139,0,83,0,255,0,51,0,0,0,73,0,206,0,180,0,0,0,240,0,224,0,81,0,0,0,94,0,191,0,120,0,13,0,60,0,76,0,0,0,119,0,0,0,81,0,116,0,32,0,0,0,113,0,0,0,76,0,116,0,167,0,25,0,245,0,0,0,190,0,229,0,172,0,63,0,8,0,235,0,0,0,192,0,235,0,204,0,244,0,237,0,199,0,97,0,0,0,86,0,136,0,119,0,177,0,155,0,209,0,89,0,0,0,226,0,108,0,179,0,94,0,77,0,12,0,85,0,231,0,0,0,0,0,30,0,73,0,103,0,63,0,211,0,54,0,10,0,219,0,243,0,0,0,0,0,96,0,243,0,165,0,0,0,113,0,47,0,118,0,6,0,0,0,0,0,219,0,0,0,231,0,0,0,171,0,76,0,51,0,0,0,88,0,188,0,95,0,15,0,208,0,187,0,188,0,46,0,45,0,53,0,0,0,143,0,63,0,132,0,236,0,103,0,0,0,78,0,181,0,60,0,0,0,137,0,79,0,191,0,55,0,0,0,75,0,105,0,152,0,0,0,242,0,109,0,238,0,34,0,200,0,0,0,98,0,0,0,239,0,40,0,247,0,148,0,0,0,15,0,213,0,0,0,0,0,191,0,108,0,0,0,157,0,223,0,12,0,248,0,10,0,22,0,28,0,50,0,0,0,112,0,0,0,42,0,28,0,0,0,214,0,215,0,86,0,116,0,0,0,153,0,0,0,0,0,12,0,216,0,7,0,50,0,0,0,64,0,0,0,239,0,0,0,194,0,214,0,187,0,112,0,0,0,182,0,179,0,249,0,106,0,201,0,73,0,246,0,255,0,206,0,107,0,164,0,145,0,24,0,0,0,165,0,123,0,135,0,0,0,225,0,145,0,136,0,193,0,243,0,75,0,0,0,155,0,70,0,184,0,231,0,0,0,96,0,216,0,0,0,0,0,25,0,212,0,171,0,210,0,219,0,226,0,0,0,36,0,0,0,161,0,179,0,220,0,0,0,0,0,53,0,181,0,147,0,249,0,132,0,0,0,162,0,191,0,173,0,9,0,107,0,245,0,54,0,253,0,193,0,0,0,0,0,0,0,41,0,225,0,69,0,169,0,0,0,81,0,109,0,100,0,166,0,61,0,0,0,179,0,0,0,254,0,221,0,45,0,119,0,165,0,67,0,78,0,176,0,235,0,19,0,86,0,95,0,170,0,0,0,118,0,0,0,89,0,47,0,0,0,127,0,0,0,3,0,0,0,129,0,79,0,202,0,205,0,28,0,51,0,79,0,198,0,190,0,0,0,81,0,65,0,101,0,88,0,0,0);
signal scenario_full  : scenario_type := (39,31,39,30,126,31,126,30,193,31,100,31,182,31,183,31,234,31,77,31,60,31,70,31,70,30,243,31,229,31,61,31,119,31,25,31,214,31,214,30,231,31,239,31,147,31,93,31,241,31,94,31,94,30,188,31,6,31,100,31,100,30,212,31,251,31,251,30,174,31,212,31,205,31,196,31,81,31,130,31,84,31,12,31,12,30,111,31,15,31,15,30,135,31,17,31,91,31,69,31,68,31,161,31,189,31,106,31,106,30,181,31,73,31,40,31,5,31,5,30,5,29,205,31,227,31,227,30,163,31,163,30,235,31,235,30,104,31,145,31,137,31,60,31,139,31,107,31,41,31,184,31,223,31,223,30,77,31,158,31,158,30,231,31,44,31,24,31,24,30,71,31,237,31,138,31,36,31,46,31,141,31,82,31,159,31,72,31,240,31,152,31,76,31,21,31,73,31,89,31,89,30,116,31,116,30,103,31,103,30,20,31,224,31,137,31,137,30,151,31,152,31,152,30,25,31,56,31,52,31,93,31,239,31,11,31,240,31,240,30,240,29,183,31,191,31,165,31,252,31,18,31,18,30,164,31,129,31,129,30,216,31,216,30,216,29,8,31,240,31,240,30,40,31,56,31,197,31,138,31,208,31,71,31,95,31,214,31,16,31,129,31,150,31,197,31,132,31,174,31,179,31,204,31,194,31,167,31,147,31,75,31,152,31,86,31,104,31,196,31,180,31,180,30,52,31,193,31,114,31,114,30,194,31,117,31,212,31,238,31,29,31,151,31,48,31,210,31,127,31,45,31,17,31,176,31,176,30,78,31,83,31,83,30,42,31,203,31,158,31,177,31,235,31,170,31,204,31,126,31,231,31,4,31,87,31,36,31,77,31,16,31,27,31,183,31,5,31,38,31,189,31,189,30,53,31,176,31,13,31,64,31,64,31,181,31,181,30,68,31,107,31,81,31,184,31,222,31,154,31,65,31,185,31,29,31,8,31,101,31,76,31,91,31,90,31,250,31,114,31,146,31,230,31,25,31,25,30,25,29,64,31,64,30,140,31,188,31,134,31,163,31,215,31,195,31,195,30,96,31,93,31,52,31,53,31,254,31,6,31,99,31,67,31,85,31,85,30,238,31,146,31,87,31,87,30,211,31,229,31,229,30,145,31,233,31,135,31,169,31,252,31,172,31,73,31,73,30,173,31,173,30,125,31,215,31,215,30,220,31,178,31,131,31,95,31,3,31,32,31,41,31,32,31,32,30,197,31,197,30,81,31,151,31,30,31,24,31,254,31,24,31,227,31,115,31,79,31,79,30,113,31,126,31,16,31,194,31,6,31,139,31,87,31,117,31,210,31,225,31,247,31,143,31,143,30,33,31,33,30,104,31,32,31,46,31,227,31,28,31,248,31,62,31,62,30,174,31,83,31,245,31,43,31,175,31,250,31,250,30,250,29,223,31,154,31,28,31,220,31,220,30,40,31,59,31,15,31,245,31,212,31,212,30,164,31,241,31,129,31,129,30,168,31,114,31,119,31,142,31,231,31,228,31,198,31,105,31,80,31,49,31,1,31,219,31,63,31,219,31,137,31,227,31,62,31,230,31,135,31,135,30,106,31,78,31,76,31,76,30,76,29,120,31,63,31,56,31,94,31,94,30,208,31,208,30,120,31,60,31,71,31,199,31,199,30,156,31,58,31,122,31,124,31,206,31,8,31,151,31,180,31,180,30,180,29,39,31,61,31,25,31,25,30,25,29,19,31,19,30,132,31,85,31,238,31,253,31,165,31,54,31,154,31,154,30,101,31,126,31,159,31,195,31,97,31,206,31,235,31,161,31,214,31,113,31,217,31,83,31,167,31,237,31,246,31,11,31,135,31,135,30,199,31,199,30,50,31,3,31,222,31,100,31,105,31,79,31,79,30,30,31,209,31,227,31,227,30,218,31,144,31,151,31,95,31,173,31,27,31,245,31,172,31,28,31,114,31,124,31,124,30,100,31,100,30,174,31,66,31,178,31,139,31,83,31,255,31,51,31,51,30,73,31,206,31,180,31,180,30,240,31,224,31,81,31,81,30,94,31,191,31,120,31,13,31,60,31,76,31,76,30,119,31,119,30,81,31,116,31,32,31,32,30,113,31,113,30,76,31,116,31,167,31,25,31,245,31,245,30,190,31,229,31,172,31,63,31,8,31,235,31,235,30,192,31,235,31,204,31,244,31,237,31,199,31,97,31,97,30,86,31,136,31,119,31,177,31,155,31,209,31,89,31,89,30,226,31,108,31,179,31,94,31,77,31,12,31,85,31,231,31,231,30,231,29,30,31,73,31,103,31,63,31,211,31,54,31,10,31,219,31,243,31,243,30,243,29,96,31,243,31,165,31,165,30,113,31,47,31,118,31,6,31,6,30,6,29,219,31,219,30,231,31,231,30,171,31,76,31,51,31,51,30,88,31,188,31,95,31,15,31,208,31,187,31,188,31,46,31,45,31,53,31,53,30,143,31,63,31,132,31,236,31,103,31,103,30,78,31,181,31,60,31,60,30,137,31,79,31,191,31,55,31,55,30,75,31,105,31,152,31,152,30,242,31,109,31,238,31,34,31,200,31,200,30,98,31,98,30,239,31,40,31,247,31,148,31,148,30,15,31,213,31,213,30,213,29,191,31,108,31,108,30,157,31,223,31,12,31,248,31,10,31,22,31,28,31,50,31,50,30,112,31,112,30,42,31,28,31,28,30,214,31,215,31,86,31,116,31,116,30,153,31,153,30,153,29,12,31,216,31,7,31,50,31,50,30,64,31,64,30,239,31,239,30,194,31,214,31,187,31,112,31,112,30,182,31,179,31,249,31,106,31,201,31,73,31,246,31,255,31,206,31,107,31,164,31,145,31,24,31,24,30,165,31,123,31,135,31,135,30,225,31,145,31,136,31,193,31,243,31,75,31,75,30,155,31,70,31,184,31,231,31,231,30,96,31,216,31,216,30,216,29,25,31,212,31,171,31,210,31,219,31,226,31,226,30,36,31,36,30,161,31,179,31,220,31,220,30,220,29,53,31,181,31,147,31,249,31,132,31,132,30,162,31,191,31,173,31,9,31,107,31,245,31,54,31,253,31,193,31,193,30,193,29,193,28,41,31,225,31,69,31,169,31,169,30,81,31,109,31,100,31,166,31,61,31,61,30,179,31,179,30,254,31,221,31,45,31,119,31,165,31,67,31,78,31,176,31,235,31,19,31,86,31,95,31,170,31,170,30,118,31,118,30,89,31,47,31,47,30,127,31,127,30,3,31,3,30,129,31,79,31,202,31,205,31,28,31,51,31,79,31,198,31,190,31,190,30,81,31,65,31,101,31,88,31,88,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
