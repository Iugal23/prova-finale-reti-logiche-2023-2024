-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 244;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,65,0,0,0,251,0,108,0,119,0,241,0,242,0,80,0,18,0,71,0,0,0,0,0,0,0,218,0,109,0,152,0,6,0,179,0,45,0,131,0,0,0,163,0,10,0,243,0,0,0,202,0,0,0,157,0,131,0,92,0,34,0,170,0,0,0,243,0,241,0,164,0,0,0,176,0,173,0,216,0,0,0,210,0,0,0,223,0,178,0,187,0,69,0,0,0,15,0,16,0,83,0,0,0,47,0,233,0,76,0,113,0,180,0,7,0,201,0,77,0,52,0,115,0,19,0,169,0,249,0,61,0,238,0,220,0,45,0,201,0,132,0,80,0,0,0,23,0,55,0,184,0,16,0,115,0,55,0,0,0,116,0,29,0,100,0,176,0,177,0,183,0,137,0,193,0,48,0,254,0,80,0,201,0,180,0,136,0,59,0,85,0,233,0,138,0,52,0,101,0,62,0,238,0,95,0,0,0,0,0,143,0,0,0,83,0,82,0,93,0,51,0,15,0,32,0,0,0,0,0,197,0,234,0,167,0,171,0,0,0,24,0,10,0,0,0,103,0,199,0,75,0,75,0,64,0,0,0,44,0,147,0,0,0,159,0,229,0,125,0,27,0,42,0,43,0,151,0,0,0,0,0,183,0,185,0,0,0,50,0,97,0,33,0,99,0,114,0,181,0,20,0,0,0,210,0,170,0,197,0,0,0,235,0,187,0,18,0,202,0,101,0,77,0,210,0,118,0,217,0,186,0,12,0,23,0,0,0,0,0,126,0,107,0,0,0,86,0,0,0,26,0,178,0,218,0,13,0,29,0,0,0,117,0,206,0,0,0,101,0,250,0,0,0,74,0,227,0,0,0,0,0,63,0,30,0,246,0,37,0,39,0,80,0,17,0,120,0,175,0,0,0,20,0,62,0,7,0,0,0,117,0,66,0,191,0,101,0,149,0,0,0,96,0,0,0,146,0,193,0,176,0,155,0,116,0,101,0,213,0,213,0,31,0,19,0,199,0,0,0,0,0,240,0,55,0,0,0,115,0,0,0,91,0,116,0,0,0,0,0,0,0,118,0,105,0,52,0,103,0,102,0,162,0,30,0);
signal scenario_full  : scenario_type := (0,0,65,31,65,30,251,31,108,31,119,31,241,31,242,31,80,31,18,31,71,31,71,30,71,29,71,28,218,31,109,31,152,31,6,31,179,31,45,31,131,31,131,30,163,31,10,31,243,31,243,30,202,31,202,30,157,31,131,31,92,31,34,31,170,31,170,30,243,31,241,31,164,31,164,30,176,31,173,31,216,31,216,30,210,31,210,30,223,31,178,31,187,31,69,31,69,30,15,31,16,31,83,31,83,30,47,31,233,31,76,31,113,31,180,31,7,31,201,31,77,31,52,31,115,31,19,31,169,31,249,31,61,31,238,31,220,31,45,31,201,31,132,31,80,31,80,30,23,31,55,31,184,31,16,31,115,31,55,31,55,30,116,31,29,31,100,31,176,31,177,31,183,31,137,31,193,31,48,31,254,31,80,31,201,31,180,31,136,31,59,31,85,31,233,31,138,31,52,31,101,31,62,31,238,31,95,31,95,30,95,29,143,31,143,30,83,31,82,31,93,31,51,31,15,31,32,31,32,30,32,29,197,31,234,31,167,31,171,31,171,30,24,31,10,31,10,30,103,31,199,31,75,31,75,31,64,31,64,30,44,31,147,31,147,30,159,31,229,31,125,31,27,31,42,31,43,31,151,31,151,30,151,29,183,31,185,31,185,30,50,31,97,31,33,31,99,31,114,31,181,31,20,31,20,30,210,31,170,31,197,31,197,30,235,31,187,31,18,31,202,31,101,31,77,31,210,31,118,31,217,31,186,31,12,31,23,31,23,30,23,29,126,31,107,31,107,30,86,31,86,30,26,31,178,31,218,31,13,31,29,31,29,30,117,31,206,31,206,30,101,31,250,31,250,30,74,31,227,31,227,30,227,29,63,31,30,31,246,31,37,31,39,31,80,31,17,31,120,31,175,31,175,30,20,31,62,31,7,31,7,30,117,31,66,31,191,31,101,31,149,31,149,30,96,31,96,30,146,31,193,31,176,31,155,31,116,31,101,31,213,31,213,31,31,31,19,31,199,31,199,30,199,29,240,31,55,31,55,30,115,31,115,30,91,31,116,31,116,30,116,29,116,28,118,31,105,31,52,31,103,31,102,31,162,31,30,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
