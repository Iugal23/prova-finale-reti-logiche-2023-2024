-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 635;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (72,0,142,0,115,0,224,0,80,0,0,0,144,0,132,0,65,0,0,0,0,0,219,0,26,0,98,0,22,0,3,0,212,0,0,0,187,0,168,0,0,0,0,0,94,0,4,0,115,0,168,0,190,0,222,0,110,0,115,0,0,0,0,0,184,0,122,0,231,0,0,0,39,0,68,0,151,0,47,0,28,0,79,0,180,0,166,0,4,0,96,0,0,0,254,0,0,0,158,0,171,0,0,0,1,0,238,0,0,0,11,0,84,0,0,0,60,0,47,0,144,0,78,0,200,0,95,0,144,0,10,0,0,0,20,0,231,0,0,0,93,0,191,0,127,0,117,0,94,0,0,0,102,0,10,0,34,0,0,0,83,0,53,0,203,0,160,0,69,0,126,0,0,0,35,0,209,0,129,0,216,0,39,0,226,0,248,0,42,0,85,0,142,0,174,0,0,0,0,0,169,0,96,0,187,0,0,0,194,0,68,0,95,0,80,0,187,0,72,0,255,0,130,0,0,0,232,0,216,0,0,0,0,0,238,0,154,0,50,0,202,0,81,0,0,0,0,0,26,0,198,0,0,0,68,0,227,0,99,0,0,0,18,0,0,0,0,0,0,0,0,0,90,0,46,0,123,0,26,0,58,0,0,0,0,0,104,0,16,0,89,0,179,0,27,0,45,0,120,0,242,0,0,0,39,0,0,0,0,0,203,0,134,0,105,0,9,0,79,0,0,0,10,0,152,0,34,0,0,0,78,0,66,0,242,0,0,0,93,0,115,0,169,0,157,0,109,0,67,0,0,0,54,0,93,0,28,0,242,0,65,0,0,0,4,0,250,0,0,0,75,0,0,0,110,0,0,0,0,0,5,0,176,0,144,0,169,0,252,0,0,0,129,0,210,0,0,0,82,0,77,0,161,0,0,0,133,0,12,0,80,0,0,0,142,0,52,0,213,0,5,0,0,0,168,0,181,0,241,0,130,0,226,0,236,0,239,0,27,0,94,0,157,0,33,0,30,0,252,0,163,0,0,0,133,0,0,0,65,0,55,0,33,0,192,0,0,0,149,0,0,0,85,0,100,0,212,0,153,0,211,0,239,0,9,0,97,0,17,0,17,0,30,0,43,0,71,0,84,0,0,0,213,0,0,0,194,0,0,0,0,0,249,0,0,0,0,0,249,0,0,0,238,0,0,0,201,0,229,0,0,0,138,0,238,0,219,0,81,0,106,0,0,0,238,0,137,0,220,0,240,0,115,0,95,0,78,0,71,0,153,0,205,0,137,0,0,0,0,0,197,0,209,0,253,0,0,0,7,0,255,0,191,0,117,0,209,0,102,0,220,0,118,0,199,0,142,0,0,0,225,0,52,0,0,0,0,0,0,0,184,0,0,0,190,0,105,0,172,0,238,0,242,0,0,0,230,0,53,0,0,0,0,0,221,0,248,0,0,0,72,0,72,0,241,0,211,0,137,0,86,0,89,0,205,0,0,0,5,0,212,0,44,0,34,0,204,0,12,0,180,0,83,0,161,0,51,0,0,0,0,0,165,0,60,0,170,0,207,0,202,0,137,0,13,0,138,0,226,0,0,0,0,0,34,0,26,0,9,0,0,0,0,0,58,0,6,0,0,0,0,0,115,0,0,0,0,0,204,0,58,0,14,0,229,0,63,0,0,0,245,0,89,0,0,0,115,0,35,0,197,0,144,0,0,0,96,0,202,0,253,0,0,0,79,0,45,0,47,0,182,0,209,0,0,0,233,0,34,0,180,0,0,0,162,0,11,0,0,0,0,0,120,0,121,0,219,0,0,0,214,0,117,0,219,0,0,0,203,0,143,0,186,0,0,0,0,0,203,0,0,0,94,0,178,0,253,0,211,0,110,0,0,0,205,0,104,0,207,0,0,0,202,0,252,0,129,0,0,0,127,0,118,0,0,0,74,0,0,0,243,0,31,0,0,0,136,0,91,0,38,0,145,0,0,0,150,0,218,0,217,0,201,0,214,0,157,0,76,0,150,0,182,0,137,0,2,0,208,0,210,0,11,0,237,0,162,0,36,0,98,0,181,0,20,0,34,0,84,0,106,0,80,0,0,0,228,0,45,0,81,0,107,0,130,0,155,0,155,0,73,0,46,0,61,0,16,0,0,0,212,0,140,0,149,0,94,0,44,0,44,0,255,0,4,0,16,0,124,0,97,0,69,0,220,0,0,0,0,0,0,0,111,0,0,0,229,0,190,0,142,0,170,0,0,0,146,0,0,0,117,0,0,0,80,0,233,0,194,0,163,0,0,0,111,0,0,0,178,0,194,0,213,0,252,0,0,0,112,0,241,0,32,0,248,0,110,0,106,0,158,0,151,0,69,0,195,0,150,0,206,0,146,0,181,0,137,0,175,0,0,0,93,0,168,0,132,0,211,0,55,0,167,0,202,0,181,0,61,0,193,0,134,0,0,0,0,0,53,0,58,0,104,0,0,0,180,0,0,0,0,0,16,0,0,0,0,0,0,0,240,0,201,0,0,0,0,0,98,0,17,0,142,0,151,0,0,0,202,0,33,0,124,0,89,0,87,0,212,0,0,0,86,0,217,0,202,0,119,0,9,0,0,0,0,0,181,0,124,0,12,0,164,0,254,0,25,0,0,0,0,0,253,0,0,0,237,0,198,0,0,0,0,0,0,0,0,0,0,0,0,0,225,0,58,0,104,0,102,0,27,0,69,0,0,0,190,0,0,0,87,0,56,0,251,0,59,0,48,0,169,0,0,0,0,0,250,0,144,0,155,0,62,0,7,0,151,0,202,0,44,0,0,0,0,0,0,0,0,0,31,0,142,0,75,0,0,0,204,0,91,0,149,0,0,0,129,0,227,0);
signal scenario_full  : scenario_type := (72,31,142,31,115,31,224,31,80,31,80,30,144,31,132,31,65,31,65,30,65,29,219,31,26,31,98,31,22,31,3,31,212,31,212,30,187,31,168,31,168,30,168,29,94,31,4,31,115,31,168,31,190,31,222,31,110,31,115,31,115,30,115,29,184,31,122,31,231,31,231,30,39,31,68,31,151,31,47,31,28,31,79,31,180,31,166,31,4,31,96,31,96,30,254,31,254,30,158,31,171,31,171,30,1,31,238,31,238,30,11,31,84,31,84,30,60,31,47,31,144,31,78,31,200,31,95,31,144,31,10,31,10,30,20,31,231,31,231,30,93,31,191,31,127,31,117,31,94,31,94,30,102,31,10,31,34,31,34,30,83,31,53,31,203,31,160,31,69,31,126,31,126,30,35,31,209,31,129,31,216,31,39,31,226,31,248,31,42,31,85,31,142,31,174,31,174,30,174,29,169,31,96,31,187,31,187,30,194,31,68,31,95,31,80,31,187,31,72,31,255,31,130,31,130,30,232,31,216,31,216,30,216,29,238,31,154,31,50,31,202,31,81,31,81,30,81,29,26,31,198,31,198,30,68,31,227,31,99,31,99,30,18,31,18,30,18,29,18,28,18,27,90,31,46,31,123,31,26,31,58,31,58,30,58,29,104,31,16,31,89,31,179,31,27,31,45,31,120,31,242,31,242,30,39,31,39,30,39,29,203,31,134,31,105,31,9,31,79,31,79,30,10,31,152,31,34,31,34,30,78,31,66,31,242,31,242,30,93,31,115,31,169,31,157,31,109,31,67,31,67,30,54,31,93,31,28,31,242,31,65,31,65,30,4,31,250,31,250,30,75,31,75,30,110,31,110,30,110,29,5,31,176,31,144,31,169,31,252,31,252,30,129,31,210,31,210,30,82,31,77,31,161,31,161,30,133,31,12,31,80,31,80,30,142,31,52,31,213,31,5,31,5,30,168,31,181,31,241,31,130,31,226,31,236,31,239,31,27,31,94,31,157,31,33,31,30,31,252,31,163,31,163,30,133,31,133,30,65,31,55,31,33,31,192,31,192,30,149,31,149,30,85,31,100,31,212,31,153,31,211,31,239,31,9,31,97,31,17,31,17,31,30,31,43,31,71,31,84,31,84,30,213,31,213,30,194,31,194,30,194,29,249,31,249,30,249,29,249,31,249,30,238,31,238,30,201,31,229,31,229,30,138,31,238,31,219,31,81,31,106,31,106,30,238,31,137,31,220,31,240,31,115,31,95,31,78,31,71,31,153,31,205,31,137,31,137,30,137,29,197,31,209,31,253,31,253,30,7,31,255,31,191,31,117,31,209,31,102,31,220,31,118,31,199,31,142,31,142,30,225,31,52,31,52,30,52,29,52,28,184,31,184,30,190,31,105,31,172,31,238,31,242,31,242,30,230,31,53,31,53,30,53,29,221,31,248,31,248,30,72,31,72,31,241,31,211,31,137,31,86,31,89,31,205,31,205,30,5,31,212,31,44,31,34,31,204,31,12,31,180,31,83,31,161,31,51,31,51,30,51,29,165,31,60,31,170,31,207,31,202,31,137,31,13,31,138,31,226,31,226,30,226,29,34,31,26,31,9,31,9,30,9,29,58,31,6,31,6,30,6,29,115,31,115,30,115,29,204,31,58,31,14,31,229,31,63,31,63,30,245,31,89,31,89,30,115,31,35,31,197,31,144,31,144,30,96,31,202,31,253,31,253,30,79,31,45,31,47,31,182,31,209,31,209,30,233,31,34,31,180,31,180,30,162,31,11,31,11,30,11,29,120,31,121,31,219,31,219,30,214,31,117,31,219,31,219,30,203,31,143,31,186,31,186,30,186,29,203,31,203,30,94,31,178,31,253,31,211,31,110,31,110,30,205,31,104,31,207,31,207,30,202,31,252,31,129,31,129,30,127,31,118,31,118,30,74,31,74,30,243,31,31,31,31,30,136,31,91,31,38,31,145,31,145,30,150,31,218,31,217,31,201,31,214,31,157,31,76,31,150,31,182,31,137,31,2,31,208,31,210,31,11,31,237,31,162,31,36,31,98,31,181,31,20,31,34,31,84,31,106,31,80,31,80,30,228,31,45,31,81,31,107,31,130,31,155,31,155,31,73,31,46,31,61,31,16,31,16,30,212,31,140,31,149,31,94,31,44,31,44,31,255,31,4,31,16,31,124,31,97,31,69,31,220,31,220,30,220,29,220,28,111,31,111,30,229,31,190,31,142,31,170,31,170,30,146,31,146,30,117,31,117,30,80,31,233,31,194,31,163,31,163,30,111,31,111,30,178,31,194,31,213,31,252,31,252,30,112,31,241,31,32,31,248,31,110,31,106,31,158,31,151,31,69,31,195,31,150,31,206,31,146,31,181,31,137,31,175,31,175,30,93,31,168,31,132,31,211,31,55,31,167,31,202,31,181,31,61,31,193,31,134,31,134,30,134,29,53,31,58,31,104,31,104,30,180,31,180,30,180,29,16,31,16,30,16,29,16,28,240,31,201,31,201,30,201,29,98,31,17,31,142,31,151,31,151,30,202,31,33,31,124,31,89,31,87,31,212,31,212,30,86,31,217,31,202,31,119,31,9,31,9,30,9,29,181,31,124,31,12,31,164,31,254,31,25,31,25,30,25,29,253,31,253,30,237,31,198,31,198,30,198,29,198,28,198,27,198,26,198,25,225,31,58,31,104,31,102,31,27,31,69,31,69,30,190,31,190,30,87,31,56,31,251,31,59,31,48,31,169,31,169,30,169,29,250,31,144,31,155,31,62,31,7,31,151,31,202,31,44,31,44,30,44,29,44,28,44,27,31,31,142,31,75,31,75,30,204,31,91,31,149,31,149,30,129,31,227,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
