-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 935;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (204,0,228,0,99,0,30,0,168,0,190,0,29,0,237,0,216,0,76,0,90,0,29,0,26,0,252,0,102,0,0,0,239,0,0,0,235,0,44,0,48,0,13,0,0,0,168,0,166,0,183,0,175,0,44,0,253,0,68,0,234,0,94,0,251,0,144,0,7,0,46,0,26,0,16,0,65,0,121,0,0,0,200,0,25,0,189,0,89,0,0,0,233,0,212,0,26,0,124,0,17,0,153,0,230,0,0,0,0,0,207,0,140,0,117,0,193,0,0,0,111,0,95,0,0,0,79,0,99,0,0,0,0,0,132,0,124,0,166,0,239,0,0,0,30,0,0,0,95,0,0,0,27,0,241,0,0,0,237,0,0,0,149,0,145,0,238,0,232,0,0,0,50,0,198,0,221,0,153,0,87,0,0,0,215,0,214,0,18,0,1,0,155,0,87,0,113,0,160,0,32,0,231,0,80,0,75,0,0,0,206,0,175,0,0,0,218,0,0,0,0,0,89,0,76,0,142,0,41,0,0,0,143,0,78,0,161,0,0,0,195,0,208,0,36,0,238,0,158,0,154,0,34,0,23,0,0,0,219,0,38,0,218,0,94,0,14,0,88,0,0,0,245,0,0,0,15,0,232,0,100,0,97,0,0,0,160,0,0,0,94,0,185,0,192,0,93,0,238,0,77,0,106,0,0,0,0,0,176,0,0,0,0,0,0,0,68,0,236,0,110,0,0,0,225,0,56,0,18,0,0,0,0,0,134,0,147,0,0,0,123,0,160,0,206,0,102,0,253,0,166,0,0,0,155,0,150,0,218,0,89,0,250,0,85,0,0,0,220,0,34,0,0,0,140,0,135,0,178,0,254,0,175,0,41,0,206,0,0,0,0,0,198,0,184,0,0,0,67,0,158,0,224,0,50,0,161,0,0,0,0,0,252,0,234,0,0,0,152,0,28,0,208,0,0,0,98,0,138,0,217,0,128,0,0,0,221,0,78,0,0,0,197,0,204,0,0,0,0,0,167,0,40,0,26,0,174,0,225,0,81,0,91,0,235,0,164,0,0,0,0,0,166,0,191,0,0,0,153,0,75,0,9,0,232,0,233,0,0,0,164,0,0,0,0,0,229,0,126,0,245,0,199,0,133,0,167,0,202,0,147,0,2,0,0,0,122,0,82,0,41,0,83,0,0,0,181,0,238,0,0,0,216,0,202,0,93,0,150,0,101,0,41,0,0,0,0,0,210,0,46,0,62,0,50,0,247,0,177,0,56,0,164,0,81,0,0,0,163,0,0,0,68,0,104,0,221,0,0,0,217,0,0,0,222,0,19,0,18,0,194,0,53,0,235,0,255,0,197,0,140,0,0,0,60,0,122,0,229,0,94,0,63,0,23,0,0,0,110,0,193,0,0,0,0,0,41,0,0,0,52,0,148,0,0,0,236,0,215,0,83,0,183,0,174,0,90,0,39,0,55,0,0,0,86,0,160,0,187,0,18,0,238,0,241,0,225,0,85,0,0,0,202,0,151,0,196,0,231,0,43,0,217,0,0,0,253,0,82,0,159,0,247,0,116,0,26,0,52,0,108,0,93,0,9,0,184,0,180,0,204,0,162,0,95,0,0,0,229,0,3,0,68,0,0,0,82,0,185,0,229,0,12,0,56,0,137,0,0,0,0,0,210,0,123,0,0,0,22,0,208,0,18,0,0,0,0,0,214,0,148,0,215,0,186,0,105,0,84,0,250,0,65,0,40,0,79,0,29,0,208,0,89,0,253,0,118,0,236,0,24,0,36,0,0,0,139,0,32,0,149,0,158,0,220,0,0,0,218,0,69,0,226,0,147,0,33,0,0,0,158,0,150,0,52,0,0,0,143,0,94,0,0,0,96,0,144,0,0,0,151,0,175,0,66,0,66,0,4,0,189,0,107,0,16,0,0,0,36,0,160,0,124,0,203,0,37,0,204,0,3,0,0,0,103,0,0,0,22,0,236,0,163,0,84,0,0,0,43,0,166,0,91,0,0,0,0,0,57,0,0,0,99,0,0,0,36,0,227,0,15,0,27,0,161,0,192,0,222,0,0,0,0,0,0,0,26,0,227,0,189,0,97,0,0,0,211,0,123,0,191,0,0,0,0,0,78,0,81,0,0,0,0,0,152,0,175,0,28,0,183,0,159,0,246,0,49,0,90,0,202,0,138,0,0,0,239,0,121,0,176,0,106,0,200,0,139,0,138,0,0,0,0,0,0,0,0,0,108,0,150,0,172,0,228,0,231,0,205,0,137,0,0,0,36,0,42,0,97,0,0,0,197,0,0,0,0,0,231,0,204,0,161,0,184,0,0,0,99,0,123,0,188,0,87,0,178,0,0,0,201,0,246,0,62,0,49,0,79,0,215,0,77,0,5,0,173,0,162,0,43,0,167,0,0,0,189,0,243,0,110,0,34,0,238,0,111,0,64,0,109,0,83,0,77,0,184,0,0,0,26,0,186,0,175,0,40,0,97,0,206,0,116,0,0,0,35,0,119,0,215,0,239,0,107,0,194,0,40,0,110,0,27,0,154,0,60,0,218,0,183,0,38,0,40,0,126,0,155,0,158,0,0,0,0,0,0,0,37,0,0,0,232,0,0,0,122,0,58,0,0,0,202,0,111,0,0,0,0,0,156,0,178,0,51,0,243,0,85,0,0,0,1,0,178,0,249,0,3,0,199,0,239,0,86,0,105,0,213,0,0,0,36,0,0,0,0,0,0,0,233,0,62,0,108,0,190,0,67,0,0,0,14,0,219,0,22,0,0,0,142,0,242,0,119,0,0,0,155,0,0,0,138,0,214,0,0,0,0,0,187,0,0,0,0,0,94,0,217,0,151,0,0,0,41,0,72,0,0,0,215,0,0,0,55,0,44,0,20,0,189,0,97,0,199,0,178,0,17,0,95,0,57,0,63,0,129,0,76,0,127,0,183,0,0,0,0,0,96,0,51,0,117,0,14,0,126,0,0,0,175,0,0,0,142,0,248,0,65,0,90,0,121,0,0,0,79,0,89,0,97,0,0,0,163,0,11,0,64,0,84,0,159,0,220,0,242,0,0,0,222,0,40,0,251,0,170,0,0,0,0,0,251,0,115,0,29,0,0,0,155,0,121,0,59,0,182,0,0,0,114,0,137,0,86,0,213,0,136,0,86,0,151,0,128,0,249,0,155,0,77,0,211,0,0,0,246,0,119,0,58,0,152,0,245,0,151,0,64,0,0,0,167,0,243,0,97,0,97,0,207,0,153,0,0,0,184,0,159,0,26,0,46,0,59,0,140,0,133,0,78,0,0,0,0,0,212,0,121,0,0,0,92,0,59,0,100,0,78,0,87,0,0,0,0,0,150,0,32,0,206,0,161,0,0,0,0,0,161,0,0,0,131,0,40,0,5,0,119,0,85,0,83,0,210,0,0,0,64,0,222,0,120,0,41,0,98,0,69,0,73,0,100,0,86,0,0,0,108,0,170,0,209,0,179,0,0,0,202,0,198,0,60,0,85,0,178,0,125,0,0,0,178,0,0,0,143,0,0,0,122,0,73,0,122,0,133,0,0,0,59,0,110,0,217,0,187,0,110,0,222,0,83,0,208,0,0,0,4,0,131,0,0,0,32,0,226,0,236,0,77,0,156,0,110,0,185,0,0,0,0,0,114,0,146,0,241,0,86,0,122,0,206,0,17,0,164,0,125,0,169,0,0,0,175,0,181,0,84,0,0,0,224,0,111,0,0,0,65,0,26,0,84,0,0,0,0,0,233,0,0,0,112,0,60,0,0,0,33,0,175,0,254,0,120,0,40,0,150,0,42,0,112,0,187,0,183,0,0,0,59,0,166,0,246,0,242,0,0,0,0,0,150,0,190,0,225,0,43,0,227,0,0,0,0,0,218,0,103,0,129,0,21,0,176,0,117,0,206,0,102,0,24,0,16,0,0,0,6,0,23,0,2,0,198,0,102,0,67,0,0,0,153,0,152,0,0,0,5,0,226,0,0,0,141,0,76,0,119,0,236,0,0,0,243,0,94,0,188,0,0,0,9,0,66,0,216,0,175,0,180,0,0,0,213,0,52,0,111,0,183,0,212,0,163,0,0,0,153,0,251,0,32,0,200,0,56,0,0,0,185,0,9,0,25,0,165,0,159,0,222,0,254,0,66,0,164,0,0,0,68,0,55,0,0,0,251,0,77,0);
signal scenario_full  : scenario_type := (204,31,228,31,99,31,30,31,168,31,190,31,29,31,237,31,216,31,76,31,90,31,29,31,26,31,252,31,102,31,102,30,239,31,239,30,235,31,44,31,48,31,13,31,13,30,168,31,166,31,183,31,175,31,44,31,253,31,68,31,234,31,94,31,251,31,144,31,7,31,46,31,26,31,16,31,65,31,121,31,121,30,200,31,25,31,189,31,89,31,89,30,233,31,212,31,26,31,124,31,17,31,153,31,230,31,230,30,230,29,207,31,140,31,117,31,193,31,193,30,111,31,95,31,95,30,79,31,99,31,99,30,99,29,132,31,124,31,166,31,239,31,239,30,30,31,30,30,95,31,95,30,27,31,241,31,241,30,237,31,237,30,149,31,145,31,238,31,232,31,232,30,50,31,198,31,221,31,153,31,87,31,87,30,215,31,214,31,18,31,1,31,155,31,87,31,113,31,160,31,32,31,231,31,80,31,75,31,75,30,206,31,175,31,175,30,218,31,218,30,218,29,89,31,76,31,142,31,41,31,41,30,143,31,78,31,161,31,161,30,195,31,208,31,36,31,238,31,158,31,154,31,34,31,23,31,23,30,219,31,38,31,218,31,94,31,14,31,88,31,88,30,245,31,245,30,15,31,232,31,100,31,97,31,97,30,160,31,160,30,94,31,185,31,192,31,93,31,238,31,77,31,106,31,106,30,106,29,176,31,176,30,176,29,176,28,68,31,236,31,110,31,110,30,225,31,56,31,18,31,18,30,18,29,134,31,147,31,147,30,123,31,160,31,206,31,102,31,253,31,166,31,166,30,155,31,150,31,218,31,89,31,250,31,85,31,85,30,220,31,34,31,34,30,140,31,135,31,178,31,254,31,175,31,41,31,206,31,206,30,206,29,198,31,184,31,184,30,67,31,158,31,224,31,50,31,161,31,161,30,161,29,252,31,234,31,234,30,152,31,28,31,208,31,208,30,98,31,138,31,217,31,128,31,128,30,221,31,78,31,78,30,197,31,204,31,204,30,204,29,167,31,40,31,26,31,174,31,225,31,81,31,91,31,235,31,164,31,164,30,164,29,166,31,191,31,191,30,153,31,75,31,9,31,232,31,233,31,233,30,164,31,164,30,164,29,229,31,126,31,245,31,199,31,133,31,167,31,202,31,147,31,2,31,2,30,122,31,82,31,41,31,83,31,83,30,181,31,238,31,238,30,216,31,202,31,93,31,150,31,101,31,41,31,41,30,41,29,210,31,46,31,62,31,50,31,247,31,177,31,56,31,164,31,81,31,81,30,163,31,163,30,68,31,104,31,221,31,221,30,217,31,217,30,222,31,19,31,18,31,194,31,53,31,235,31,255,31,197,31,140,31,140,30,60,31,122,31,229,31,94,31,63,31,23,31,23,30,110,31,193,31,193,30,193,29,41,31,41,30,52,31,148,31,148,30,236,31,215,31,83,31,183,31,174,31,90,31,39,31,55,31,55,30,86,31,160,31,187,31,18,31,238,31,241,31,225,31,85,31,85,30,202,31,151,31,196,31,231,31,43,31,217,31,217,30,253,31,82,31,159,31,247,31,116,31,26,31,52,31,108,31,93,31,9,31,184,31,180,31,204,31,162,31,95,31,95,30,229,31,3,31,68,31,68,30,82,31,185,31,229,31,12,31,56,31,137,31,137,30,137,29,210,31,123,31,123,30,22,31,208,31,18,31,18,30,18,29,214,31,148,31,215,31,186,31,105,31,84,31,250,31,65,31,40,31,79,31,29,31,208,31,89,31,253,31,118,31,236,31,24,31,36,31,36,30,139,31,32,31,149,31,158,31,220,31,220,30,218,31,69,31,226,31,147,31,33,31,33,30,158,31,150,31,52,31,52,30,143,31,94,31,94,30,96,31,144,31,144,30,151,31,175,31,66,31,66,31,4,31,189,31,107,31,16,31,16,30,36,31,160,31,124,31,203,31,37,31,204,31,3,31,3,30,103,31,103,30,22,31,236,31,163,31,84,31,84,30,43,31,166,31,91,31,91,30,91,29,57,31,57,30,99,31,99,30,36,31,227,31,15,31,27,31,161,31,192,31,222,31,222,30,222,29,222,28,26,31,227,31,189,31,97,31,97,30,211,31,123,31,191,31,191,30,191,29,78,31,81,31,81,30,81,29,152,31,175,31,28,31,183,31,159,31,246,31,49,31,90,31,202,31,138,31,138,30,239,31,121,31,176,31,106,31,200,31,139,31,138,31,138,30,138,29,138,28,138,27,108,31,150,31,172,31,228,31,231,31,205,31,137,31,137,30,36,31,42,31,97,31,97,30,197,31,197,30,197,29,231,31,204,31,161,31,184,31,184,30,99,31,123,31,188,31,87,31,178,31,178,30,201,31,246,31,62,31,49,31,79,31,215,31,77,31,5,31,173,31,162,31,43,31,167,31,167,30,189,31,243,31,110,31,34,31,238,31,111,31,64,31,109,31,83,31,77,31,184,31,184,30,26,31,186,31,175,31,40,31,97,31,206,31,116,31,116,30,35,31,119,31,215,31,239,31,107,31,194,31,40,31,110,31,27,31,154,31,60,31,218,31,183,31,38,31,40,31,126,31,155,31,158,31,158,30,158,29,158,28,37,31,37,30,232,31,232,30,122,31,58,31,58,30,202,31,111,31,111,30,111,29,156,31,178,31,51,31,243,31,85,31,85,30,1,31,178,31,249,31,3,31,199,31,239,31,86,31,105,31,213,31,213,30,36,31,36,30,36,29,36,28,233,31,62,31,108,31,190,31,67,31,67,30,14,31,219,31,22,31,22,30,142,31,242,31,119,31,119,30,155,31,155,30,138,31,214,31,214,30,214,29,187,31,187,30,187,29,94,31,217,31,151,31,151,30,41,31,72,31,72,30,215,31,215,30,55,31,44,31,20,31,189,31,97,31,199,31,178,31,17,31,95,31,57,31,63,31,129,31,76,31,127,31,183,31,183,30,183,29,96,31,51,31,117,31,14,31,126,31,126,30,175,31,175,30,142,31,248,31,65,31,90,31,121,31,121,30,79,31,89,31,97,31,97,30,163,31,11,31,64,31,84,31,159,31,220,31,242,31,242,30,222,31,40,31,251,31,170,31,170,30,170,29,251,31,115,31,29,31,29,30,155,31,121,31,59,31,182,31,182,30,114,31,137,31,86,31,213,31,136,31,86,31,151,31,128,31,249,31,155,31,77,31,211,31,211,30,246,31,119,31,58,31,152,31,245,31,151,31,64,31,64,30,167,31,243,31,97,31,97,31,207,31,153,31,153,30,184,31,159,31,26,31,46,31,59,31,140,31,133,31,78,31,78,30,78,29,212,31,121,31,121,30,92,31,59,31,100,31,78,31,87,31,87,30,87,29,150,31,32,31,206,31,161,31,161,30,161,29,161,31,161,30,131,31,40,31,5,31,119,31,85,31,83,31,210,31,210,30,64,31,222,31,120,31,41,31,98,31,69,31,73,31,100,31,86,31,86,30,108,31,170,31,209,31,179,31,179,30,202,31,198,31,60,31,85,31,178,31,125,31,125,30,178,31,178,30,143,31,143,30,122,31,73,31,122,31,133,31,133,30,59,31,110,31,217,31,187,31,110,31,222,31,83,31,208,31,208,30,4,31,131,31,131,30,32,31,226,31,236,31,77,31,156,31,110,31,185,31,185,30,185,29,114,31,146,31,241,31,86,31,122,31,206,31,17,31,164,31,125,31,169,31,169,30,175,31,181,31,84,31,84,30,224,31,111,31,111,30,65,31,26,31,84,31,84,30,84,29,233,31,233,30,112,31,60,31,60,30,33,31,175,31,254,31,120,31,40,31,150,31,42,31,112,31,187,31,183,31,183,30,59,31,166,31,246,31,242,31,242,30,242,29,150,31,190,31,225,31,43,31,227,31,227,30,227,29,218,31,103,31,129,31,21,31,176,31,117,31,206,31,102,31,24,31,16,31,16,30,6,31,23,31,2,31,198,31,102,31,67,31,67,30,153,31,152,31,152,30,5,31,226,31,226,30,141,31,76,31,119,31,236,31,236,30,243,31,94,31,188,31,188,30,9,31,66,31,216,31,175,31,180,31,180,30,213,31,52,31,111,31,183,31,212,31,163,31,163,30,153,31,251,31,32,31,200,31,56,31,56,30,185,31,9,31,25,31,165,31,159,31,222,31,254,31,66,31,164,31,164,30,68,31,55,31,55,30,251,31,77,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
