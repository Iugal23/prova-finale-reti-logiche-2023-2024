-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_468 is
end project_tb_468;

architecture project_tb_arch_468 of project_tb_468 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 589;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (153,0,150,0,0,0,214,0,0,0,76,0,106,0,48,0,208,0,159,0,0,0,65,0,151,0,0,0,0,0,254,0,151,0,175,0,24,0,28,0,83,0,184,0,231,0,230,0,138,0,184,0,42,0,0,0,216,0,0,0,174,0,26,0,92,0,0,0,118,0,0,0,40,0,0,0,154,0,0,0,0,0,192,0,88,0,124,0,235,0,0,0,136,0,218,0,17,0,5,0,0,0,0,0,160,0,247,0,107,0,170,0,111,0,63,0,3,0,129,0,0,0,0,0,58,0,0,0,54,0,82,0,0,0,109,0,0,0,71,0,63,0,89,0,140,0,112,0,175,0,21,0,200,0,176,0,11,0,0,0,128,0,31,0,23,0,241,0,81,0,3,0,166,0,0,0,53,0,68,0,234,0,77,0,243,0,125,0,0,0,0,0,68,0,0,0,217,0,0,0,32,0,54,0,0,0,26,0,173,0,78,0,39,0,151,0,0,0,253,0,202,0,166,0,124,0,24,0,148,0,233,0,113,0,77,0,23,0,225,0,54,0,17,0,0,0,13,0,235,0,0,0,203,0,89,0,0,0,78,0,0,0,234,0,180,0,0,0,84,0,242,0,0,0,0,0,249,0,64,0,0,0,0,0,0,0,0,0,236,0,242,0,188,0,228,0,0,0,240,0,171,0,127,0,0,0,0,0,100,0,0,0,221,0,214,0,120,0,144,0,0,0,35,0,74,0,33,0,250,0,204,0,6,0,231,0,14,0,99,0,53,0,127,0,79,0,44,0,167,0,0,0,83,0,62,0,67,0,214,0,148,0,61,0,0,0,20,0,142,0,4,0,223,0,67,0,235,0,72,0,170,0,69,0,161,0,148,0,0,0,0,0,51,0,0,0,2,0,208,0,222,0,0,0,253,0,33,0,176,0,68,0,240,0,197,0,34,0,208,0,0,0,0,0,245,0,191,0,0,0,80,0,0,0,0,0,56,0,24,0,241,0,0,0,20,0,0,0,81,0,0,0,138,0,235,0,188,0,192,0,36,0,104,0,65,0,221,0,194,0,203,0,10,0,22,0,209,0,131,0,0,0,62,0,57,0,46,0,101,0,27,0,167,0,0,0,0,0,182,0,29,0,21,0,0,0,185,0,199,0,42,0,167,0,15,0,49,0,240,0,39,0,171,0,74,0,147,0,214,0,131,0,165,0,15,0,0,0,28,0,91,0,0,0,69,0,0,0,177,0,191,0,95,0,47,0,0,0,15,0,22,0,0,0,97,0,123,0,238,0,99,0,163,0,0,0,0,0,132,0,141,0,228,0,99,0,228,0,55,0,73,0,227,0,69,0,177,0,0,0,191,0,156,0,26,0,214,0,221,0,0,0,109,0,10,0,169,0,234,0,1,0,10,0,56,0,60,0,230,0,0,0,0,0,134,0,0,0,80,0,0,0,175,0,1,0,230,0,46,0,120,0,120,0,151,0,140,0,0,0,0,0,234,0,216,0,181,0,76,0,195,0,150,0,102,0,41,0,158,0,152,0,247,0,29,0,141,0,7,0,0,0,89,0,72,0,0,0,28,0,60,0,0,0,20,0,200,0,136,0,35,0,126,0,207,0,90,0,141,0,216,0,15,0,168,0,192,0,23,0,158,0,4,0,79,0,112,0,122,0,224,0,130,0,140,0,0,0,166,0,50,0,0,0,39,0,48,0,0,0,10,0,145,0,0,0,53,0,0,0,81,0,166,0,38,0,175,0,166,0,194,0,50,0,152,0,93,0,227,0,0,0,56,0,51,0,71,0,0,0,181,0,66,0,184,0,35,0,213,0,152,0,190,0,7,0,59,0,99,0,194,0,252,0,102,0,0,0,0,0,182,0,148,0,169,0,203,0,47,0,7,0,206,0,100,0,9,0,48,0,95,0,63,0,0,0,71,0,200,0,0,0,0,0,29,0,16,0,76,0,0,0,246,0,54,0,0,0,155,0,233,0,0,0,11,0,94,0,38,0,0,0,109,0,0,0,0,0,10,0,159,0,35,0,167,0,7,0,181,0,76,0,155,0,8,0,168,0,153,0,165,0,238,0,82,0,5,0,82,0,103,0,0,0,209,0,59,0,94,0,0,0,212,0,94,0,21,0,0,0,158,0,23,0,116,0,0,0,49,0,81,0,7,0,121,0,114,0,120,0,94,0,63,0,0,0,14,0,122,0,141,0,0,0,21,0,114,0,92,0,83,0,14,0,107,0,201,0,140,0,179,0,235,0,156,0,248,0,0,0,142,0,210,0,0,0,109,0,253,0,118,0,187,0,0,0,176,0,182,0,54,0,75,0,222,0,44,0,24,0,0,0,0,0,233,0,0,0,137,0,62,0,144,0,161,0,123,0,186,0,26,0,93,0,146,0,0,0,70,0,121,0,230,0,116,0,175,0,67,0,109,0,91,0,0,0,144,0,241,0,59,0,129,0,251,0,200,0,0,0,61,0,178,0,11,0,0,0,68,0,215,0,250,0,95,0,151,0,157,0,218,0,139,0,128,0,96,0,175,0,223,0,112,0,192,0,0,0,0,0,218,0,227,0,33,0,7,0,196,0,0,0,255,0,165,0,162,0,71,0,0,0,204,0,187,0,116,0,183,0,31,0,170,0,0,0,0,0);
signal scenario_full  : scenario_type := (153,31,150,31,150,30,214,31,214,30,76,31,106,31,48,31,208,31,159,31,159,30,65,31,151,31,151,30,151,29,254,31,151,31,175,31,24,31,28,31,83,31,184,31,231,31,230,31,138,31,184,31,42,31,42,30,216,31,216,30,174,31,26,31,92,31,92,30,118,31,118,30,40,31,40,30,154,31,154,30,154,29,192,31,88,31,124,31,235,31,235,30,136,31,218,31,17,31,5,31,5,30,5,29,160,31,247,31,107,31,170,31,111,31,63,31,3,31,129,31,129,30,129,29,58,31,58,30,54,31,82,31,82,30,109,31,109,30,71,31,63,31,89,31,140,31,112,31,175,31,21,31,200,31,176,31,11,31,11,30,128,31,31,31,23,31,241,31,81,31,3,31,166,31,166,30,53,31,68,31,234,31,77,31,243,31,125,31,125,30,125,29,68,31,68,30,217,31,217,30,32,31,54,31,54,30,26,31,173,31,78,31,39,31,151,31,151,30,253,31,202,31,166,31,124,31,24,31,148,31,233,31,113,31,77,31,23,31,225,31,54,31,17,31,17,30,13,31,235,31,235,30,203,31,89,31,89,30,78,31,78,30,234,31,180,31,180,30,84,31,242,31,242,30,242,29,249,31,64,31,64,30,64,29,64,28,64,27,236,31,242,31,188,31,228,31,228,30,240,31,171,31,127,31,127,30,127,29,100,31,100,30,221,31,214,31,120,31,144,31,144,30,35,31,74,31,33,31,250,31,204,31,6,31,231,31,14,31,99,31,53,31,127,31,79,31,44,31,167,31,167,30,83,31,62,31,67,31,214,31,148,31,61,31,61,30,20,31,142,31,4,31,223,31,67,31,235,31,72,31,170,31,69,31,161,31,148,31,148,30,148,29,51,31,51,30,2,31,208,31,222,31,222,30,253,31,33,31,176,31,68,31,240,31,197,31,34,31,208,31,208,30,208,29,245,31,191,31,191,30,80,31,80,30,80,29,56,31,24,31,241,31,241,30,20,31,20,30,81,31,81,30,138,31,235,31,188,31,192,31,36,31,104,31,65,31,221,31,194,31,203,31,10,31,22,31,209,31,131,31,131,30,62,31,57,31,46,31,101,31,27,31,167,31,167,30,167,29,182,31,29,31,21,31,21,30,185,31,199,31,42,31,167,31,15,31,49,31,240,31,39,31,171,31,74,31,147,31,214,31,131,31,165,31,15,31,15,30,28,31,91,31,91,30,69,31,69,30,177,31,191,31,95,31,47,31,47,30,15,31,22,31,22,30,97,31,123,31,238,31,99,31,163,31,163,30,163,29,132,31,141,31,228,31,99,31,228,31,55,31,73,31,227,31,69,31,177,31,177,30,191,31,156,31,26,31,214,31,221,31,221,30,109,31,10,31,169,31,234,31,1,31,10,31,56,31,60,31,230,31,230,30,230,29,134,31,134,30,80,31,80,30,175,31,1,31,230,31,46,31,120,31,120,31,151,31,140,31,140,30,140,29,234,31,216,31,181,31,76,31,195,31,150,31,102,31,41,31,158,31,152,31,247,31,29,31,141,31,7,31,7,30,89,31,72,31,72,30,28,31,60,31,60,30,20,31,200,31,136,31,35,31,126,31,207,31,90,31,141,31,216,31,15,31,168,31,192,31,23,31,158,31,4,31,79,31,112,31,122,31,224,31,130,31,140,31,140,30,166,31,50,31,50,30,39,31,48,31,48,30,10,31,145,31,145,30,53,31,53,30,81,31,166,31,38,31,175,31,166,31,194,31,50,31,152,31,93,31,227,31,227,30,56,31,51,31,71,31,71,30,181,31,66,31,184,31,35,31,213,31,152,31,190,31,7,31,59,31,99,31,194,31,252,31,102,31,102,30,102,29,182,31,148,31,169,31,203,31,47,31,7,31,206,31,100,31,9,31,48,31,95,31,63,31,63,30,71,31,200,31,200,30,200,29,29,31,16,31,76,31,76,30,246,31,54,31,54,30,155,31,233,31,233,30,11,31,94,31,38,31,38,30,109,31,109,30,109,29,10,31,159,31,35,31,167,31,7,31,181,31,76,31,155,31,8,31,168,31,153,31,165,31,238,31,82,31,5,31,82,31,103,31,103,30,209,31,59,31,94,31,94,30,212,31,94,31,21,31,21,30,158,31,23,31,116,31,116,30,49,31,81,31,7,31,121,31,114,31,120,31,94,31,63,31,63,30,14,31,122,31,141,31,141,30,21,31,114,31,92,31,83,31,14,31,107,31,201,31,140,31,179,31,235,31,156,31,248,31,248,30,142,31,210,31,210,30,109,31,253,31,118,31,187,31,187,30,176,31,182,31,54,31,75,31,222,31,44,31,24,31,24,30,24,29,233,31,233,30,137,31,62,31,144,31,161,31,123,31,186,31,26,31,93,31,146,31,146,30,70,31,121,31,230,31,116,31,175,31,67,31,109,31,91,31,91,30,144,31,241,31,59,31,129,31,251,31,200,31,200,30,61,31,178,31,11,31,11,30,68,31,215,31,250,31,95,31,151,31,157,31,218,31,139,31,128,31,96,31,175,31,223,31,112,31,192,31,192,30,192,29,218,31,227,31,33,31,7,31,196,31,196,30,255,31,165,31,162,31,71,31,71,30,204,31,187,31,116,31,183,31,31,31,170,31,170,30,170,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
