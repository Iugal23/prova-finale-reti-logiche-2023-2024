-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 653;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (29,0,0,0,0,0,68,0,137,0,182,0,128,0,177,0,199,0,32,0,205,0,228,0,14,0,91,0,40,0,0,0,71,0,53,0,84,0,94,0,0,0,0,0,93,0,9,0,0,0,218,0,101,0,254,0,86,0,0,0,169,0,163,0,149,0,71,0,89,0,69,0,0,0,53,0,94,0,189,0,254,0,0,0,0,0,1,0,130,0,47,0,133,0,201,0,167,0,40,0,0,0,0,0,141,0,171,0,129,0,43,0,217,0,90,0,216,0,0,0,0,0,210,0,219,0,144,0,0,0,0,0,142,0,60,0,158,0,0,0,25,0,178,0,0,0,0,0,0,0,0,0,5,0,91,0,68,0,95,0,198,0,28,0,87,0,10,0,0,0,12,0,106,0,0,0,27,0,0,0,81,0,115,0,104,0,94,0,180,0,174,0,201,0,0,0,39,0,36,0,47,0,93,0,114,0,196,0,31,0,242,0,19,0,235,0,216,0,8,0,154,0,170,0,194,0,220,0,39,0,66,0,85,0,116,0,29,0,39,0,224,0,0,0,246,0,240,0,139,0,202,0,118,0,66,0,0,0,181,0,26,0,0,0,27,0,91,0,38,0,32,0,57,0,170,0,12,0,31,0,144,0,148,0,0,0,68,0,248,0,110,0,142,0,247,0,31,0,0,0,233,0,89,0,240,0,9,0,129,0,167,0,193,0,72,0,66,0,103,0,187,0,0,0,27,0,0,0,78,0,100,0,165,0,0,0,97,0,201,0,41,0,26,0,194,0,255,0,0,0,140,0,169,0,0,0,0,0,0,0,13,0,0,0,0,0,150,0,146,0,0,0,177,0,151,0,176,0,23,0,84,0,127,0,179,0,3,0,11,0,112,0,154,0,180,0,0,0,127,0,0,0,145,0,77,0,5,0,121,0,108,0,251,0,253,0,128,0,100,0,17,0,207,0,0,0,0,0,173,0,128,0,4,0,0,0,227,0,233,0,178,0,0,0,0,0,197,0,146,0,246,0,187,0,0,0,210,0,94,0,91,0,83,0,16,0,189,0,103,0,233,0,26,0,144,0,0,0,152,0,234,0,87,0,33,0,27,0,244,0,50,0,149,0,0,0,220,0,16,0,95,0,106,0,252,0,120,0,170,0,202,0,72,0,141,0,0,0,24,0,0,0,79,0,0,0,20,0,0,0,109,0,232,0,117,0,90,0,221,0,108,0,83,0,208,0,254,0,232,0,0,0,207,0,39,0,213,0,0,0,115,0,0,0,111,0,29,0,218,0,222,0,123,0,177,0,0,0,117,0,0,0,0,0,172,0,0,0,232,0,0,0,0,0,0,0,0,0,0,0,181,0,249,0,1,0,126,0,124,0,0,0,195,0,58,0,199,0,161,0,0,0,0,0,142,0,0,0,0,0,203,0,100,0,196,0,121,0,0,0,0,0,251,0,136,0,73,0,211,0,116,0,164,0,139,0,192,0,230,0,39,0,0,0,0,0,26,0,87,0,136,0,0,0,121,0,111,0,150,0,0,0,117,0,0,0,0,0,255,0,124,0,0,0,0,0,35,0,0,0,144,0,114,0,216,0,118,0,142,0,0,0,0,0,217,0,0,0,0,0,123,0,151,0,236,0,49,0,14,0,239,0,94,0,15,0,108,0,0,0,49,0,147,0,0,0,52,0,229,0,168,0,253,0,196,0,241,0,65,0,0,0,0,0,0,0,0,0,142,0,0,0,190,0,0,0,193,0,195,0,0,0,0,0,147,0,166,0,187,0,0,0,62,0,0,0,127,0,151,0,0,0,136,0,122,0,70,0,32,0,89,0,0,0,43,0,188,0,139,0,145,0,71,0,33,0,0,0,0,0,104,0,8,0,57,0,0,0,130,0,155,0,0,0,170,0,0,0,139,0,137,0,146,0,194,0,82,0,10,0,118,0,184,0,0,0,220,0,67,0,234,0,177,0,0,0,0,0,201,0,16,0,6,0,124,0,191,0,0,0,79,0,70,0,26,0,95,0,118,0,215,0,28,0,0,0,82,0,127,0,0,0,254,0,0,0,243,0,0,0,0,0,240,0,162,0,23,0,75,0,229,0,78,0,122,0,170,0,0,0,0,0,220,0,217,0,105,0,0,0,210,0,27,0,9,0,167,0,0,0,0,0,255,0,111,0,241,0,169,0,45,0,201,0,159,0,0,0,100,0,144,0,43,0,0,0,0,0,0,0,0,0,59,0,117,0,234,0,149,0,55,0,20,0,157,0,196,0,99,0,45,0,0,0,47,0,55,0,64,0,126,0,211,0,153,0,34,0,32,0,0,0,180,0,0,0,0,0,0,0,0,0,223,0,22,0,87,0,182,0,0,0,184,0,250,0,158,0,119,0,85,0,0,0,99,0,70,0,0,0,0,0,124,0,163,0,0,0,95,0,161,0,39,0,12,0,55,0,246,0,212,0,194,0,75,0,22,0,143,0,129,0,212,0,111,0,7,0,74,0,82,0,136,0,16,0,153,0,24,0,93,0,231,0,53,0,252,0,81,0,221,0,234,0,0,0,62,0,25,0,5,0,0,0,0,0,0,0,148,0,201,0,0,0,5,0,54,0,0,0,149,0,78,0,240,0,255,0,209,0,231,0,117,0,72,0,242,0,158,0,153,0,9,0,180,0,0,0,0,0,50,0,0,0,0,0,37,0,228,0,200,0,0,0,133,0,33,0,0,0,6,0,103,0,0,0,36,0,0,0,9,0,36,0,195,0,11,0,149,0,0,0,58,0,46,0,145,0,0,0,0,0,223,0,148,0,226,0,0,0,235,0,87,0,0,0,143,0,191,0,174,0,0,0,40,0,14,0,0,0,134,0,224,0,103,0,231,0,241,0,49,0,139,0,124,0,202,0,58,0,98,0,248,0,7,0,158,0,35,0,0,0,146,0,223,0);
signal scenario_full  : scenario_type := (29,31,29,30,29,29,68,31,137,31,182,31,128,31,177,31,199,31,32,31,205,31,228,31,14,31,91,31,40,31,40,30,71,31,53,31,84,31,94,31,94,30,94,29,93,31,9,31,9,30,218,31,101,31,254,31,86,31,86,30,169,31,163,31,149,31,71,31,89,31,69,31,69,30,53,31,94,31,189,31,254,31,254,30,254,29,1,31,130,31,47,31,133,31,201,31,167,31,40,31,40,30,40,29,141,31,171,31,129,31,43,31,217,31,90,31,216,31,216,30,216,29,210,31,219,31,144,31,144,30,144,29,142,31,60,31,158,31,158,30,25,31,178,31,178,30,178,29,178,28,178,27,5,31,91,31,68,31,95,31,198,31,28,31,87,31,10,31,10,30,12,31,106,31,106,30,27,31,27,30,81,31,115,31,104,31,94,31,180,31,174,31,201,31,201,30,39,31,36,31,47,31,93,31,114,31,196,31,31,31,242,31,19,31,235,31,216,31,8,31,154,31,170,31,194,31,220,31,39,31,66,31,85,31,116,31,29,31,39,31,224,31,224,30,246,31,240,31,139,31,202,31,118,31,66,31,66,30,181,31,26,31,26,30,27,31,91,31,38,31,32,31,57,31,170,31,12,31,31,31,144,31,148,31,148,30,68,31,248,31,110,31,142,31,247,31,31,31,31,30,233,31,89,31,240,31,9,31,129,31,167,31,193,31,72,31,66,31,103,31,187,31,187,30,27,31,27,30,78,31,100,31,165,31,165,30,97,31,201,31,41,31,26,31,194,31,255,31,255,30,140,31,169,31,169,30,169,29,169,28,13,31,13,30,13,29,150,31,146,31,146,30,177,31,151,31,176,31,23,31,84,31,127,31,179,31,3,31,11,31,112,31,154,31,180,31,180,30,127,31,127,30,145,31,77,31,5,31,121,31,108,31,251,31,253,31,128,31,100,31,17,31,207,31,207,30,207,29,173,31,128,31,4,31,4,30,227,31,233,31,178,31,178,30,178,29,197,31,146,31,246,31,187,31,187,30,210,31,94,31,91,31,83,31,16,31,189,31,103,31,233,31,26,31,144,31,144,30,152,31,234,31,87,31,33,31,27,31,244,31,50,31,149,31,149,30,220,31,16,31,95,31,106,31,252,31,120,31,170,31,202,31,72,31,141,31,141,30,24,31,24,30,79,31,79,30,20,31,20,30,109,31,232,31,117,31,90,31,221,31,108,31,83,31,208,31,254,31,232,31,232,30,207,31,39,31,213,31,213,30,115,31,115,30,111,31,29,31,218,31,222,31,123,31,177,31,177,30,117,31,117,30,117,29,172,31,172,30,232,31,232,30,232,29,232,28,232,27,232,26,181,31,249,31,1,31,126,31,124,31,124,30,195,31,58,31,199,31,161,31,161,30,161,29,142,31,142,30,142,29,203,31,100,31,196,31,121,31,121,30,121,29,251,31,136,31,73,31,211,31,116,31,164,31,139,31,192,31,230,31,39,31,39,30,39,29,26,31,87,31,136,31,136,30,121,31,111,31,150,31,150,30,117,31,117,30,117,29,255,31,124,31,124,30,124,29,35,31,35,30,144,31,114,31,216,31,118,31,142,31,142,30,142,29,217,31,217,30,217,29,123,31,151,31,236,31,49,31,14,31,239,31,94,31,15,31,108,31,108,30,49,31,147,31,147,30,52,31,229,31,168,31,253,31,196,31,241,31,65,31,65,30,65,29,65,28,65,27,142,31,142,30,190,31,190,30,193,31,195,31,195,30,195,29,147,31,166,31,187,31,187,30,62,31,62,30,127,31,151,31,151,30,136,31,122,31,70,31,32,31,89,31,89,30,43,31,188,31,139,31,145,31,71,31,33,31,33,30,33,29,104,31,8,31,57,31,57,30,130,31,155,31,155,30,170,31,170,30,139,31,137,31,146,31,194,31,82,31,10,31,118,31,184,31,184,30,220,31,67,31,234,31,177,31,177,30,177,29,201,31,16,31,6,31,124,31,191,31,191,30,79,31,70,31,26,31,95,31,118,31,215,31,28,31,28,30,82,31,127,31,127,30,254,31,254,30,243,31,243,30,243,29,240,31,162,31,23,31,75,31,229,31,78,31,122,31,170,31,170,30,170,29,220,31,217,31,105,31,105,30,210,31,27,31,9,31,167,31,167,30,167,29,255,31,111,31,241,31,169,31,45,31,201,31,159,31,159,30,100,31,144,31,43,31,43,30,43,29,43,28,43,27,59,31,117,31,234,31,149,31,55,31,20,31,157,31,196,31,99,31,45,31,45,30,47,31,55,31,64,31,126,31,211,31,153,31,34,31,32,31,32,30,180,31,180,30,180,29,180,28,180,27,223,31,22,31,87,31,182,31,182,30,184,31,250,31,158,31,119,31,85,31,85,30,99,31,70,31,70,30,70,29,124,31,163,31,163,30,95,31,161,31,39,31,12,31,55,31,246,31,212,31,194,31,75,31,22,31,143,31,129,31,212,31,111,31,7,31,74,31,82,31,136,31,16,31,153,31,24,31,93,31,231,31,53,31,252,31,81,31,221,31,234,31,234,30,62,31,25,31,5,31,5,30,5,29,5,28,148,31,201,31,201,30,5,31,54,31,54,30,149,31,78,31,240,31,255,31,209,31,231,31,117,31,72,31,242,31,158,31,153,31,9,31,180,31,180,30,180,29,50,31,50,30,50,29,37,31,228,31,200,31,200,30,133,31,33,31,33,30,6,31,103,31,103,30,36,31,36,30,9,31,36,31,195,31,11,31,149,31,149,30,58,31,46,31,145,31,145,30,145,29,223,31,148,31,226,31,226,30,235,31,87,31,87,30,143,31,191,31,174,31,174,30,40,31,14,31,14,30,134,31,224,31,103,31,231,31,241,31,49,31,139,31,124,31,202,31,58,31,98,31,248,31,7,31,158,31,35,31,35,30,146,31,223,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
