-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_12 is
end project_tb_12;

architecture project_tb_arch_12 of project_tb_12 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 172;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (245,0,72,0,42,0,45,0,41,0,228,0,100,0,214,0,0,0,217,0,176,0,199,0,73,0,50,0,246,0,194,0,78,0,152,0,209,0,86,0,5,0,0,0,187,0,249,0,0,0,168,0,58,0,53,0,62,0,131,0,0,0,0,0,251,0,46,0,0,0,133,0,174,0,148,0,180,0,0,0,129,0,68,0,152,0,159,0,249,0,15,0,175,0,58,0,152,0,0,0,247,0,20,0,170,0,0,0,57,0,32,0,224,0,0,0,39,0,0,0,0,0,47,0,111,0,0,0,0,0,0,0,140,0,0,0,46,0,0,0,150,0,0,0,8,0,155,0,217,0,155,0,53,0,156,0,0,0,209,0,36,0,110,0,168,0,0,0,201,0,23,0,208,0,0,0,170,0,0,0,160,0,69,0,75,0,0,0,0,0,80,0,65,0,94,0,115,0,253,0,178,0,200,0,0,0,169,0,0,0,131,0,32,0,120,0,106,0,79,0,169,0,88,0,4,0,0,0,29,0,118,0,197,0,0,0,254,0,0,0,63,0,182,0,252,0,49,0,117,0,0,0,137,0,0,0,0,0,96,0,0,0,142,0,168,0,225,0,161,0,96,0,28,0,140,0,231,0,87,0,183,0,204,0,52,0,11,0,199,0,0,0,0,0,226,0,98,0,187,0,145,0,217,0,214,0,135,0,226,0,128,0,106,0,0,0,177,0,0,0,0,0,227,0,34,0,135,0,78,0,231,0,197,0,151,0,0,0,0,0,212,0,66,0);
signal scenario_full  : scenario_type := (245,31,72,31,42,31,45,31,41,31,228,31,100,31,214,31,214,30,217,31,176,31,199,31,73,31,50,31,246,31,194,31,78,31,152,31,209,31,86,31,5,31,5,30,187,31,249,31,249,30,168,31,58,31,53,31,62,31,131,31,131,30,131,29,251,31,46,31,46,30,133,31,174,31,148,31,180,31,180,30,129,31,68,31,152,31,159,31,249,31,15,31,175,31,58,31,152,31,152,30,247,31,20,31,170,31,170,30,57,31,32,31,224,31,224,30,39,31,39,30,39,29,47,31,111,31,111,30,111,29,111,28,140,31,140,30,46,31,46,30,150,31,150,30,8,31,155,31,217,31,155,31,53,31,156,31,156,30,209,31,36,31,110,31,168,31,168,30,201,31,23,31,208,31,208,30,170,31,170,30,160,31,69,31,75,31,75,30,75,29,80,31,65,31,94,31,115,31,253,31,178,31,200,31,200,30,169,31,169,30,131,31,32,31,120,31,106,31,79,31,169,31,88,31,4,31,4,30,29,31,118,31,197,31,197,30,254,31,254,30,63,31,182,31,252,31,49,31,117,31,117,30,137,31,137,30,137,29,96,31,96,30,142,31,168,31,225,31,161,31,96,31,28,31,140,31,231,31,87,31,183,31,204,31,52,31,11,31,199,31,199,30,199,29,226,31,98,31,187,31,145,31,217,31,214,31,135,31,226,31,128,31,106,31,106,30,177,31,177,30,177,29,227,31,34,31,135,31,78,31,231,31,197,31,151,31,151,30,151,29,212,31,66,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
