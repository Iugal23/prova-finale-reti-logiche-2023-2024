-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 844;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (127,0,248,0,221,0,28,0,185,0,7,0,99,0,127,0,27,0,0,0,244,0,0,0,31,0,143,0,181,0,0,0,0,0,0,0,235,0,0,0,4,0,0,0,56,0,155,0,120,0,49,0,0,0,0,0,62,0,199,0,220,0,48,0,59,0,0,0,113,0,0,0,71,0,20,0,159,0,42,0,45,0,146,0,74,0,127,0,92,0,0,0,121,0,212,0,162,0,1,0,181,0,0,0,107,0,72,0,82,0,80,0,127,0,208,0,49,0,40,0,130,0,138,0,223,0,0,0,0,0,253,0,3,0,0,0,0,0,0,0,118,0,100,0,0,0,208,0,236,0,39,0,245,0,54,0,198,0,217,0,78,0,128,0,104,0,89,0,0,0,53,0,0,0,109,0,0,0,0,0,207,0,172,0,210,0,0,0,148,0,148,0,220,0,32,0,0,0,45,0,0,0,89,0,15,0,172,0,115,0,0,0,104,0,202,0,206,0,129,0,26,0,180,0,95,0,56,0,228,0,240,0,29,0,137,0,198,0,22,0,168,0,235,0,0,0,219,0,198,0,43,0,65,0,199,0,226,0,14,0,0,0,171,0,242,0,229,0,220,0,30,0,0,0,79,0,0,0,65,0,57,0,119,0,211,0,133,0,222,0,181,0,126,0,53,0,0,0,72,0,169,0,0,0,147,0,92,0,200,0,166,0,217,0,0,0,7,0,11,0,37,0,98,0,191,0,191,0,129,0,86,0,0,0,108,0,0,0,220,0,193,0,124,0,78,0,162,0,69,0,190,0,150,0,15,0,230,0,0,0,0,0,0,0,112,0,0,0,171,0,82,0,181,0,58,0,0,0,216,0,0,0,19,0,240,0,219,0,105,0,33,0,0,0,98,0,248,0,211,0,149,0,0,0,156,0,26,0,86,0,151,0,214,0,107,0,93,0,0,0,120,0,123,0,224,0,90,0,82,0,0,0,45,0,192,0,0,0,41,0,1,0,187,0,154,0,101,0,0,0,0,0,122,0,195,0,8,0,8,0,38,0,223,0,0,0,199,0,227,0,164,0,166,0,40,0,0,0,0,0,226,0,139,0,226,0,189,0,0,0,0,0,137,0,0,0,157,0,167,0,15,0,201,0,61,0,0,0,186,0,238,0,129,0,172,0,42,0,104,0,170,0,36,0,96,0,165,0,165,0,68,0,112,0,69,0,0,0,50,0,166,0,1,0,76,0,88,0,111,0,38,0,117,0,194,0,85,0,32,0,209,0,146,0,148,0,199,0,53,0,72,0,173,0,8,0,195,0,191,0,106,0,0,0,136,0,0,0,189,0,27,0,107,0,141,0,0,0,46,0,207,0,255,0,222,0,0,0,235,0,235,0,29,0,241,0,145,0,11,0,188,0,0,0,240,0,82,0,191,0,68,0,46,0,121,0,55,0,31,0,251,0,5,0,230,0,103,0,42,0,110,0,137,0,93,0,0,0,192,0,189,0,157,0,177,0,11,0,119,0,36,0,1,0,71,0,0,0,0,0,120,0,233,0,135,0,0,0,0,0,0,0,248,0,204,0,4,0,0,0,232,0,149,0,189,0,240,0,102,0,227,0,62,0,146,0,226,0,242,0,2,0,52,0,35,0,131,0,157,0,251,0,106,0,0,0,19,0,0,0,219,0,0,0,90,0,99,0,110,0,173,0,72,0,215,0,130,0,236,0,90,0,205,0,111,0,131,0,0,0,192,0,118,0,90,0,225,0,253,0,101,0,216,0,126,0,160,0,0,0,51,0,119,0,115,0,102,0,62,0,0,0,226,0,31,0,179,0,144,0,229,0,116,0,22,0,11,0,37,0,0,0,200,0,200,0,125,0,12,0,160,0,0,0,91,0,230,0,101,0,11,0,86,0,145,0,211,0,246,0,0,0,80,0,73,0,83,0,210,0,0,0,131,0,0,0,236,0,238,0,0,0,253,0,0,0,157,0,252,0,238,0,134,0,9,0,0,0,39,0,0,0,100,0,0,0,88,0,0,0,73,0,56,0,224,0,138,0,232,0,133,0,94,0,0,0,10,0,254,0,0,0,136,0,100,0,253,0,0,0,217,0,0,0,200,0,11,0,61,0,237,0,195,0,106,0,8,0,245,0,0,0,163,0,78,0,186,0,83,0,97,0,136,0,82,0,205,0,131,0,0,0,46,0,73,0,0,0,123,0,55,0,104,0,84,0,213,0,201,0,1,0,216,0,0,0,108,0,0,0,0,0,38,0,186,0,123,0,47,0,7,0,0,0,0,0,79,0,0,0,254,0,0,0,0,0,197,0,94,0,27,0,0,0,149,0,233,0,0,0,172,0,207,0,190,0,60,0,0,0,0,0,51,0,0,0,57,0,80,0,157,0,0,0,36,0,167,0,40,0,0,0,204,0,46,0,129,0,0,0,199,0,150,0,229,0,226,0,0,0,71,0,0,0,236,0,90,0,0,0,23,0,0,0,0,0,158,0,42,0,124,0,116,0,211,0,0,0,140,0,59,0,0,0,132,0,141,0,0,0,0,0,6,0,180,0,95,0,133,0,0,0,255,0,114,0,0,0,0,0,236,0,146,0,121,0,121,0,223,0,137,0,67,0,72,0,21,0,16,0,177,0,124,0,0,0,0,0,181,0,145,0,148,0,101,0,0,0,107,0,184,0,25,0,0,0,0,0,66,0,0,0,229,0,177,0,207,0,151,0,225,0,0,0,0,0,57,0,0,0,6,0,183,0,174,0,177,0,153,0,197,0,139,0,11,0,226,0,0,0,95,0,89,0,223,0,37,0,186,0,177,0,59,0,74,0,3,0,126,0,242,0,0,0,0,0,0,0,120,0,16,0,243,0,175,0,95,0,138,0,227,0,103,0,140,0,141,0,46,0,92,0,36,0,0,0,221,0,67,0,34,0,154,0,244,0,0,0,90,0,4,0,202,0,185,0,201,0,231,0,70,0,177,0,0,0,44,0,0,0,117,0,0,0,73,0,206,0,0,0,141,0,179,0,232,0,209,0,0,0,188,0,108,0,67,0,168,0,0,0,69,0,73,0,170,0,186,0,7,0,157,0,169,0,37,0,71,0,6,0,97,0,223,0,135,0,90,0,174,0,0,0,0,0,237,0,41,0,134,0,64,0,214,0,4,0,26,0,0,0,171,0,204,0,182,0,189,0,136,0,176,0,0,0,75,0,135,0,78,0,116,0,45,0,219,0,253,0,66,0,39,0,50,0,0,0,13,0,170,0,49,0,117,0,166,0,215,0,248,0,59,0,0,0,231,0,0,0,225,0,138,0,239,0,60,0,0,0,250,0,254,0,22,0,217,0,162,0,98,0,123,0,172,0,112,0,29,0,110,0,201,0,98,0,171,0,0,0,177,0,117,0,231,0,92,0,241,0,119,0,214,0,0,0,232,0,158,0,0,0,0,0,124,0,48,0,163,0,173,0,201,0,109,0,104,0,175,0,230,0,12,0,0,0,178,0,240,0,114,0,229,0,0,0,184,0,237,0,26,0,0,0,65,0,60,0,166,0,208,0,200,0,238,0,78,0,240,0,107,0,1,0,0,0,174,0,0,0,143,0,47,0,81,0,253,0,233,0,62,0,83,0,103,0,0,0,61,0,0,0,174,0,60,0,0,0,203,0,201,0,73,0,213,0,174,0,186,0,30,0,145,0,105,0,160,0,128,0,212,0,106,0,114,0,108,0,0,0,36,0,156,0,243,0,96,0,0,0,245,0,100,0,69,0,0,0,237,0,235,0,204,0,0,0,121,0,51,0);
signal scenario_full  : scenario_type := (127,31,248,31,221,31,28,31,185,31,7,31,99,31,127,31,27,31,27,30,244,31,244,30,31,31,143,31,181,31,181,30,181,29,181,28,235,31,235,30,4,31,4,30,56,31,155,31,120,31,49,31,49,30,49,29,62,31,199,31,220,31,48,31,59,31,59,30,113,31,113,30,71,31,20,31,159,31,42,31,45,31,146,31,74,31,127,31,92,31,92,30,121,31,212,31,162,31,1,31,181,31,181,30,107,31,72,31,82,31,80,31,127,31,208,31,49,31,40,31,130,31,138,31,223,31,223,30,223,29,253,31,3,31,3,30,3,29,3,28,118,31,100,31,100,30,208,31,236,31,39,31,245,31,54,31,198,31,217,31,78,31,128,31,104,31,89,31,89,30,53,31,53,30,109,31,109,30,109,29,207,31,172,31,210,31,210,30,148,31,148,31,220,31,32,31,32,30,45,31,45,30,89,31,15,31,172,31,115,31,115,30,104,31,202,31,206,31,129,31,26,31,180,31,95,31,56,31,228,31,240,31,29,31,137,31,198,31,22,31,168,31,235,31,235,30,219,31,198,31,43,31,65,31,199,31,226,31,14,31,14,30,171,31,242,31,229,31,220,31,30,31,30,30,79,31,79,30,65,31,57,31,119,31,211,31,133,31,222,31,181,31,126,31,53,31,53,30,72,31,169,31,169,30,147,31,92,31,200,31,166,31,217,31,217,30,7,31,11,31,37,31,98,31,191,31,191,31,129,31,86,31,86,30,108,31,108,30,220,31,193,31,124,31,78,31,162,31,69,31,190,31,150,31,15,31,230,31,230,30,230,29,230,28,112,31,112,30,171,31,82,31,181,31,58,31,58,30,216,31,216,30,19,31,240,31,219,31,105,31,33,31,33,30,98,31,248,31,211,31,149,31,149,30,156,31,26,31,86,31,151,31,214,31,107,31,93,31,93,30,120,31,123,31,224,31,90,31,82,31,82,30,45,31,192,31,192,30,41,31,1,31,187,31,154,31,101,31,101,30,101,29,122,31,195,31,8,31,8,31,38,31,223,31,223,30,199,31,227,31,164,31,166,31,40,31,40,30,40,29,226,31,139,31,226,31,189,31,189,30,189,29,137,31,137,30,157,31,167,31,15,31,201,31,61,31,61,30,186,31,238,31,129,31,172,31,42,31,104,31,170,31,36,31,96,31,165,31,165,31,68,31,112,31,69,31,69,30,50,31,166,31,1,31,76,31,88,31,111,31,38,31,117,31,194,31,85,31,32,31,209,31,146,31,148,31,199,31,53,31,72,31,173,31,8,31,195,31,191,31,106,31,106,30,136,31,136,30,189,31,27,31,107,31,141,31,141,30,46,31,207,31,255,31,222,31,222,30,235,31,235,31,29,31,241,31,145,31,11,31,188,31,188,30,240,31,82,31,191,31,68,31,46,31,121,31,55,31,31,31,251,31,5,31,230,31,103,31,42,31,110,31,137,31,93,31,93,30,192,31,189,31,157,31,177,31,11,31,119,31,36,31,1,31,71,31,71,30,71,29,120,31,233,31,135,31,135,30,135,29,135,28,248,31,204,31,4,31,4,30,232,31,149,31,189,31,240,31,102,31,227,31,62,31,146,31,226,31,242,31,2,31,52,31,35,31,131,31,157,31,251,31,106,31,106,30,19,31,19,30,219,31,219,30,90,31,99,31,110,31,173,31,72,31,215,31,130,31,236,31,90,31,205,31,111,31,131,31,131,30,192,31,118,31,90,31,225,31,253,31,101,31,216,31,126,31,160,31,160,30,51,31,119,31,115,31,102,31,62,31,62,30,226,31,31,31,179,31,144,31,229,31,116,31,22,31,11,31,37,31,37,30,200,31,200,31,125,31,12,31,160,31,160,30,91,31,230,31,101,31,11,31,86,31,145,31,211,31,246,31,246,30,80,31,73,31,83,31,210,31,210,30,131,31,131,30,236,31,238,31,238,30,253,31,253,30,157,31,252,31,238,31,134,31,9,31,9,30,39,31,39,30,100,31,100,30,88,31,88,30,73,31,56,31,224,31,138,31,232,31,133,31,94,31,94,30,10,31,254,31,254,30,136,31,100,31,253,31,253,30,217,31,217,30,200,31,11,31,61,31,237,31,195,31,106,31,8,31,245,31,245,30,163,31,78,31,186,31,83,31,97,31,136,31,82,31,205,31,131,31,131,30,46,31,73,31,73,30,123,31,55,31,104,31,84,31,213,31,201,31,1,31,216,31,216,30,108,31,108,30,108,29,38,31,186,31,123,31,47,31,7,31,7,30,7,29,79,31,79,30,254,31,254,30,254,29,197,31,94,31,27,31,27,30,149,31,233,31,233,30,172,31,207,31,190,31,60,31,60,30,60,29,51,31,51,30,57,31,80,31,157,31,157,30,36,31,167,31,40,31,40,30,204,31,46,31,129,31,129,30,199,31,150,31,229,31,226,31,226,30,71,31,71,30,236,31,90,31,90,30,23,31,23,30,23,29,158,31,42,31,124,31,116,31,211,31,211,30,140,31,59,31,59,30,132,31,141,31,141,30,141,29,6,31,180,31,95,31,133,31,133,30,255,31,114,31,114,30,114,29,236,31,146,31,121,31,121,31,223,31,137,31,67,31,72,31,21,31,16,31,177,31,124,31,124,30,124,29,181,31,145,31,148,31,101,31,101,30,107,31,184,31,25,31,25,30,25,29,66,31,66,30,229,31,177,31,207,31,151,31,225,31,225,30,225,29,57,31,57,30,6,31,183,31,174,31,177,31,153,31,197,31,139,31,11,31,226,31,226,30,95,31,89,31,223,31,37,31,186,31,177,31,59,31,74,31,3,31,126,31,242,31,242,30,242,29,242,28,120,31,16,31,243,31,175,31,95,31,138,31,227,31,103,31,140,31,141,31,46,31,92,31,36,31,36,30,221,31,67,31,34,31,154,31,244,31,244,30,90,31,4,31,202,31,185,31,201,31,231,31,70,31,177,31,177,30,44,31,44,30,117,31,117,30,73,31,206,31,206,30,141,31,179,31,232,31,209,31,209,30,188,31,108,31,67,31,168,31,168,30,69,31,73,31,170,31,186,31,7,31,157,31,169,31,37,31,71,31,6,31,97,31,223,31,135,31,90,31,174,31,174,30,174,29,237,31,41,31,134,31,64,31,214,31,4,31,26,31,26,30,171,31,204,31,182,31,189,31,136,31,176,31,176,30,75,31,135,31,78,31,116,31,45,31,219,31,253,31,66,31,39,31,50,31,50,30,13,31,170,31,49,31,117,31,166,31,215,31,248,31,59,31,59,30,231,31,231,30,225,31,138,31,239,31,60,31,60,30,250,31,254,31,22,31,217,31,162,31,98,31,123,31,172,31,112,31,29,31,110,31,201,31,98,31,171,31,171,30,177,31,117,31,231,31,92,31,241,31,119,31,214,31,214,30,232,31,158,31,158,30,158,29,124,31,48,31,163,31,173,31,201,31,109,31,104,31,175,31,230,31,12,31,12,30,178,31,240,31,114,31,229,31,229,30,184,31,237,31,26,31,26,30,65,31,60,31,166,31,208,31,200,31,238,31,78,31,240,31,107,31,1,31,1,30,174,31,174,30,143,31,47,31,81,31,253,31,233,31,62,31,83,31,103,31,103,30,61,31,61,30,174,31,60,31,60,30,203,31,201,31,73,31,213,31,174,31,186,31,30,31,145,31,105,31,160,31,128,31,212,31,106,31,114,31,108,31,108,30,36,31,156,31,243,31,96,31,96,30,245,31,100,31,69,31,69,30,237,31,235,31,204,31,204,30,121,31,51,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
