-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_47 is
end project_tb_47;

architecture project_tb_arch_47 of project_tb_47 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 425;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (2,0,123,0,6,0,23,0,64,0,211,0,194,0,181,0,74,0,92,0,104,0,158,0,88,0,190,0,95,0,252,0,0,0,156,0,155,0,238,0,0,0,237,0,14,0,54,0,0,0,43,0,194,0,137,0,117,0,0,0,189,0,15,0,217,0,0,0,53,0,0,0,0,0,30,0,34,0,159,0,222,0,145,0,0,0,98,0,207,0,148,0,114,0,14,0,125,0,209,0,254,0,229,0,217,0,0,0,80,0,254,0,0,0,99,0,142,0,93,0,228,0,50,0,143,0,48,0,3,0,226,0,185,0,161,0,246,0,234,0,0,0,184,0,92,0,107,0,159,0,214,0,45,0,111,0,0,0,0,0,197,0,233,0,247,0,4,0,0,0,14,0,246,0,0,0,153,0,148,0,0,0,198,0,162,0,27,0,147,0,42,0,140,0,65,0,36,0,101,0,83,0,193,0,125,0,31,0,93,0,212,0,254,0,250,0,246,0,72,0,35,0,178,0,64,0,0,0,73,0,161,0,166,0,86,0,203,0,192,0,78,0,6,0,186,0,0,0,84,0,87,0,0,0,101,0,0,0,26,0,0,0,111,0,49,0,68,0,0,0,113,0,162,0,196,0,21,0,247,0,1,0,0,0,120,0,153,0,246,0,41,0,0,0,226,0,99,0,234,0,206,0,149,0,193,0,142,0,234,0,92,0,251,0,65,0,223,0,80,0,231,0,0,0,180,0,145,0,27,0,14,0,17,0,0,0,107,0,89,0,86,0,17,0,168,0,34,0,214,0,35,0,236,0,76,0,10,0,50,0,0,0,119,0,139,0,136,0,91,0,14,0,15,0,30,0,148,0,50,0,0,0,0,0,207,0,1,0,47,0,68,0,82,0,105,0,154,0,0,0,88,0,93,0,200,0,191,0,239,0,120,0,0,0,114,0,181,0,102,0,15,0,16,0,0,0,0,0,34,0,0,0,201,0,214,0,220,0,172,0,39,0,197,0,0,0,162,0,173,0,148,0,153,0,43,0,21,0,61,0,73,0,38,0,0,0,166,0,141,0,218,0,126,0,157,0,63,0,61,0,197,0,32,0,96,0,247,0,0,0,115,0,26,0,220,0,69,0,0,0,0,0,157,0,0,0,157,0,70,0,0,0,40,0,22,0,0,0,232,0,197,0,28,0,0,0,79,0,130,0,23,0,212,0,94,0,212,0,131,0,90,0,192,0,93,0,116,0,98,0,101,0,181,0,176,0,23,0,16,0,10,0,242,0,173,0,22,0,46,0,0,0,180,0,227,0,0,0,47,0,0,0,244,0,55,0,97,0,10,0,115,0,153,0,213,0,90,0,0,0,78,0,24,0,101,0,112,0,81,0,252,0,255,0,120,0,185,0,63,0,196,0,104,0,0,0,0,0,123,0,0,0,157,0,60,0,21,0,45,0,0,0,180,0,20,0,142,0,33,0,111,0,162,0,0,0,162,0,0,0,218,0,168,0,85,0,0,0,241,0,70,0,215,0,249,0,0,0,0,0,0,0,182,0,0,0,0,0,177,0,0,0,236,0,0,0,96,0,0,0,204,0,99,0,170,0,102,0,34,0,0,0,137,0,174,0,233,0,111,0,38,0,0,0,240,0,0,0,11,0,64,0,45,0,79,0,7,0,222,0,0,0,18,0,98,0,183,0,178,0,12,0,255,0,72,0,0,0,0,0,0,0,152,0,180,0,0,0,137,0,36,0,163,0,0,0,0,0,3,0,145,0,0,0,29,0,188,0,20,0,126,0,23,0,22,0,80,0,181,0,102,0,63,0,243,0,62,0,0,0,57,0,32,0,0,0,246,0,71,0,0,0,0,0,0,0,32,0,130,0,166,0,0,0,228,0,0,0,90,0,130,0,2,0,202,0,204,0,174,0);
signal scenario_full  : scenario_type := (2,31,123,31,6,31,23,31,64,31,211,31,194,31,181,31,74,31,92,31,104,31,158,31,88,31,190,31,95,31,252,31,252,30,156,31,155,31,238,31,238,30,237,31,14,31,54,31,54,30,43,31,194,31,137,31,117,31,117,30,189,31,15,31,217,31,217,30,53,31,53,30,53,29,30,31,34,31,159,31,222,31,145,31,145,30,98,31,207,31,148,31,114,31,14,31,125,31,209,31,254,31,229,31,217,31,217,30,80,31,254,31,254,30,99,31,142,31,93,31,228,31,50,31,143,31,48,31,3,31,226,31,185,31,161,31,246,31,234,31,234,30,184,31,92,31,107,31,159,31,214,31,45,31,111,31,111,30,111,29,197,31,233,31,247,31,4,31,4,30,14,31,246,31,246,30,153,31,148,31,148,30,198,31,162,31,27,31,147,31,42,31,140,31,65,31,36,31,101,31,83,31,193,31,125,31,31,31,93,31,212,31,254,31,250,31,246,31,72,31,35,31,178,31,64,31,64,30,73,31,161,31,166,31,86,31,203,31,192,31,78,31,6,31,186,31,186,30,84,31,87,31,87,30,101,31,101,30,26,31,26,30,111,31,49,31,68,31,68,30,113,31,162,31,196,31,21,31,247,31,1,31,1,30,120,31,153,31,246,31,41,31,41,30,226,31,99,31,234,31,206,31,149,31,193,31,142,31,234,31,92,31,251,31,65,31,223,31,80,31,231,31,231,30,180,31,145,31,27,31,14,31,17,31,17,30,107,31,89,31,86,31,17,31,168,31,34,31,214,31,35,31,236,31,76,31,10,31,50,31,50,30,119,31,139,31,136,31,91,31,14,31,15,31,30,31,148,31,50,31,50,30,50,29,207,31,1,31,47,31,68,31,82,31,105,31,154,31,154,30,88,31,93,31,200,31,191,31,239,31,120,31,120,30,114,31,181,31,102,31,15,31,16,31,16,30,16,29,34,31,34,30,201,31,214,31,220,31,172,31,39,31,197,31,197,30,162,31,173,31,148,31,153,31,43,31,21,31,61,31,73,31,38,31,38,30,166,31,141,31,218,31,126,31,157,31,63,31,61,31,197,31,32,31,96,31,247,31,247,30,115,31,26,31,220,31,69,31,69,30,69,29,157,31,157,30,157,31,70,31,70,30,40,31,22,31,22,30,232,31,197,31,28,31,28,30,79,31,130,31,23,31,212,31,94,31,212,31,131,31,90,31,192,31,93,31,116,31,98,31,101,31,181,31,176,31,23,31,16,31,10,31,242,31,173,31,22,31,46,31,46,30,180,31,227,31,227,30,47,31,47,30,244,31,55,31,97,31,10,31,115,31,153,31,213,31,90,31,90,30,78,31,24,31,101,31,112,31,81,31,252,31,255,31,120,31,185,31,63,31,196,31,104,31,104,30,104,29,123,31,123,30,157,31,60,31,21,31,45,31,45,30,180,31,20,31,142,31,33,31,111,31,162,31,162,30,162,31,162,30,218,31,168,31,85,31,85,30,241,31,70,31,215,31,249,31,249,30,249,29,249,28,182,31,182,30,182,29,177,31,177,30,236,31,236,30,96,31,96,30,204,31,99,31,170,31,102,31,34,31,34,30,137,31,174,31,233,31,111,31,38,31,38,30,240,31,240,30,11,31,64,31,45,31,79,31,7,31,222,31,222,30,18,31,98,31,183,31,178,31,12,31,255,31,72,31,72,30,72,29,72,28,152,31,180,31,180,30,137,31,36,31,163,31,163,30,163,29,3,31,145,31,145,30,29,31,188,31,20,31,126,31,23,31,22,31,80,31,181,31,102,31,63,31,243,31,62,31,62,30,57,31,32,31,32,30,246,31,71,31,71,30,71,29,71,28,32,31,130,31,166,31,166,30,228,31,228,30,90,31,130,31,2,31,202,31,204,31,174,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
