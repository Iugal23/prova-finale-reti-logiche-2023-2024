-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 976;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (37,0,41,0,0,0,0,0,192,0,229,0,182,0,91,0,17,0,149,0,40,0,38,0,0,0,215,0,69,0,43,0,56,0,0,0,244,0,25,0,84,0,159,0,168,0,99,0,157,0,222,0,190,0,0,0,37,0,104,0,214,0,143,0,216,0,172,0,151,0,11,0,0,0,194,0,0,0,231,0,213,0,212,0,234,0,188,0,204,0,0,0,231,0,162,0,123,0,108,0,114,0,16,0,165,0,3,0,0,0,128,0,217,0,0,0,253,0,18,0,196,0,11,0,0,0,110,0,190,0,16,0,207,0,0,0,84,0,38,0,0,0,5,0,106,0,0,0,220,0,10,0,168,0,35,0,230,0,149,0,100,0,0,0,0,0,0,0,188,0,116,0,208,0,18,0,87,0,0,0,234,0,107,0,131,0,157,0,0,0,245,0,0,0,0,0,62,0,164,0,171,0,179,0,207,0,234,0,119,0,198,0,0,0,208,0,115,0,73,0,91,0,156,0,0,0,209,0,126,0,5,0,52,0,80,0,21,0,128,0,0,0,196,0,102,0,0,0,63,0,54,0,0,0,211,0,0,0,91,0,136,0,0,0,0,0,0,0,180,0,208,0,230,0,134,0,100,0,0,0,0,0,99,0,79,0,65,0,203,0,0,0,52,0,14,0,115,0,215,0,0,0,255,0,190,0,145,0,95,0,224,0,0,0,126,0,0,0,54,0,87,0,0,0,82,0,0,0,0,0,27,0,170,0,105,0,79,0,25,0,0,0,0,0,0,0,186,0,141,0,0,0,81,0,0,0,114,0,0,0,233,0,196,0,174,0,31,0,246,0,159,0,81,0,96,0,176,0,237,0,245,0,35,0,198,0,60,0,16,0,0,0,155,0,144,0,0,0,24,0,11,0,199,0,157,0,157,0,0,0,6,0,182,0,154,0,0,0,89,0,21,0,122,0,163,0,173,0,169,0,10,0,32,0,103,0,0,0,210,0,232,0,32,0,148,0,212,0,247,0,135,0,4,0,0,0,0,0,149,0,254,0,0,0,123,0,170,0,21,0,82,0,168,0,0,0,231,0,203,0,8,0,0,0,242,0,226,0,0,0,2,0,40,0,187,0,112,0,52,0,67,0,72,0,0,0,0,0,229,0,149,0,0,0,85,0,141,0,103,0,114,0,44,0,126,0,135,0,241,0,7,0,163,0,61,0,183,0,26,0,0,0,114,0,31,0,190,0,69,0,123,0,222,0,47,0,158,0,17,0,187,0,129,0,92,0,252,0,0,0,120,0,0,0,117,0,196,0,177,0,186,0,212,0,232,0,235,0,212,0,90,0,17,0,41,0,128,0,201,0,0,0,94,0,147,0,171,0,0,0,70,0,116,0,90,0,169,0,66,0,165,0,22,0,248,0,28,0,34,0,75,0,89,0,0,0,0,0,20,0,100,0,19,0,197,0,0,0,215,0,255,0,134,0,0,0,63,0,240,0,0,0,70,0,228,0,142,0,103,0,46,0,192,0,213,0,0,0,132,0,37,0,84,0,53,0,0,0,209,0,123,0,0,0,168,0,244,0,39,0,158,0,1,0,0,0,214,0,214,0,95,0,241,0,74,0,43,0,0,0,11,0,251,0,0,0,239,0,62,0,135,0,108,0,29,0,250,0,81,0,255,0,110,0,0,0,50,0,94,0,246,0,144,0,0,0,0,0,0,0,72,0,0,0,166,0,231,0,0,0,34,0,0,0,0,0,174,0,237,0,237,0,146,0,47,0,196,0,2,0,208,0,0,0,157,0,176,0,19,0,33,0,108,0,139,0,29,0,234,0,240,0,51,0,136,0,29,0,0,0,151,0,0,0,126,0,151,0,110,0,6,0,133,0,0,0,0,0,0,0,172,0,31,0,74,0,0,0,195,0,0,0,0,0,203,0,0,0,171,0,236,0,34,0,23,0,181,0,0,0,222,0,89,0,159,0,0,0,75,0,244,0,201,0,172,0,67,0,0,0,236,0,159,0,208,0,87,0,138,0,0,0,69,0,131,0,190,0,175,0,108,0,37,0,8,0,232,0,152,0,0,0,11,0,79,0,0,0,0,0,0,0,73,0,113,0,172,0,18,0,0,0,100,0,138,0,9,0,208,0,206,0,70,0,124,0,0,0,211,0,59,0,0,0,150,0,0,0,0,0,17,0,248,0,214,0,196,0,8,0,0,0,0,0,137,0,38,0,13,0,249,0,181,0,135,0,25,0,5,0,216,0,32,0,68,0,0,0,0,0,0,0,76,0,0,0,209,0,83,0,165,0,10,0,22,0,0,0,120,0,0,0,81,0,0,0,32,0,0,0,0,0,153,0,228,0,0,0,240,0,230,0,40,0,228,0,163,0,226,0,2,0,131,0,95,0,147,0,0,0,114,0,210,0,157,0,113,0,63,0,87,0,156,0,0,0,0,0,0,0,221,0,231,0,72,0,182,0,0,0,229,0,95,0,122,0,0,0,0,0,162,0,78,0,0,0,153,0,236,0,254,0,117,0,40,0,19,0,0,0,253,0,20,0,38,0,114,0,49,0,0,0,185,0,0,0,0,0,0,0,40,0,224,0,164,0,0,0,30,0,93,0,229,0,63,0,210,0,185,0,94,0,52,0,109,0,138,0,0,0,156,0,93,0,142,0,250,0,0,0,104,0,92,0,122,0,4,0,214,0,247,0,157,0,88,0,70,0,0,0,0,0,240,0,81,0,93,0,10,0,0,0,193,0,212,0,0,0,235,0,7,0,0,0,107,0,0,0,0,0,112,0,18,0,14,0,93,0,8,0,232,0,84,0,195,0,52,0,0,0,209,0,117,0,164,0,254,0,251,0,68,0,119,0,23,0,135,0,0,0,112,0,201,0,127,0,230,0,0,0,68,0,38,0,30,0,178,0,64,0,0,0,96,0,192,0,0,0,221,0,119,0,151,0,192,0,189,0,100,0,74,0,77,0,17,0,73,0,210,0,83,0,161,0,0,0,99,0,2,0,0,0,0,0,212,0,204,0,29,0,194,0,109,0,207,0,205,0,0,0,6,0,113,0,82,0,145,0,206,0,64,0,249,0,202,0,38,0,0,0,0,0,16,0,218,0,0,0,175,0,0,0,131,0,12,0,80,0,110,0,0,0,0,0,61,0,0,0,57,0,0,0,0,0,6,0,69,0,0,0,197,0,146,0,2,0,0,0,189,0,5,0,0,0,18,0,246,0,160,0,107,0,237,0,174,0,171,0,194,0,12,0,0,0,135,0,0,0,0,0,147,0,0,0,84,0,133,0,0,0,0,0,90,0,243,0,240,0,175,0,254,0,208,0,127,0,162,0,206,0,0,0,48,0,181,0,157,0,126,0,110,0,39,0,126,0,0,0,0,0,167,0,11,0,242,0,3,0,208,0,37,0,78,0,234,0,142,0,250,0,242,0,169,0,37,0,120,0,150,0,0,0,0,0,0,0,168,0,0,0,0,0,97,0,62,0,118,0,0,0,185,0,0,0,0,0,202,0,0,0,96,0,186,0,83,0,0,0,90,0,98,0,102,0,31,0,138,0,68,0,0,0,63,0,0,0,24,0,158,0,8,0,215,0,146,0,80,0,98,0,163,0,93,0,242,0,0,0,166,0,39,0,148,0,0,0,72,0,102,0,4,0,107,0,44,0,234,0,184,0,175,0,183,0,49,0,0,0,98,0,34,0,0,0,55,0,227,0,251,0,6,0,223,0,3,0,0,0,90,0,8,0,0,0,140,0,52,0,25,0,75,0,0,0,48,0,234,0,154,0,243,0,70,0,59,0,14,0,0,0,121,0,88,0,198,0,113,0,231,0,101,0,58,0,0,0,218,0,153,0,156,0,41,0,240,0,5,0,0,0,87,0,249,0,152,0,94,0,132,0,7,0,181,0,58,0,19,0,7,0,209,0,149,0,156,0,53,0,205,0,94,0,63,0,7,0,90,0,108,0,27,0,0,0,126,0,49,0,202,0,0,0,195,0,47,0,67,0,255,0,77,0,64,0,0,0,0,0,17,0,169,0,226,0,220,0,200,0,252,0,11,0,0,0,0,0,34,0,235,0,0,0,216,0,19,0,245,0,211,0,29,0,63,0,26,0,123,0,196,0,61,0,182,0,0,0,235,0,210,0,41,0,218,0,89,0,164,0,0,0,119,0,155,0,151,0,164,0,2,0,216,0,94,0,136,0,86,0,165,0,212,0,0,0,170,0,64,0,61,0,153,0,117,0,0,0,240,0,44,0,20,0,49,0,78,0,70,0,35,0,77,0,187,0,65,0,117,0,251,0,0,0,207,0,139,0,227,0,15,0,2,0,96,0,112,0,91,0,0,0,239,0,27,0,115,0,37,0,12,0,42,0);
signal scenario_full  : scenario_type := (37,31,41,31,41,30,41,29,192,31,229,31,182,31,91,31,17,31,149,31,40,31,38,31,38,30,215,31,69,31,43,31,56,31,56,30,244,31,25,31,84,31,159,31,168,31,99,31,157,31,222,31,190,31,190,30,37,31,104,31,214,31,143,31,216,31,172,31,151,31,11,31,11,30,194,31,194,30,231,31,213,31,212,31,234,31,188,31,204,31,204,30,231,31,162,31,123,31,108,31,114,31,16,31,165,31,3,31,3,30,128,31,217,31,217,30,253,31,18,31,196,31,11,31,11,30,110,31,190,31,16,31,207,31,207,30,84,31,38,31,38,30,5,31,106,31,106,30,220,31,10,31,168,31,35,31,230,31,149,31,100,31,100,30,100,29,100,28,188,31,116,31,208,31,18,31,87,31,87,30,234,31,107,31,131,31,157,31,157,30,245,31,245,30,245,29,62,31,164,31,171,31,179,31,207,31,234,31,119,31,198,31,198,30,208,31,115,31,73,31,91,31,156,31,156,30,209,31,126,31,5,31,52,31,80,31,21,31,128,31,128,30,196,31,102,31,102,30,63,31,54,31,54,30,211,31,211,30,91,31,136,31,136,30,136,29,136,28,180,31,208,31,230,31,134,31,100,31,100,30,100,29,99,31,79,31,65,31,203,31,203,30,52,31,14,31,115,31,215,31,215,30,255,31,190,31,145,31,95,31,224,31,224,30,126,31,126,30,54,31,87,31,87,30,82,31,82,30,82,29,27,31,170,31,105,31,79,31,25,31,25,30,25,29,25,28,186,31,141,31,141,30,81,31,81,30,114,31,114,30,233,31,196,31,174,31,31,31,246,31,159,31,81,31,96,31,176,31,237,31,245,31,35,31,198,31,60,31,16,31,16,30,155,31,144,31,144,30,24,31,11,31,199,31,157,31,157,31,157,30,6,31,182,31,154,31,154,30,89,31,21,31,122,31,163,31,173,31,169,31,10,31,32,31,103,31,103,30,210,31,232,31,32,31,148,31,212,31,247,31,135,31,4,31,4,30,4,29,149,31,254,31,254,30,123,31,170,31,21,31,82,31,168,31,168,30,231,31,203,31,8,31,8,30,242,31,226,31,226,30,2,31,40,31,187,31,112,31,52,31,67,31,72,31,72,30,72,29,229,31,149,31,149,30,85,31,141,31,103,31,114,31,44,31,126,31,135,31,241,31,7,31,163,31,61,31,183,31,26,31,26,30,114,31,31,31,190,31,69,31,123,31,222,31,47,31,158,31,17,31,187,31,129,31,92,31,252,31,252,30,120,31,120,30,117,31,196,31,177,31,186,31,212,31,232,31,235,31,212,31,90,31,17,31,41,31,128,31,201,31,201,30,94,31,147,31,171,31,171,30,70,31,116,31,90,31,169,31,66,31,165,31,22,31,248,31,28,31,34,31,75,31,89,31,89,30,89,29,20,31,100,31,19,31,197,31,197,30,215,31,255,31,134,31,134,30,63,31,240,31,240,30,70,31,228,31,142,31,103,31,46,31,192,31,213,31,213,30,132,31,37,31,84,31,53,31,53,30,209,31,123,31,123,30,168,31,244,31,39,31,158,31,1,31,1,30,214,31,214,31,95,31,241,31,74,31,43,31,43,30,11,31,251,31,251,30,239,31,62,31,135,31,108,31,29,31,250,31,81,31,255,31,110,31,110,30,50,31,94,31,246,31,144,31,144,30,144,29,144,28,72,31,72,30,166,31,231,31,231,30,34,31,34,30,34,29,174,31,237,31,237,31,146,31,47,31,196,31,2,31,208,31,208,30,157,31,176,31,19,31,33,31,108,31,139,31,29,31,234,31,240,31,51,31,136,31,29,31,29,30,151,31,151,30,126,31,151,31,110,31,6,31,133,31,133,30,133,29,133,28,172,31,31,31,74,31,74,30,195,31,195,30,195,29,203,31,203,30,171,31,236,31,34,31,23,31,181,31,181,30,222,31,89,31,159,31,159,30,75,31,244,31,201,31,172,31,67,31,67,30,236,31,159,31,208,31,87,31,138,31,138,30,69,31,131,31,190,31,175,31,108,31,37,31,8,31,232,31,152,31,152,30,11,31,79,31,79,30,79,29,79,28,73,31,113,31,172,31,18,31,18,30,100,31,138,31,9,31,208,31,206,31,70,31,124,31,124,30,211,31,59,31,59,30,150,31,150,30,150,29,17,31,248,31,214,31,196,31,8,31,8,30,8,29,137,31,38,31,13,31,249,31,181,31,135,31,25,31,5,31,216,31,32,31,68,31,68,30,68,29,68,28,76,31,76,30,209,31,83,31,165,31,10,31,22,31,22,30,120,31,120,30,81,31,81,30,32,31,32,30,32,29,153,31,228,31,228,30,240,31,230,31,40,31,228,31,163,31,226,31,2,31,131,31,95,31,147,31,147,30,114,31,210,31,157,31,113,31,63,31,87,31,156,31,156,30,156,29,156,28,221,31,231,31,72,31,182,31,182,30,229,31,95,31,122,31,122,30,122,29,162,31,78,31,78,30,153,31,236,31,254,31,117,31,40,31,19,31,19,30,253,31,20,31,38,31,114,31,49,31,49,30,185,31,185,30,185,29,185,28,40,31,224,31,164,31,164,30,30,31,93,31,229,31,63,31,210,31,185,31,94,31,52,31,109,31,138,31,138,30,156,31,93,31,142,31,250,31,250,30,104,31,92,31,122,31,4,31,214,31,247,31,157,31,88,31,70,31,70,30,70,29,240,31,81,31,93,31,10,31,10,30,193,31,212,31,212,30,235,31,7,31,7,30,107,31,107,30,107,29,112,31,18,31,14,31,93,31,8,31,232,31,84,31,195,31,52,31,52,30,209,31,117,31,164,31,254,31,251,31,68,31,119,31,23,31,135,31,135,30,112,31,201,31,127,31,230,31,230,30,68,31,38,31,30,31,178,31,64,31,64,30,96,31,192,31,192,30,221,31,119,31,151,31,192,31,189,31,100,31,74,31,77,31,17,31,73,31,210,31,83,31,161,31,161,30,99,31,2,31,2,30,2,29,212,31,204,31,29,31,194,31,109,31,207,31,205,31,205,30,6,31,113,31,82,31,145,31,206,31,64,31,249,31,202,31,38,31,38,30,38,29,16,31,218,31,218,30,175,31,175,30,131,31,12,31,80,31,110,31,110,30,110,29,61,31,61,30,57,31,57,30,57,29,6,31,69,31,69,30,197,31,146,31,2,31,2,30,189,31,5,31,5,30,18,31,246,31,160,31,107,31,237,31,174,31,171,31,194,31,12,31,12,30,135,31,135,30,135,29,147,31,147,30,84,31,133,31,133,30,133,29,90,31,243,31,240,31,175,31,254,31,208,31,127,31,162,31,206,31,206,30,48,31,181,31,157,31,126,31,110,31,39,31,126,31,126,30,126,29,167,31,11,31,242,31,3,31,208,31,37,31,78,31,234,31,142,31,250,31,242,31,169,31,37,31,120,31,150,31,150,30,150,29,150,28,168,31,168,30,168,29,97,31,62,31,118,31,118,30,185,31,185,30,185,29,202,31,202,30,96,31,186,31,83,31,83,30,90,31,98,31,102,31,31,31,138,31,68,31,68,30,63,31,63,30,24,31,158,31,8,31,215,31,146,31,80,31,98,31,163,31,93,31,242,31,242,30,166,31,39,31,148,31,148,30,72,31,102,31,4,31,107,31,44,31,234,31,184,31,175,31,183,31,49,31,49,30,98,31,34,31,34,30,55,31,227,31,251,31,6,31,223,31,3,31,3,30,90,31,8,31,8,30,140,31,52,31,25,31,75,31,75,30,48,31,234,31,154,31,243,31,70,31,59,31,14,31,14,30,121,31,88,31,198,31,113,31,231,31,101,31,58,31,58,30,218,31,153,31,156,31,41,31,240,31,5,31,5,30,87,31,249,31,152,31,94,31,132,31,7,31,181,31,58,31,19,31,7,31,209,31,149,31,156,31,53,31,205,31,94,31,63,31,7,31,90,31,108,31,27,31,27,30,126,31,49,31,202,31,202,30,195,31,47,31,67,31,255,31,77,31,64,31,64,30,64,29,17,31,169,31,226,31,220,31,200,31,252,31,11,31,11,30,11,29,34,31,235,31,235,30,216,31,19,31,245,31,211,31,29,31,63,31,26,31,123,31,196,31,61,31,182,31,182,30,235,31,210,31,41,31,218,31,89,31,164,31,164,30,119,31,155,31,151,31,164,31,2,31,216,31,94,31,136,31,86,31,165,31,212,31,212,30,170,31,64,31,61,31,153,31,117,31,117,30,240,31,44,31,20,31,49,31,78,31,70,31,35,31,77,31,187,31,65,31,117,31,251,31,251,30,207,31,139,31,227,31,15,31,2,31,96,31,112,31,91,31,91,30,239,31,27,31,115,31,37,31,12,31,42,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
