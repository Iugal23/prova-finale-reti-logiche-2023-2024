-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_693 is
end project_tb_693;

architecture project_tb_arch_693 of project_tb_693 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 793;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (135,0,93,0,106,0,103,0,0,0,231,0,0,0,64,0,253,0,234,0,72,0,194,0,209,0,250,0,247,0,29,0,13,0,68,0,0,0,161,0,195,0,67,0,112,0,19,0,251,0,146,0,37,0,0,0,239,0,153,0,34,0,66,0,0,0,0,0,148,0,128,0,239,0,77,0,186,0,183,0,0,0,121,0,198,0,38,0,54,0,131,0,156,0,238,0,212,0,97,0,128,0,25,0,59,0,5,0,34,0,63,0,191,0,201,0,53,0,172,0,0,0,111,0,249,0,0,0,12,0,243,0,6,0,26,0,67,0,139,0,233,0,0,0,0,0,36,0,0,0,180,0,252,0,141,0,240,0,13,0,141,0,0,0,167,0,0,0,124,0,53,0,163,0,92,0,0,0,2,0,9,0,220,0,13,0,0,0,233,0,228,0,0,0,99,0,162,0,193,0,9,0,20,0,9,0,108,0,45,0,60,0,199,0,81,0,0,0,45,0,161,0,154,0,30,0,78,0,124,0,244,0,169,0,35,0,173,0,209,0,48,0,22,0,0,0,226,0,241,0,156,0,174,0,232,0,1,0,0,0,46,0,24,0,220,0,132,0,180,0,148,0,0,0,28,0,138,0,189,0,0,0,125,0,9,0,135,0,187,0,145,0,17,0,0,0,79,0,150,0,191,0,73,0,123,0,199,0,0,0,0,0,0,0,55,0,73,0,94,0,186,0,0,0,0,0,0,0,0,0,0,0,180,0,0,0,27,0,153,0,134,0,95,0,140,0,105,0,70,0,53,0,174,0,130,0,251,0,14,0,155,0,2,0,76,0,12,0,207,0,27,0,27,0,0,0,43,0,157,0,62,0,183,0,113,0,0,0,227,0,160,0,0,0,0,0,134,0,135,0,58,0,223,0,30,0,0,0,179,0,0,0,34,0,226,0,250,0,0,0,116,0,187,0,109,0,179,0,103,0,10,0,180,0,94,0,120,0,128,0,107,0,67,0,75,0,0,0,146,0,177,0,66,0,79,0,248,0,16,0,67,0,235,0,65,0,13,0,130,0,147,0,146,0,228,0,0,0,30,0,60,0,229,0,236,0,62,0,13,0,9,0,185,0,255,0,98,0,27,0,17,0,192,0,244,0,221,0,160,0,0,0,0,0,74,0,54,0,101,0,197,0,113,0,0,0,108,0,154,0,0,0,138,0,0,0,60,0,90,0,18,0,234,0,134,0,26,0,152,0,44,0,153,0,154,0,117,0,0,0,237,0,61,0,148,0,35,0,210,0,53,0,36,0,0,0,14,0,5,0,30,0,0,0,141,0,77,0,19,0,201,0,162,0,228,0,59,0,159,0,118,0,245,0,53,0,223,0,10,0,64,0,43,0,88,0,27,0,251,0,170,0,123,0,59,0,228,0,202,0,226,0,235,0,143,0,122,0,43,0,185,0,170,0,78,0,0,0,113,0,191,0,0,0,75,0,191,0,181,0,236,0,0,0,0,0,104,0,157,0,20,0,142,0,0,0,223,0,236,0,115,0,0,0,240,0,198,0,60,0,129,0,116,0,49,0,11,0,226,0,75,0,123,0,0,0,241,0,159,0,0,0,66,0,221,0,0,0,161,0,227,0,17,0,36,0,134,0,87,0,233,0,18,0,48,0,0,0,80,0,0,0,0,0,194,0,83,0,213,0,137,0,94,0,152,0,0,0,0,0,71,0,34,0,113,0,59,0,25,0,111,0,0,0,132,0,157,0,0,0,0,0,122,0,92,0,128,0,76,0,0,0,185,0,163,0,222,0,186,0,140,0,73,0,0,0,240,0,114,0,137,0,195,0,8,0,253,0,0,0,56,0,29,0,95,0,61,0,234,0,151,0,0,0,250,0,0,0,65,0,70,0,159,0,12,0,79,0,0,0,93,0,22,0,49,0,0,0,106,0,126,0,159,0,249,0,81,0,0,0,121,0,45,0,230,0,145,0,199,0,9,0,183,0,165,0,171,0,45,0,230,0,231,0,254,0,178,0,36,0,241,0,0,0,191,0,172,0,105,0,164,0,2,0,59,0,170,0,103,0,17,0,22,0,0,0,230,0,132,0,109,0,90,0,0,0,124,0,208,0,85,0,133,0,0,0,160,0,153,0,94,0,41,0,11,0,180,0,133,0,184,0,48,0,245,0,0,0,57,0,16,0,236,0,250,0,42,0,36,0,0,0,120,0,162,0,199,0,0,0,227,0,230,0,235,0,0,0,21,0,206,0,174,0,0,0,0,0,115,0,108,0,77,0,0,0,80,0,59,0,34,0,0,0,239,0,155,0,0,0,146,0,38,0,0,0,0,0,59,0,77,0,0,0,0,0,194,0,253,0,207,0,199,0,185,0,84,0,134,0,128,0,164,0,43,0,0,0,19,0,213,0,0,0,0,0,140,0,17,0,0,0,48,0,0,0,211,0,176,0,225,0,252,0,210,0,243,0,23,0,71,0,74,0,116,0,62,0,173,0,0,0,0,0,176,0,245,0,106,0,80,0,73,0,18,0,183,0,0,0,67,0,0,0,47,0,33,0,1,0,220,0,151,0,12,0,230,0,137,0,131,0,168,0,89,0,187,0,0,0,218,0,8,0,82,0,32,0,203,0,143,0,5,0,138,0,225,0,185,0,0,0,29,0,0,0,128,0,50,0,0,0,120,0,128,0,55,0,192,0,100,0,210,0,199,0,67,0,229,0,37,0,86,0,154,0,55,0,198,0,244,0,97,0,36,0,215,0,95,0,0,0,26,0,0,0,74,0,111,0,36,0,0,0,0,0,161,0,13,0,136,0,60,0,0,0,138,0,0,0,159,0,0,0,67,0,209,0,0,0,147,0,236,0,222,0,22,0,195,0,0,0,205,0,185,0,59,0,151,0,118,0,111,0,11,0,241,0,75,0,221,0,35,0,17,0,0,0,247,0,0,0,0,0,89,0,93,0,253,0,70,0,157,0,170,0,245,0,132,0,125,0,53,0,243,0,92,0,0,0,0,0,214,0,134,0,62,0,63,0,174,0,202,0,28,0,158,0,8,0,231,0,227,0,223,0,35,0,220,0,21,0,123,0,45,0,0,0,51,0,251,0,146,0,114,0,213,0,224,0,0,0,219,0,242,0,96,0,150,0,209,0,34,0,28,0,38,0,224,0,0,0,68,0,0,0,0,0,64,0,0,0,239,0,0,0,0,0,95,0,130,0,202,0,142,0,104,0,33,0,0,0,240,0,17,0,157,0,170,0,0,0,0,0,221,0,115,0,48,0,125,0,11,0,0,0,138,0,63,0,34,0,157,0,0,0,0,0,208,0,238,0,90,0,199,0,0,0,0,0,78,0,108,0,0,0,203,0,55,0,188,0,140,0,75,0,7,0,187,0,128,0,0,0,31,0,44,0,46,0,75,0,254,0,0,0,115,0,110,0,73,0,102,0,0,0,214,0,235,0,141,0,154,0,161,0,230,0,34,0,134,0,0,0,18,0,40,0,0,0,185,0,0,0,111,0,153,0,17,0,0,0,193,0,230,0,83,0,233,0,78,0,166,0,224,0);
signal scenario_full  : scenario_type := (135,31,93,31,106,31,103,31,103,30,231,31,231,30,64,31,253,31,234,31,72,31,194,31,209,31,250,31,247,31,29,31,13,31,68,31,68,30,161,31,195,31,67,31,112,31,19,31,251,31,146,31,37,31,37,30,239,31,153,31,34,31,66,31,66,30,66,29,148,31,128,31,239,31,77,31,186,31,183,31,183,30,121,31,198,31,38,31,54,31,131,31,156,31,238,31,212,31,97,31,128,31,25,31,59,31,5,31,34,31,63,31,191,31,201,31,53,31,172,31,172,30,111,31,249,31,249,30,12,31,243,31,6,31,26,31,67,31,139,31,233,31,233,30,233,29,36,31,36,30,180,31,252,31,141,31,240,31,13,31,141,31,141,30,167,31,167,30,124,31,53,31,163,31,92,31,92,30,2,31,9,31,220,31,13,31,13,30,233,31,228,31,228,30,99,31,162,31,193,31,9,31,20,31,9,31,108,31,45,31,60,31,199,31,81,31,81,30,45,31,161,31,154,31,30,31,78,31,124,31,244,31,169,31,35,31,173,31,209,31,48,31,22,31,22,30,226,31,241,31,156,31,174,31,232,31,1,31,1,30,46,31,24,31,220,31,132,31,180,31,148,31,148,30,28,31,138,31,189,31,189,30,125,31,9,31,135,31,187,31,145,31,17,31,17,30,79,31,150,31,191,31,73,31,123,31,199,31,199,30,199,29,199,28,55,31,73,31,94,31,186,31,186,30,186,29,186,28,186,27,186,26,180,31,180,30,27,31,153,31,134,31,95,31,140,31,105,31,70,31,53,31,174,31,130,31,251,31,14,31,155,31,2,31,76,31,12,31,207,31,27,31,27,31,27,30,43,31,157,31,62,31,183,31,113,31,113,30,227,31,160,31,160,30,160,29,134,31,135,31,58,31,223,31,30,31,30,30,179,31,179,30,34,31,226,31,250,31,250,30,116,31,187,31,109,31,179,31,103,31,10,31,180,31,94,31,120,31,128,31,107,31,67,31,75,31,75,30,146,31,177,31,66,31,79,31,248,31,16,31,67,31,235,31,65,31,13,31,130,31,147,31,146,31,228,31,228,30,30,31,60,31,229,31,236,31,62,31,13,31,9,31,185,31,255,31,98,31,27,31,17,31,192,31,244,31,221,31,160,31,160,30,160,29,74,31,54,31,101,31,197,31,113,31,113,30,108,31,154,31,154,30,138,31,138,30,60,31,90,31,18,31,234,31,134,31,26,31,152,31,44,31,153,31,154,31,117,31,117,30,237,31,61,31,148,31,35,31,210,31,53,31,36,31,36,30,14,31,5,31,30,31,30,30,141,31,77,31,19,31,201,31,162,31,228,31,59,31,159,31,118,31,245,31,53,31,223,31,10,31,64,31,43,31,88,31,27,31,251,31,170,31,123,31,59,31,228,31,202,31,226,31,235,31,143,31,122,31,43,31,185,31,170,31,78,31,78,30,113,31,191,31,191,30,75,31,191,31,181,31,236,31,236,30,236,29,104,31,157,31,20,31,142,31,142,30,223,31,236,31,115,31,115,30,240,31,198,31,60,31,129,31,116,31,49,31,11,31,226,31,75,31,123,31,123,30,241,31,159,31,159,30,66,31,221,31,221,30,161,31,227,31,17,31,36,31,134,31,87,31,233,31,18,31,48,31,48,30,80,31,80,30,80,29,194,31,83,31,213,31,137,31,94,31,152,31,152,30,152,29,71,31,34,31,113,31,59,31,25,31,111,31,111,30,132,31,157,31,157,30,157,29,122,31,92,31,128,31,76,31,76,30,185,31,163,31,222,31,186,31,140,31,73,31,73,30,240,31,114,31,137,31,195,31,8,31,253,31,253,30,56,31,29,31,95,31,61,31,234,31,151,31,151,30,250,31,250,30,65,31,70,31,159,31,12,31,79,31,79,30,93,31,22,31,49,31,49,30,106,31,126,31,159,31,249,31,81,31,81,30,121,31,45,31,230,31,145,31,199,31,9,31,183,31,165,31,171,31,45,31,230,31,231,31,254,31,178,31,36,31,241,31,241,30,191,31,172,31,105,31,164,31,2,31,59,31,170,31,103,31,17,31,22,31,22,30,230,31,132,31,109,31,90,31,90,30,124,31,208,31,85,31,133,31,133,30,160,31,153,31,94,31,41,31,11,31,180,31,133,31,184,31,48,31,245,31,245,30,57,31,16,31,236,31,250,31,42,31,36,31,36,30,120,31,162,31,199,31,199,30,227,31,230,31,235,31,235,30,21,31,206,31,174,31,174,30,174,29,115,31,108,31,77,31,77,30,80,31,59,31,34,31,34,30,239,31,155,31,155,30,146,31,38,31,38,30,38,29,59,31,77,31,77,30,77,29,194,31,253,31,207,31,199,31,185,31,84,31,134,31,128,31,164,31,43,31,43,30,19,31,213,31,213,30,213,29,140,31,17,31,17,30,48,31,48,30,211,31,176,31,225,31,252,31,210,31,243,31,23,31,71,31,74,31,116,31,62,31,173,31,173,30,173,29,176,31,245,31,106,31,80,31,73,31,18,31,183,31,183,30,67,31,67,30,47,31,33,31,1,31,220,31,151,31,12,31,230,31,137,31,131,31,168,31,89,31,187,31,187,30,218,31,8,31,82,31,32,31,203,31,143,31,5,31,138,31,225,31,185,31,185,30,29,31,29,30,128,31,50,31,50,30,120,31,128,31,55,31,192,31,100,31,210,31,199,31,67,31,229,31,37,31,86,31,154,31,55,31,198,31,244,31,97,31,36,31,215,31,95,31,95,30,26,31,26,30,74,31,111,31,36,31,36,30,36,29,161,31,13,31,136,31,60,31,60,30,138,31,138,30,159,31,159,30,67,31,209,31,209,30,147,31,236,31,222,31,22,31,195,31,195,30,205,31,185,31,59,31,151,31,118,31,111,31,11,31,241,31,75,31,221,31,35,31,17,31,17,30,247,31,247,30,247,29,89,31,93,31,253,31,70,31,157,31,170,31,245,31,132,31,125,31,53,31,243,31,92,31,92,30,92,29,214,31,134,31,62,31,63,31,174,31,202,31,28,31,158,31,8,31,231,31,227,31,223,31,35,31,220,31,21,31,123,31,45,31,45,30,51,31,251,31,146,31,114,31,213,31,224,31,224,30,219,31,242,31,96,31,150,31,209,31,34,31,28,31,38,31,224,31,224,30,68,31,68,30,68,29,64,31,64,30,239,31,239,30,239,29,95,31,130,31,202,31,142,31,104,31,33,31,33,30,240,31,17,31,157,31,170,31,170,30,170,29,221,31,115,31,48,31,125,31,11,31,11,30,138,31,63,31,34,31,157,31,157,30,157,29,208,31,238,31,90,31,199,31,199,30,199,29,78,31,108,31,108,30,203,31,55,31,188,31,140,31,75,31,7,31,187,31,128,31,128,30,31,31,44,31,46,31,75,31,254,31,254,30,115,31,110,31,73,31,102,31,102,30,214,31,235,31,141,31,154,31,161,31,230,31,34,31,134,31,134,30,18,31,40,31,40,30,185,31,185,30,111,31,153,31,17,31,17,30,193,31,230,31,83,31,233,31,78,31,166,31,224,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
