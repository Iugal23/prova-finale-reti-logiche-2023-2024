-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 183;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (102,0,252,0,150,0,185,0,191,0,0,0,66,0,85,0,143,0,245,0,0,0,138,0,56,0,246,0,135,0,0,0,60,0,239,0,89,0,128,0,204,0,161,0,241,0,254,0,0,0,120,0,246,0,0,0,7,0,42,0,126,0,30,0,13,0,49,0,121,0,243,0,85,0,0,0,0,0,17,0,0,0,59,0,143,0,245,0,43,0,217,0,127,0,237,0,211,0,0,0,0,0,0,0,54,0,0,0,133,0,177,0,0,0,246,0,217,0,75,0,68,0,16,0,237,0,223,0,236,0,128,0,32,0,0,0,70,0,133,0,28,0,226,0,0,0,55,0,208,0,70,0,193,0,0,0,45,0,0,0,207,0,116,0,239,0,0,0,236,0,0,0,6,0,175,0,0,0,123,0,176,0,227,0,129,0,0,0,124,0,180,0,32,0,103,0,103,0,21,0,31,0,243,0,121,0,105,0,5,0,251,0,41,0,100,0,82,0,22,0,132,0,190,0,93,0,232,0,211,0,32,0,11,0,0,0,201,0,183,0,193,0,20,0,235,0,225,0,0,0,91,0,0,0,119,0,179,0,95,0,148,0,0,0,7,0,19,0,245,0,0,0,243,0,184,0,255,0,129,0,0,0,247,0,154,0,203,0,53,0,7,0,190,0,22,0,163,0,222,0,209,0,1,0,0,0,111,0,147,0,177,0,191,0,25,0,80,0,227,0,197,0,198,0,193,0,219,0,1,0,53,0,196,0,10,0,106,0,157,0,0,0,4,0,0,0,0,0,139,0,203,0,0,0,217,0,178,0,144,0,125,0,218,0,80,0);
signal scenario_full  : scenario_type := (102,31,252,31,150,31,185,31,191,31,191,30,66,31,85,31,143,31,245,31,245,30,138,31,56,31,246,31,135,31,135,30,60,31,239,31,89,31,128,31,204,31,161,31,241,31,254,31,254,30,120,31,246,31,246,30,7,31,42,31,126,31,30,31,13,31,49,31,121,31,243,31,85,31,85,30,85,29,17,31,17,30,59,31,143,31,245,31,43,31,217,31,127,31,237,31,211,31,211,30,211,29,211,28,54,31,54,30,133,31,177,31,177,30,246,31,217,31,75,31,68,31,16,31,237,31,223,31,236,31,128,31,32,31,32,30,70,31,133,31,28,31,226,31,226,30,55,31,208,31,70,31,193,31,193,30,45,31,45,30,207,31,116,31,239,31,239,30,236,31,236,30,6,31,175,31,175,30,123,31,176,31,227,31,129,31,129,30,124,31,180,31,32,31,103,31,103,31,21,31,31,31,243,31,121,31,105,31,5,31,251,31,41,31,100,31,82,31,22,31,132,31,190,31,93,31,232,31,211,31,32,31,11,31,11,30,201,31,183,31,193,31,20,31,235,31,225,31,225,30,91,31,91,30,119,31,179,31,95,31,148,31,148,30,7,31,19,31,245,31,245,30,243,31,184,31,255,31,129,31,129,30,247,31,154,31,203,31,53,31,7,31,190,31,22,31,163,31,222,31,209,31,1,31,1,30,111,31,147,31,177,31,191,31,25,31,80,31,227,31,197,31,198,31,193,31,219,31,1,31,53,31,196,31,10,31,106,31,157,31,157,30,4,31,4,30,4,29,139,31,203,31,203,30,217,31,178,31,144,31,125,31,218,31,80,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
