-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_339 is
end project_tb_339;

architecture project_tb_arch_339 of project_tb_339 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 629;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (197,0,0,0,0,0,85,0,177,0,74,0,109,0,95,0,193,0,0,0,122,0,184,0,88,0,204,0,222,0,71,0,226,0,110,0,0,0,221,0,176,0,160,0,37,0,122,0,173,0,109,0,69,0,10,0,61,0,54,0,0,0,111,0,0,0,117,0,0,0,189,0,200,0,0,0,43,0,0,0,251,0,206,0,0,0,159,0,124,0,207,0,0,0,175,0,58,0,170,0,75,0,78,0,227,0,0,0,43,0,237,0,7,0,237,0,57,0,245,0,0,0,0,0,17,0,179,0,51,0,157,0,107,0,158,0,22,0,66,0,109,0,88,0,134,0,191,0,223,0,224,0,240,0,0,0,144,0,232,0,0,0,70,0,113,0,200,0,37,0,244,0,46,0,168,0,48,0,80,0,130,0,228,0,115,0,171,0,0,0,23,0,160,0,237,0,167,0,123,0,91,0,17,0,99,0,88,0,114,0,90,0,40,0,0,0,137,0,65,0,48,0,0,0,24,0,184,0,34,0,165,0,193,0,0,0,33,0,221,0,202,0,233,0,190,0,106,0,126,0,217,0,194,0,22,0,100,0,56,0,83,0,0,0,241,0,136,0,18,0,135,0,116,0,11,0,0,0,207,0,0,0,75,0,230,0,168,0,244,0,23,0,156,0,177,0,177,0,0,0,151,0,232,0,151,0,149,0,146,0,0,0,78,0,208,0,91,0,158,0,118,0,110,0,249,0,232,0,191,0,217,0,47,0,82,0,0,0,0,0,185,0,240,0,0,0,96,0,10,0,0,0,118,0,42,0,84,0,0,0,156,0,33,0,127,0,247,0,129,0,0,0,174,0,40,0,187,0,249,0,9,0,147,0,0,0,162,0,76,0,0,0,67,0,31,0,0,0,102,0,235,0,245,0,67,0,223,0,97,0,205,0,186,0,152,0,0,0,217,0,0,0,161,0,13,0,138,0,0,0,189,0,0,0,222,0,74,0,101,0,147,0,69,0,45,0,0,0,247,0,236,0,123,0,150,0,66,0,207,0,212,0,82,0,206,0,122,0,126,0,149,0,47,0,202,0,0,0,219,0,237,0,24,0,74,0,204,0,94,0,181,0,234,0,0,0,96,0,160,0,103,0,224,0,5,0,0,0,39,0,202,0,106,0,251,0,0,0,231,0,101,0,206,0,182,0,137,0,201,0,63,0,0,0,164,0,0,0,149,0,10,0,200,0,0,0,127,0,192,0,228,0,60,0,238,0,255,0,38,0,156,0,85,0,244,0,182,0,37,0,21,0,149,0,82,0,192,0,125,0,220,0,0,0,5,0,123,0,178,0,198,0,0,0,164,0,0,0,155,0,61,0,0,0,81,0,67,0,13,0,96,0,0,0,8,0,76,0,169,0,168,0,7,0,112,0,185,0,0,0,240,0,105,0,114,0,62,0,129,0,44,0,0,0,218,0,139,0,198,0,98,0,121,0,41,0,151,0,0,0,105,0,149,0,253,0,89,0,191,0,0,0,0,0,29,0,0,0,0,0,0,0,226,0,66,0,52,0,174,0,119,0,112,0,228,0,237,0,0,0,231,0,0,0,0,0,102,0,0,0,26,0,117,0,236,0,234,0,102,0,0,0,141,0,0,0,246,0,177,0,128,0,0,0,0,0,215,0,25,0,144,0,123,0,37,0,228,0,31,0,0,0,133,0,0,0,137,0,21,0,0,0,120,0,201,0,106,0,4,0,241,0,16,0,97,0,204,0,53,0,235,0,134,0,171,0,193,0,24,0,192,0,0,0,42,0,244,0,177,0,187,0,0,0,0,0,232,0,84,0,9,0,0,0,214,0,84,0,247,0,220,0,0,0,119,0,245,0,147,0,0,0,241,0,255,0,33,0,0,0,23,0,211,0,0,0,225,0,88,0,98,0,115,0,181,0,173,0,0,0,39,0,97,0,197,0,171,0,80,0,0,0,179,0,90,0,232,0,57,0,0,0,0,0,214,0,167,0,28,0,124,0,71,0,0,0,248,0,8,0,225,0,0,0,3,0,131,0,0,0,200,0,3,0,51,0,244,0,193,0,247,0,109,0,225,0,220,0,0,0,0,0,23,0,193,0,91,0,93,0,167,0,0,0,164,0,0,0,235,0,56,0,35,0,10,0,0,0,173,0,25,0,123,0,95,0,49,0,131,0,148,0,243,0,175,0,130,0,0,0,0,0,0,0,13,0,0,0,235,0,87,0,15,0,0,0,137,0,1,0,14,0,225,0,189,0,238,0,0,0,83,0,27,0,0,0,182,0,157,0,173,0,174,0,5,0,240,0,86,0,0,0,152,0,224,0,232,0,64,0,166,0,204,0,96,0,13,0,222,0,0,0,0,0,221,0,73,0,97,0,4,0,0,0,9,0,246,0,86,0,177,0,49,0,142,0,63,0,157,0,0,0,32,0,0,0,89,0,230,0,62,0,46,0,180,0,213,0,61,0,233,0,141,0,0,0,112,0,83,0,25,0,189,0,180,0,58,0,254,0,35,0,111,0,93,0,0,0,172,0,221,0,0,0,0,0,14,0,93,0,0,0,92,0,24,0,214,0,22,0,51,0,124,0,0,0,0,0,13,0,16,0,163,0,45,0,26,0,174,0,246,0,41,0,118,0,206,0,236,0,248,0,135,0,0,0,141,0,145,0,145,0,138,0,228,0,64,0,242,0,0,0,78,0,252,0,115,0,137,0,16,0,221,0,52,0,202,0,0,0,169,0,136,0,173,0,125,0,195,0,39,0,255,0,44,0,53,0,153,0,163,0,89,0,54,0,188,0,213,0,81,0,44,0,47,0,17,0);
signal scenario_full  : scenario_type := (197,31,197,30,197,29,85,31,177,31,74,31,109,31,95,31,193,31,193,30,122,31,184,31,88,31,204,31,222,31,71,31,226,31,110,31,110,30,221,31,176,31,160,31,37,31,122,31,173,31,109,31,69,31,10,31,61,31,54,31,54,30,111,31,111,30,117,31,117,30,189,31,200,31,200,30,43,31,43,30,251,31,206,31,206,30,159,31,124,31,207,31,207,30,175,31,58,31,170,31,75,31,78,31,227,31,227,30,43,31,237,31,7,31,237,31,57,31,245,31,245,30,245,29,17,31,179,31,51,31,157,31,107,31,158,31,22,31,66,31,109,31,88,31,134,31,191,31,223,31,224,31,240,31,240,30,144,31,232,31,232,30,70,31,113,31,200,31,37,31,244,31,46,31,168,31,48,31,80,31,130,31,228,31,115,31,171,31,171,30,23,31,160,31,237,31,167,31,123,31,91,31,17,31,99,31,88,31,114,31,90,31,40,31,40,30,137,31,65,31,48,31,48,30,24,31,184,31,34,31,165,31,193,31,193,30,33,31,221,31,202,31,233,31,190,31,106,31,126,31,217,31,194,31,22,31,100,31,56,31,83,31,83,30,241,31,136,31,18,31,135,31,116,31,11,31,11,30,207,31,207,30,75,31,230,31,168,31,244,31,23,31,156,31,177,31,177,31,177,30,151,31,232,31,151,31,149,31,146,31,146,30,78,31,208,31,91,31,158,31,118,31,110,31,249,31,232,31,191,31,217,31,47,31,82,31,82,30,82,29,185,31,240,31,240,30,96,31,10,31,10,30,118,31,42,31,84,31,84,30,156,31,33,31,127,31,247,31,129,31,129,30,174,31,40,31,187,31,249,31,9,31,147,31,147,30,162,31,76,31,76,30,67,31,31,31,31,30,102,31,235,31,245,31,67,31,223,31,97,31,205,31,186,31,152,31,152,30,217,31,217,30,161,31,13,31,138,31,138,30,189,31,189,30,222,31,74,31,101,31,147,31,69,31,45,31,45,30,247,31,236,31,123,31,150,31,66,31,207,31,212,31,82,31,206,31,122,31,126,31,149,31,47,31,202,31,202,30,219,31,237,31,24,31,74,31,204,31,94,31,181,31,234,31,234,30,96,31,160,31,103,31,224,31,5,31,5,30,39,31,202,31,106,31,251,31,251,30,231,31,101,31,206,31,182,31,137,31,201,31,63,31,63,30,164,31,164,30,149,31,10,31,200,31,200,30,127,31,192,31,228,31,60,31,238,31,255,31,38,31,156,31,85,31,244,31,182,31,37,31,21,31,149,31,82,31,192,31,125,31,220,31,220,30,5,31,123,31,178,31,198,31,198,30,164,31,164,30,155,31,61,31,61,30,81,31,67,31,13,31,96,31,96,30,8,31,76,31,169,31,168,31,7,31,112,31,185,31,185,30,240,31,105,31,114,31,62,31,129,31,44,31,44,30,218,31,139,31,198,31,98,31,121,31,41,31,151,31,151,30,105,31,149,31,253,31,89,31,191,31,191,30,191,29,29,31,29,30,29,29,29,28,226,31,66,31,52,31,174,31,119,31,112,31,228,31,237,31,237,30,231,31,231,30,231,29,102,31,102,30,26,31,117,31,236,31,234,31,102,31,102,30,141,31,141,30,246,31,177,31,128,31,128,30,128,29,215,31,25,31,144,31,123,31,37,31,228,31,31,31,31,30,133,31,133,30,137,31,21,31,21,30,120,31,201,31,106,31,4,31,241,31,16,31,97,31,204,31,53,31,235,31,134,31,171,31,193,31,24,31,192,31,192,30,42,31,244,31,177,31,187,31,187,30,187,29,232,31,84,31,9,31,9,30,214,31,84,31,247,31,220,31,220,30,119,31,245,31,147,31,147,30,241,31,255,31,33,31,33,30,23,31,211,31,211,30,225,31,88,31,98,31,115,31,181,31,173,31,173,30,39,31,97,31,197,31,171,31,80,31,80,30,179,31,90,31,232,31,57,31,57,30,57,29,214,31,167,31,28,31,124,31,71,31,71,30,248,31,8,31,225,31,225,30,3,31,131,31,131,30,200,31,3,31,51,31,244,31,193,31,247,31,109,31,225,31,220,31,220,30,220,29,23,31,193,31,91,31,93,31,167,31,167,30,164,31,164,30,235,31,56,31,35,31,10,31,10,30,173,31,25,31,123,31,95,31,49,31,131,31,148,31,243,31,175,31,130,31,130,30,130,29,130,28,13,31,13,30,235,31,87,31,15,31,15,30,137,31,1,31,14,31,225,31,189,31,238,31,238,30,83,31,27,31,27,30,182,31,157,31,173,31,174,31,5,31,240,31,86,31,86,30,152,31,224,31,232,31,64,31,166,31,204,31,96,31,13,31,222,31,222,30,222,29,221,31,73,31,97,31,4,31,4,30,9,31,246,31,86,31,177,31,49,31,142,31,63,31,157,31,157,30,32,31,32,30,89,31,230,31,62,31,46,31,180,31,213,31,61,31,233,31,141,31,141,30,112,31,83,31,25,31,189,31,180,31,58,31,254,31,35,31,111,31,93,31,93,30,172,31,221,31,221,30,221,29,14,31,93,31,93,30,92,31,24,31,214,31,22,31,51,31,124,31,124,30,124,29,13,31,16,31,163,31,45,31,26,31,174,31,246,31,41,31,118,31,206,31,236,31,248,31,135,31,135,30,141,31,145,31,145,31,138,31,228,31,64,31,242,31,242,30,78,31,252,31,115,31,137,31,16,31,221,31,52,31,202,31,202,30,169,31,136,31,173,31,125,31,195,31,39,31,255,31,44,31,53,31,153,31,163,31,89,31,54,31,188,31,213,31,81,31,44,31,47,31,17,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
