-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_703 is
end project_tb_703;

architecture project_tb_arch_703 of project_tb_703 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 292;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,174,0,123,0,187,0,0,0,27,0,207,0,72,0,36,0,151,0,0,0,228,0,0,0,186,0,100,0,152,0,0,0,56,0,234,0,27,0,150,0,44,0,131,0,0,0,233,0,0,0,187,0,140,0,6,0,69,0,6,0,158,0,0,0,0,0,160,0,244,0,207,0,245,0,232,0,206,0,124,0,0,0,25,0,123,0,112,0,216,0,0,0,0,0,127,0,110,0,147,0,0,0,25,0,69,0,0,0,0,0,0,0,0,0,239,0,245,0,146,0,55,0,201,0,0,0,42,0,97,0,33,0,202,0,36,0,147,0,235,0,118,0,65,0,177,0,0,0,79,0,237,0,88,0,45,0,160,0,240,0,6,0,76,0,114,0,61,0,2,0,225,0,187,0,198,0,61,0,154,0,141,0,147,0,98,0,159,0,51,0,128,0,93,0,3,0,121,0,149,0,207,0,175,0,98,0,165,0,183,0,221,0,188,0,0,0,193,0,84,0,126,0,96,0,43,0,29,0,0,0,34,0,211,0,38,0,0,0,111,0,13,0,49,0,18,0,101,0,72,0,115,0,0,0,200,0,146,0,80,0,204,0,142,0,46,0,246,0,0,0,99,0,43,0,217,0,204,0,184,0,0,0,92,0,55,0,255,0,93,0,0,0,140,0,0,0,222,0,0,0,18,0,31,0,180,0,3,0,232,0,67,0,183,0,177,0,69,0,0,0,47,0,0,0,0,0,205,0,0,0,0,0,169,0,200,0,0,0,59,0,28,0,223,0,131,0,65,0,0,0,199,0,0,0,246,0,215,0,125,0,77,0,0,0,0,0,0,0,192,0,35,0,51,0,240,0,36,0,0,0,0,0,0,0,113,0,73,0,0,0,0,0,51,0,201,0,0,0,55,0,23,0,52,0,46,0,237,0,169,0,167,0,0,0,207,0,0,0,0,0,142,0,112,0,0,0,214,0,58,0,163,0,55,0,154,0,198,0,244,0,83,0,89,0,64,0,0,0,252,0,6,0,140,0,188,0,0,0,54,0,243,0,119,0,143,0,67,0,153,0,87,0,157,0,106,0,83,0,60,0,112,0,180,0,114,0,0,0,231,0,154,0,0,0,177,0,81,0,0,0,234,0,192,0,210,0,116,0,106,0,149,0,35,0,89,0,0,0,227,0,160,0,45,0,186,0,75,0,214,0,0,0,2,0,239,0,0,0,159,0,0,0,8,0,232,0,132,0,150,0,101,0,64,0,204,0,60,0,0,0,193,0,244,0,154,0,0,0,201,0,0,0,0,0,245,0,105,0,134,0,41,0);
signal scenario_full  : scenario_type := (0,0,174,31,123,31,187,31,187,30,27,31,207,31,72,31,36,31,151,31,151,30,228,31,228,30,186,31,100,31,152,31,152,30,56,31,234,31,27,31,150,31,44,31,131,31,131,30,233,31,233,30,187,31,140,31,6,31,69,31,6,31,158,31,158,30,158,29,160,31,244,31,207,31,245,31,232,31,206,31,124,31,124,30,25,31,123,31,112,31,216,31,216,30,216,29,127,31,110,31,147,31,147,30,25,31,69,31,69,30,69,29,69,28,69,27,239,31,245,31,146,31,55,31,201,31,201,30,42,31,97,31,33,31,202,31,36,31,147,31,235,31,118,31,65,31,177,31,177,30,79,31,237,31,88,31,45,31,160,31,240,31,6,31,76,31,114,31,61,31,2,31,225,31,187,31,198,31,61,31,154,31,141,31,147,31,98,31,159,31,51,31,128,31,93,31,3,31,121,31,149,31,207,31,175,31,98,31,165,31,183,31,221,31,188,31,188,30,193,31,84,31,126,31,96,31,43,31,29,31,29,30,34,31,211,31,38,31,38,30,111,31,13,31,49,31,18,31,101,31,72,31,115,31,115,30,200,31,146,31,80,31,204,31,142,31,46,31,246,31,246,30,99,31,43,31,217,31,204,31,184,31,184,30,92,31,55,31,255,31,93,31,93,30,140,31,140,30,222,31,222,30,18,31,31,31,180,31,3,31,232,31,67,31,183,31,177,31,69,31,69,30,47,31,47,30,47,29,205,31,205,30,205,29,169,31,200,31,200,30,59,31,28,31,223,31,131,31,65,31,65,30,199,31,199,30,246,31,215,31,125,31,77,31,77,30,77,29,77,28,192,31,35,31,51,31,240,31,36,31,36,30,36,29,36,28,113,31,73,31,73,30,73,29,51,31,201,31,201,30,55,31,23,31,52,31,46,31,237,31,169,31,167,31,167,30,207,31,207,30,207,29,142,31,112,31,112,30,214,31,58,31,163,31,55,31,154,31,198,31,244,31,83,31,89,31,64,31,64,30,252,31,6,31,140,31,188,31,188,30,54,31,243,31,119,31,143,31,67,31,153,31,87,31,157,31,106,31,83,31,60,31,112,31,180,31,114,31,114,30,231,31,154,31,154,30,177,31,81,31,81,30,234,31,192,31,210,31,116,31,106,31,149,31,35,31,89,31,89,30,227,31,160,31,45,31,186,31,75,31,214,31,214,30,2,31,239,31,239,30,159,31,159,30,8,31,232,31,132,31,150,31,101,31,64,31,204,31,60,31,60,30,193,31,244,31,154,31,154,30,201,31,201,30,201,29,245,31,105,31,134,31,41,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
