-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_215 is
end project_tb_215;

architecture project_tb_arch_215 of project_tb_215 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 838;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (60,0,4,0,170,0,90,0,159,0,0,0,198,0,0,0,0,0,0,0,185,0,221,0,75,0,216,0,48,0,35,0,240,0,227,0,144,0,0,0,211,0,195,0,155,0,0,0,0,0,87,0,79,0,150,0,124,0,33,0,57,0,0,0,85,0,0,0,0,0,101,0,65,0,0,0,157,0,147,0,237,0,0,0,194,0,0,0,118,0,151,0,188,0,236,0,14,0,89,0,0,0,54,0,238,0,214,0,215,0,0,0,0,0,193,0,148,0,0,0,172,0,109,0,2,0,0,0,63,0,0,0,23,0,48,0,147,0,124,0,0,0,2,0,204,0,71,0,0,0,17,0,127,0,133,0,4,0,179,0,178,0,0,0,4,0,215,0,0,0,153,0,138,0,0,0,195,0,91,0,0,0,115,0,0,0,0,0,45,0,0,0,85,0,243,0,0,0,143,0,227,0,162,0,239,0,0,0,51,0,0,0,0,0,0,0,136,0,64,0,100,0,25,0,235,0,66,0,0,0,0,0,130,0,137,0,39,0,57,0,0,0,180,0,0,0,185,0,0,0,38,0,2,0,237,0,155,0,169,0,206,0,0,0,23,0,56,0,202,0,0,0,112,0,0,0,19,0,166,0,185,0,119,0,102,0,247,0,65,0,8,0,160,0,92,0,160,0,58,0,0,0,0,0,46,0,151,0,93,0,2,0,0,0,174,0,0,0,207,0,171,0,37,0,45,0,162,0,117,0,47,0,0,0,96,0,25,0,38,0,0,0,252,0,36,0,139,0,0,0,179,0,0,0,192,0,8,0,56,0,235,0,200,0,237,0,62,0,160,0,3,0,218,0,65,0,99,0,189,0,55,0,80,0,14,0,74,0,140,0,204,0,0,0,59,0,0,0,167,0,146,0,68,0,194,0,158,0,60,0,112,0,164,0,172,0,116,0,124,0,0,0,51,0,60,0,242,0,157,0,245,0,183,0,0,0,0,0,31,0,219,0,187,0,0,0,229,0,15,0,0,0,0,0,223,0,221,0,244,0,204,0,227,0,0,0,142,0,20,0,0,0,0,0,92,0,243,0,197,0,252,0,0,0,19,0,0,0,59,0,229,0,171,0,36,0,0,0,226,0,26,0,95,0,44,0,0,0,106,0,0,0,57,0,0,0,184,0,129,0,218,0,75,0,0,0,176,0,0,0,108,0,187,0,170,0,75,0,58,0,227,0,18,0,0,0,205,0,109,0,77,0,45,0,93,0,29,0,176,0,124,0,56,0,38,0,166,0,189,0,0,0,0,0,9,0,36,0,0,0,0,0,0,0,0,0,0,0,49,0,207,0,208,0,51,0,163,0,18,0,31,0,149,0,102,0,39,0,72,0,37,0,220,0,112,0,64,0,148,0,6,0,238,0,159,0,197,0,228,0,118,0,210,0,124,0,0,0,99,0,68,0,243,0,132,0,229,0,0,0,77,0,0,0,0,0,203,0,58,0,102,0,201,0,24,0,129,0,15,0,47,0,0,0,118,0,123,0,47,0,180,0,151,0,37,0,0,0,242,0,13,0,76,0,213,0,113,0,174,0,198,0,195,0,113,0,213,0,0,0,172,0,31,0,223,0,126,0,110,0,131,0,73,0,103,0,123,0,0,0,87,0,99,0,40,0,98,0,248,0,248,0,0,0,69,0,83,0,0,0,58,0,0,0,95,0,237,0,194,0,136,0,236,0,157,0,248,0,190,0,72,0,234,0,216,0,0,0,0,0,142,0,115,0,0,0,0,0,255,0,0,0,0,0,149,0,142,0,0,0,239,0,0,0,23,0,42,0,0,0,246,0,115,0,193,0,122,0,187,0,126,0,0,0,147,0,51,0,219,0,0,0,64,0,255,0,0,0,29,0,144,0,196,0,0,0,68,0,67,0,12,0,151,0,163,0,239,0,169,0,32,0,246,0,0,0,110,0,176,0,16,0,134,0,233,0,95,0,61,0,32,0,104,0,1,0,98,0,10,0,255,0,249,0,68,0,45,0,180,0,3,0,0,0,129,0,89,0,139,0,14,0,0,0,192,0,241,0,0,0,0,0,92,0,0,0,105,0,107,0,80,0,0,0,97,0,0,0,222,0,0,0,94,0,162,0,107,0,0,0,64,0,192,0,0,0,0,0,152,0,169,0,77,0,25,0,122,0,13,0,176,0,220,0,221,0,143,0,0,0,0,0,35,0,0,0,17,0,255,0,230,0,191,0,71,0,0,0,213,0,128,0,215,0,8,0,143,0,193,0,0,0,55,0,38,0,0,0,175,0,162,0,158,0,0,0,59,0,62,0,82,0,66,0,209,0,167,0,26,0,61,0,20,0,252,0,131,0,83,0,153,0,221,0,0,0,240,0,42,0,0,0,232,0,75,0,0,0,138,0,0,0,187,0,129,0,218,0,114,0,219,0,255,0,0,0,234,0,49,0,0,0,0,0,12,0,108,0,105,0,0,0,160,0,51,0,207,0,42,0,127,0,246,0,92,0,0,0,0,0,72,0,107,0,255,0,78,0,118,0,30,0,0,0,146,0,200,0,114,0,0,0,0,0,144,0,162,0,3,0,45,0,207,0,0,0,9,0,0,0,173,0,159,0,101,0,55,0,188,0,127,0,176,0,51,0,89,0,42,0,116,0,52,0,161,0,124,0,148,0,19,0,2,0,188,0,0,0,0,0,0,0,0,0,0,0,0,0,173,0,60,0,224,0,0,0,193,0,226,0,99,0,186,0,221,0,10,0,100,0,25,0,26,0,144,0,180,0,112,0,5,0,88,0,0,0,16,0,89,0,0,0,247,0,132,0,248,0,90,0,101,0,0,0,34,0,141,0,181,0,152,0,183,0,163,0,89,0,195,0,49,0,5,0,203,0,89,0,156,0,122,0,223,0,0,0,45,0,70,0,82,0,10,0,226,0,130,0,117,0,151,0,0,0,77,0,57,0,162,0,198,0,13,0,69,0,110,0,85,0,0,0,51,0,22,0,30,0,212,0,141,0,178,0,0,0,206,0,170,0,113,0,220,0,0,0,0,0,103,0,67,0,242,0,4,0,6,0,63,0,0,0,184,0,251,0,225,0,23,0,194,0,227,0,0,0,0,0,0,0,155,0,77,0,146,0,109,0,16,0,92,0,0,0,195,0,125,0,234,0,176,0,0,0,179,0,0,0,31,0,83,0,0,0,233,0,210,0,61,0,0,0,189,0,0,0,244,0,213,0,240,0,76,0,0,0,170,0,164,0,0,0,0,0,0,0,31,0,28,0,0,0,92,0,0,0,214,0,24,0,227,0,185,0,248,0,77,0,37,0,109,0,0,0,73,0,169,0,169,0,42,0,11,0,5,0,122,0,251,0,208,0,0,0,188,0,135,0,136,0,7,0,77,0,0,0,189,0,213,0,247,0,132,0,29,0,19,0,240,0,83,0,0,0,0,0,23,0,110,0,63,0,0,0,59,0,59,0,164,0,244,0,110,0,8,0,159,0,0,0,0,0,243,0,97,0,199,0,128,0,0,0,218,0,69,0,0,0,222,0,0,0,222,0,21,0,0,0,44,0,247,0,34,0,220,0,23,0,0,0,13,0,240,0,117,0,0,0,12,0,0,0,78,0,80,0,55,0,138,0,230,0,13,0,60,0,127,0,80,0,114,0,53,0,144,0,142,0,48,0,86,0,182,0,111,0,252,0,0,0,221,0,101,0,190,0,0,0,0,0,0,0,0,0,160,0,0,0,110,0,158,0,234,0,89,0);
signal scenario_full  : scenario_type := (60,31,4,31,170,31,90,31,159,31,159,30,198,31,198,30,198,29,198,28,185,31,221,31,75,31,216,31,48,31,35,31,240,31,227,31,144,31,144,30,211,31,195,31,155,31,155,30,155,29,87,31,79,31,150,31,124,31,33,31,57,31,57,30,85,31,85,30,85,29,101,31,65,31,65,30,157,31,147,31,237,31,237,30,194,31,194,30,118,31,151,31,188,31,236,31,14,31,89,31,89,30,54,31,238,31,214,31,215,31,215,30,215,29,193,31,148,31,148,30,172,31,109,31,2,31,2,30,63,31,63,30,23,31,48,31,147,31,124,31,124,30,2,31,204,31,71,31,71,30,17,31,127,31,133,31,4,31,179,31,178,31,178,30,4,31,215,31,215,30,153,31,138,31,138,30,195,31,91,31,91,30,115,31,115,30,115,29,45,31,45,30,85,31,243,31,243,30,143,31,227,31,162,31,239,31,239,30,51,31,51,30,51,29,51,28,136,31,64,31,100,31,25,31,235,31,66,31,66,30,66,29,130,31,137,31,39,31,57,31,57,30,180,31,180,30,185,31,185,30,38,31,2,31,237,31,155,31,169,31,206,31,206,30,23,31,56,31,202,31,202,30,112,31,112,30,19,31,166,31,185,31,119,31,102,31,247,31,65,31,8,31,160,31,92,31,160,31,58,31,58,30,58,29,46,31,151,31,93,31,2,31,2,30,174,31,174,30,207,31,171,31,37,31,45,31,162,31,117,31,47,31,47,30,96,31,25,31,38,31,38,30,252,31,36,31,139,31,139,30,179,31,179,30,192,31,8,31,56,31,235,31,200,31,237,31,62,31,160,31,3,31,218,31,65,31,99,31,189,31,55,31,80,31,14,31,74,31,140,31,204,31,204,30,59,31,59,30,167,31,146,31,68,31,194,31,158,31,60,31,112,31,164,31,172,31,116,31,124,31,124,30,51,31,60,31,242,31,157,31,245,31,183,31,183,30,183,29,31,31,219,31,187,31,187,30,229,31,15,31,15,30,15,29,223,31,221,31,244,31,204,31,227,31,227,30,142,31,20,31,20,30,20,29,92,31,243,31,197,31,252,31,252,30,19,31,19,30,59,31,229,31,171,31,36,31,36,30,226,31,26,31,95,31,44,31,44,30,106,31,106,30,57,31,57,30,184,31,129,31,218,31,75,31,75,30,176,31,176,30,108,31,187,31,170,31,75,31,58,31,227,31,18,31,18,30,205,31,109,31,77,31,45,31,93,31,29,31,176,31,124,31,56,31,38,31,166,31,189,31,189,30,189,29,9,31,36,31,36,30,36,29,36,28,36,27,36,26,49,31,207,31,208,31,51,31,163,31,18,31,31,31,149,31,102,31,39,31,72,31,37,31,220,31,112,31,64,31,148,31,6,31,238,31,159,31,197,31,228,31,118,31,210,31,124,31,124,30,99,31,68,31,243,31,132,31,229,31,229,30,77,31,77,30,77,29,203,31,58,31,102,31,201,31,24,31,129,31,15,31,47,31,47,30,118,31,123,31,47,31,180,31,151,31,37,31,37,30,242,31,13,31,76,31,213,31,113,31,174,31,198,31,195,31,113,31,213,31,213,30,172,31,31,31,223,31,126,31,110,31,131,31,73,31,103,31,123,31,123,30,87,31,99,31,40,31,98,31,248,31,248,31,248,30,69,31,83,31,83,30,58,31,58,30,95,31,237,31,194,31,136,31,236,31,157,31,248,31,190,31,72,31,234,31,216,31,216,30,216,29,142,31,115,31,115,30,115,29,255,31,255,30,255,29,149,31,142,31,142,30,239,31,239,30,23,31,42,31,42,30,246,31,115,31,193,31,122,31,187,31,126,31,126,30,147,31,51,31,219,31,219,30,64,31,255,31,255,30,29,31,144,31,196,31,196,30,68,31,67,31,12,31,151,31,163,31,239,31,169,31,32,31,246,31,246,30,110,31,176,31,16,31,134,31,233,31,95,31,61,31,32,31,104,31,1,31,98,31,10,31,255,31,249,31,68,31,45,31,180,31,3,31,3,30,129,31,89,31,139,31,14,31,14,30,192,31,241,31,241,30,241,29,92,31,92,30,105,31,107,31,80,31,80,30,97,31,97,30,222,31,222,30,94,31,162,31,107,31,107,30,64,31,192,31,192,30,192,29,152,31,169,31,77,31,25,31,122,31,13,31,176,31,220,31,221,31,143,31,143,30,143,29,35,31,35,30,17,31,255,31,230,31,191,31,71,31,71,30,213,31,128,31,215,31,8,31,143,31,193,31,193,30,55,31,38,31,38,30,175,31,162,31,158,31,158,30,59,31,62,31,82,31,66,31,209,31,167,31,26,31,61,31,20,31,252,31,131,31,83,31,153,31,221,31,221,30,240,31,42,31,42,30,232,31,75,31,75,30,138,31,138,30,187,31,129,31,218,31,114,31,219,31,255,31,255,30,234,31,49,31,49,30,49,29,12,31,108,31,105,31,105,30,160,31,51,31,207,31,42,31,127,31,246,31,92,31,92,30,92,29,72,31,107,31,255,31,78,31,118,31,30,31,30,30,146,31,200,31,114,31,114,30,114,29,144,31,162,31,3,31,45,31,207,31,207,30,9,31,9,30,173,31,159,31,101,31,55,31,188,31,127,31,176,31,51,31,89,31,42,31,116,31,52,31,161,31,124,31,148,31,19,31,2,31,188,31,188,30,188,29,188,28,188,27,188,26,188,25,173,31,60,31,224,31,224,30,193,31,226,31,99,31,186,31,221,31,10,31,100,31,25,31,26,31,144,31,180,31,112,31,5,31,88,31,88,30,16,31,89,31,89,30,247,31,132,31,248,31,90,31,101,31,101,30,34,31,141,31,181,31,152,31,183,31,163,31,89,31,195,31,49,31,5,31,203,31,89,31,156,31,122,31,223,31,223,30,45,31,70,31,82,31,10,31,226,31,130,31,117,31,151,31,151,30,77,31,57,31,162,31,198,31,13,31,69,31,110,31,85,31,85,30,51,31,22,31,30,31,212,31,141,31,178,31,178,30,206,31,170,31,113,31,220,31,220,30,220,29,103,31,67,31,242,31,4,31,6,31,63,31,63,30,184,31,251,31,225,31,23,31,194,31,227,31,227,30,227,29,227,28,155,31,77,31,146,31,109,31,16,31,92,31,92,30,195,31,125,31,234,31,176,31,176,30,179,31,179,30,31,31,83,31,83,30,233,31,210,31,61,31,61,30,189,31,189,30,244,31,213,31,240,31,76,31,76,30,170,31,164,31,164,30,164,29,164,28,31,31,28,31,28,30,92,31,92,30,214,31,24,31,227,31,185,31,248,31,77,31,37,31,109,31,109,30,73,31,169,31,169,31,42,31,11,31,5,31,122,31,251,31,208,31,208,30,188,31,135,31,136,31,7,31,77,31,77,30,189,31,213,31,247,31,132,31,29,31,19,31,240,31,83,31,83,30,83,29,23,31,110,31,63,31,63,30,59,31,59,31,164,31,244,31,110,31,8,31,159,31,159,30,159,29,243,31,97,31,199,31,128,31,128,30,218,31,69,31,69,30,222,31,222,30,222,31,21,31,21,30,44,31,247,31,34,31,220,31,23,31,23,30,13,31,240,31,117,31,117,30,12,31,12,30,78,31,80,31,55,31,138,31,230,31,13,31,60,31,127,31,80,31,114,31,53,31,144,31,142,31,48,31,86,31,182,31,111,31,252,31,252,30,221,31,101,31,190,31,190,30,190,29,190,28,190,27,160,31,160,30,110,31,158,31,234,31,89,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
