-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 726;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (224,0,187,0,154,0,143,0,122,0,214,0,163,0,0,0,115,0,0,0,0,0,233,0,141,0,125,0,0,0,80,0,82,0,0,0,84,0,7,0,0,0,51,0,178,0,0,0,0,0,62,0,147,0,0,0,110,0,0,0,151,0,0,0,137,0,216,0,104,0,197,0,87,0,172,0,163,0,236,0,80,0,0,0,248,0,17,0,113,0,83,0,124,0,35,0,128,0,6,0,194,0,195,0,0,0,162,0,52,0,198,0,11,0,42,0,194,0,176,0,241,0,74,0,111,0,39,0,29,0,0,0,27,0,223,0,30,0,33,0,193,0,174,0,0,0,122,0,0,0,193,0,42,0,0,0,0,0,106,0,5,0,67,0,205,0,49,0,91,0,181,0,79,0,0,0,149,0,132,0,71,0,110,0,228,0,124,0,135,0,205,0,14,0,236,0,174,0,55,0,4,0,0,0,63,0,7,0,142,0,172,0,182,0,117,0,0,0,249,0,43,0,253,0,35,0,123,0,81,0,161,0,199,0,37,0,0,0,0,0,185,0,0,0,0,0,176,0,86,0,140,0,218,0,22,0,72,0,210,0,89,0,137,0,182,0,148,0,135,0,198,0,110,0,216,0,198,0,22,0,94,0,124,0,52,0,0,0,226,0,1,0,105,0,252,0,159,0,153,0,0,0,0,0,0,0,9,0,95,0,37,0,188,0,190,0,1,0,0,0,16,0,52,0,232,0,26,0,0,0,90,0,115,0,0,0,0,0,247,0,0,0,187,0,67,0,180,0,228,0,0,0,2,0,33,0,235,0,20,0,158,0,157,0,160,0,96,0,81,0,219,0,0,0,235,0,0,0,96,0,100,0,236,0,247,0,77,0,104,0,248,0,0,0,157,0,181,0,44,0,169,0,236,0,0,0,0,0,59,0,73,0,110,0,159,0,0,0,102,0,95,0,227,0,0,0,58,0,0,0,0,0,254,0,255,0,28,0,208,0,107,0,0,0,179,0,0,0,0,0,129,0,0,0,163,0,0,0,40,0,0,0,213,0,11,0,117,0,160,0,167,0,91,0,164,0,115,0,63,0,166,0,86,0,181,0,172,0,192,0,40,0,206,0,0,0,0,0,0,0,76,0,233,0,6,0,190,0,0,0,19,0,39,0,245,0,134,0,27,0,0,0,147,0,2,0,112,0,40,0,153,0,0,0,215,0,74,0,34,0,47,0,0,0,75,0,90,0,186,0,221,0,9,0,0,0,183,0,227,0,113,0,49,0,166,0,99,0,61,0,198,0,0,0,0,0,223,0,168,0,0,0,223,0,0,0,74,0,129,0,160,0,98,0,64,0,89,0,173,0,128,0,0,0,66,0,107,0,167,0,193,0,46,0,15,0,176,0,89,0,195,0,173,0,218,0,37,0,65,0,51,0,102,0,4,0,0,0,15,0,25,0,228,0,0,0,28,0,21,0,125,0,114,0,191,0,8,0,194,0,73,0,128,0,170,0,9,0,41,0,115,0,91,0,187,0,203,0,111,0,0,0,31,0,82,0,73,0,244,0,104,0,0,0,7,0,0,0,225,0,169,0,6,0,0,0,201,0,0,0,41,0,201,0,42,0,37,0,189,0,124,0,195,0,64,0,0,0,0,0,41,0,48,0,0,0,0,0,230,0,209,0,0,0,186,0,0,0,0,0,0,0,209,0,140,0,3,0,177,0,0,0,121,0,22,0,144,0,44,0,0,0,0,0,196,0,216,0,214,0,40,0,62,0,165,0,88,0,33,0,164,0,118,0,11,0,135,0,158,0,0,0,166,0,239,0,134,0,97,0,0,0,96,0,0,0,208,0,213,0,175,0,212,0,105,0,15,0,0,0,183,0,0,0,108,0,0,0,208,0,0,0,158,0,208,0,34,0,0,0,212,0,138,0,109,0,0,0,69,0,134,0,245,0,144,0,198,0,207,0,120,0,0,0,7,0,202,0,0,0,148,0,214,0,225,0,35,0,13,0,0,0,0,0,199,0,71,0,97,0,32,0,161,0,18,0,41,0,207,0,190,0,0,0,162,0,250,0,174,0,188,0,36,0,14,0,232,0,195,0,246,0,184,0,136,0,43,0,60,0,246,0,29,0,23,0,57,0,148,0,9,0,145,0,19,0,0,0,36,0,219,0,0,0,153,0,208,0,0,0,179,0,148,0,0,0,30,0,0,0,245,0,0,0,71,0,253,0,118,0,5,0,102,0,0,0,135,0,43,0,217,0,0,0,137,0,11,0,127,0,61,0,70,0,0,0,119,0,90,0,78,0,239,0,0,0,185,0,233,0,0,0,215,0,249,0,14,0,45,0,0,0,131,0,0,0,28,0,0,0,32,0,133,0,142,0,44,0,158,0,69,0,5,0,0,0,113,0,190,0,138,0,95,0,13,0,193,0,168,0,0,0,173,0,119,0,106,0,113,0,212,0,255,0,103,0,158,0,121,0,0,0,76,0,112,0,142,0,0,0,166,0,0,0,0,0,155,0,19,0,39,0,67,0,226,0,185,0,78,0,125,0,95,0,26,0,216,0,4,0,0,0,83,0,44,0,217,0,163,0,19,0,28,0,51,0,92,0,0,0,70,0,69,0,56,0,122,0,31,0,50,0,219,0,80,0,0,0,60,0,101,0,0,0,152,0,146,0,69,0,222,0,48,0,146,0,18,0,35,0,207,0,0,0,143,0,71,0,50,0,60,0,37,0,8,0,0,0,40,0,107,0,0,0,0,0,229,0,242,0,0,0,126,0,48,0,83,0,173,0,223,0,0,0,170,0,141,0,60,0,99,0,145,0,11,0,107,0,116,0,107,0,69,0,118,0,0,0,0,0,7,0,55,0,106,0,19,0,64,0,0,0,79,0,0,0,47,0,127,0,86,0,174,0,132,0,230,0,0,0,0,0,44,0,10,0,119,0,233,0,0,0,165,0,154,0,0,0,86,0,36,0,55,0,32,0,23,0,164,0,81,0,153,0,42,0,0,0,237,0,201,0,216,0,0,0,235,0,179,0,34,0,236,0,51,0,0,0,73,0,233,0,10,0,185,0,38,0,0,0,39,0,0,0,104,0,203,0,65,0,38,0,0,0,88,0,157,0,89,0,177,0,24,0,86,0,145,0,239,0,106,0,75,0,147,0,0,0,0,0,31,0,146,0,101,0,191,0,244,0,0,0,174,0,91,0,44,0,57,0,236,0,125,0,148,0,60,0,0,0,0,0,0,0,116,0,0,0,189,0,81,0);
signal scenario_full  : scenario_type := (224,31,187,31,154,31,143,31,122,31,214,31,163,31,163,30,115,31,115,30,115,29,233,31,141,31,125,31,125,30,80,31,82,31,82,30,84,31,7,31,7,30,51,31,178,31,178,30,178,29,62,31,147,31,147,30,110,31,110,30,151,31,151,30,137,31,216,31,104,31,197,31,87,31,172,31,163,31,236,31,80,31,80,30,248,31,17,31,113,31,83,31,124,31,35,31,128,31,6,31,194,31,195,31,195,30,162,31,52,31,198,31,11,31,42,31,194,31,176,31,241,31,74,31,111,31,39,31,29,31,29,30,27,31,223,31,30,31,33,31,193,31,174,31,174,30,122,31,122,30,193,31,42,31,42,30,42,29,106,31,5,31,67,31,205,31,49,31,91,31,181,31,79,31,79,30,149,31,132,31,71,31,110,31,228,31,124,31,135,31,205,31,14,31,236,31,174,31,55,31,4,31,4,30,63,31,7,31,142,31,172,31,182,31,117,31,117,30,249,31,43,31,253,31,35,31,123,31,81,31,161,31,199,31,37,31,37,30,37,29,185,31,185,30,185,29,176,31,86,31,140,31,218,31,22,31,72,31,210,31,89,31,137,31,182,31,148,31,135,31,198,31,110,31,216,31,198,31,22,31,94,31,124,31,52,31,52,30,226,31,1,31,105,31,252,31,159,31,153,31,153,30,153,29,153,28,9,31,95,31,37,31,188,31,190,31,1,31,1,30,16,31,52,31,232,31,26,31,26,30,90,31,115,31,115,30,115,29,247,31,247,30,187,31,67,31,180,31,228,31,228,30,2,31,33,31,235,31,20,31,158,31,157,31,160,31,96,31,81,31,219,31,219,30,235,31,235,30,96,31,100,31,236,31,247,31,77,31,104,31,248,31,248,30,157,31,181,31,44,31,169,31,236,31,236,30,236,29,59,31,73,31,110,31,159,31,159,30,102,31,95,31,227,31,227,30,58,31,58,30,58,29,254,31,255,31,28,31,208,31,107,31,107,30,179,31,179,30,179,29,129,31,129,30,163,31,163,30,40,31,40,30,213,31,11,31,117,31,160,31,167,31,91,31,164,31,115,31,63,31,166,31,86,31,181,31,172,31,192,31,40,31,206,31,206,30,206,29,206,28,76,31,233,31,6,31,190,31,190,30,19,31,39,31,245,31,134,31,27,31,27,30,147,31,2,31,112,31,40,31,153,31,153,30,215,31,74,31,34,31,47,31,47,30,75,31,90,31,186,31,221,31,9,31,9,30,183,31,227,31,113,31,49,31,166,31,99,31,61,31,198,31,198,30,198,29,223,31,168,31,168,30,223,31,223,30,74,31,129,31,160,31,98,31,64,31,89,31,173,31,128,31,128,30,66,31,107,31,167,31,193,31,46,31,15,31,176,31,89,31,195,31,173,31,218,31,37,31,65,31,51,31,102,31,4,31,4,30,15,31,25,31,228,31,228,30,28,31,21,31,125,31,114,31,191,31,8,31,194,31,73,31,128,31,170,31,9,31,41,31,115,31,91,31,187,31,203,31,111,31,111,30,31,31,82,31,73,31,244,31,104,31,104,30,7,31,7,30,225,31,169,31,6,31,6,30,201,31,201,30,41,31,201,31,42,31,37,31,189,31,124,31,195,31,64,31,64,30,64,29,41,31,48,31,48,30,48,29,230,31,209,31,209,30,186,31,186,30,186,29,186,28,209,31,140,31,3,31,177,31,177,30,121,31,22,31,144,31,44,31,44,30,44,29,196,31,216,31,214,31,40,31,62,31,165,31,88,31,33,31,164,31,118,31,11,31,135,31,158,31,158,30,166,31,239,31,134,31,97,31,97,30,96,31,96,30,208,31,213,31,175,31,212,31,105,31,15,31,15,30,183,31,183,30,108,31,108,30,208,31,208,30,158,31,208,31,34,31,34,30,212,31,138,31,109,31,109,30,69,31,134,31,245,31,144,31,198,31,207,31,120,31,120,30,7,31,202,31,202,30,148,31,214,31,225,31,35,31,13,31,13,30,13,29,199,31,71,31,97,31,32,31,161,31,18,31,41,31,207,31,190,31,190,30,162,31,250,31,174,31,188,31,36,31,14,31,232,31,195,31,246,31,184,31,136,31,43,31,60,31,246,31,29,31,23,31,57,31,148,31,9,31,145,31,19,31,19,30,36,31,219,31,219,30,153,31,208,31,208,30,179,31,148,31,148,30,30,31,30,30,245,31,245,30,71,31,253,31,118,31,5,31,102,31,102,30,135,31,43,31,217,31,217,30,137,31,11,31,127,31,61,31,70,31,70,30,119,31,90,31,78,31,239,31,239,30,185,31,233,31,233,30,215,31,249,31,14,31,45,31,45,30,131,31,131,30,28,31,28,30,32,31,133,31,142,31,44,31,158,31,69,31,5,31,5,30,113,31,190,31,138,31,95,31,13,31,193,31,168,31,168,30,173,31,119,31,106,31,113,31,212,31,255,31,103,31,158,31,121,31,121,30,76,31,112,31,142,31,142,30,166,31,166,30,166,29,155,31,19,31,39,31,67,31,226,31,185,31,78,31,125,31,95,31,26,31,216,31,4,31,4,30,83,31,44,31,217,31,163,31,19,31,28,31,51,31,92,31,92,30,70,31,69,31,56,31,122,31,31,31,50,31,219,31,80,31,80,30,60,31,101,31,101,30,152,31,146,31,69,31,222,31,48,31,146,31,18,31,35,31,207,31,207,30,143,31,71,31,50,31,60,31,37,31,8,31,8,30,40,31,107,31,107,30,107,29,229,31,242,31,242,30,126,31,48,31,83,31,173,31,223,31,223,30,170,31,141,31,60,31,99,31,145,31,11,31,107,31,116,31,107,31,69,31,118,31,118,30,118,29,7,31,55,31,106,31,19,31,64,31,64,30,79,31,79,30,47,31,127,31,86,31,174,31,132,31,230,31,230,30,230,29,44,31,10,31,119,31,233,31,233,30,165,31,154,31,154,30,86,31,36,31,55,31,32,31,23,31,164,31,81,31,153,31,42,31,42,30,237,31,201,31,216,31,216,30,235,31,179,31,34,31,236,31,51,31,51,30,73,31,233,31,10,31,185,31,38,31,38,30,39,31,39,30,104,31,203,31,65,31,38,31,38,30,88,31,157,31,89,31,177,31,24,31,86,31,145,31,239,31,106,31,75,31,147,31,147,30,147,29,31,31,146,31,101,31,191,31,244,31,244,30,174,31,91,31,44,31,57,31,236,31,125,31,148,31,60,31,60,30,60,29,60,28,116,31,116,30,189,31,81,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
