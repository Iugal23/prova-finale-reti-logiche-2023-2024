-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_504 is
end project_tb_504;

architecture project_tb_arch_504 of project_tb_504 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 843;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (215,0,39,0,141,0,241,0,0,0,193,0,194,0,146,0,0,0,53,0,124,0,209,0,219,0,229,0,102,0,0,0,120,0,54,0,236,0,20,0,132,0,13,0,240,0,162,0,0,0,159,0,106,0,0,0,84,0,0,0,27,0,182,0,207,0,0,0,232,0,45,0,218,0,54,0,219,0,0,0,79,0,0,0,145,0,104,0,14,0,79,0,249,0,179,0,0,0,97,0,0,0,105,0,145,0,255,0,186,0,220,0,176,0,122,0,192,0,128,0,0,0,254,0,100,0,93,0,153,0,0,0,113,0,12,0,0,0,174,0,191,0,96,0,89,0,0,0,0,0,188,0,187,0,43,0,50,0,0,0,0,0,245,0,25,0,109,0,0,0,0,0,147,0,26,0,38,0,32,0,0,0,0,0,151,0,0,0,2,0,25,0,104,0,29,0,42,0,0,0,26,0,40,0,122,0,67,0,226,0,212,0,154,0,119,0,0,0,47,0,47,0,0,0,223,0,64,0,210,0,0,0,140,0,58,0,46,0,78,0,17,0,249,0,34,0,156,0,0,0,159,0,84,0,176,0,81,0,169,0,221,0,98,0,69,0,105,0,118,0,186,0,58,0,200,0,109,0,0,0,19,0,0,0,0,0,207,0,169,0,243,0,0,0,165,0,222,0,239,0,0,0,5,0,241,0,34,0,233,0,178,0,0,0,32,0,100,0,0,0,91,0,0,0,0,0,15,0,183,0,177,0,139,0,221,0,98,0,143,0,201,0,0,0,240,0,234,0,0,0,208,0,116,0,67,0,232,0,19,0,82,0,161,0,148,0,5,0,33,0,50,0,26,0,190,0,0,0,23,0,7,0,136,0,239,0,46,0,87,0,208,0,49,0,0,0,143,0,86,0,36,0,122,0,0,0,5,0,211,0,0,0,36,0,0,0,71,0,85,0,148,0,116,0,211,0,138,0,200,0,219,0,53,0,237,0,140,0,160,0,0,0,28,0,97,0,168,0,235,0,207,0,0,0,0,0,155,0,0,0,194,0,212,0,185,0,61,0,74,0,0,0,56,0,0,0,0,0,247,0,198,0,205,0,7,0,0,0,236,0,0,0,204,0,25,0,123,0,29,0,170,0,244,0,0,0,0,0,156,0,0,0,93,0,0,0,0,0,0,0,223,0,69,0,139,0,114,0,251,0,180,0,62,0,33,0,100,0,143,0,191,0,0,0,199,0,186,0,116,0,230,0,92,0,242,0,199,0,156,0,0,0,89,0,0,0,221,0,0,0,0,0,0,0,210,0,118,0,215,0,50,0,0,0,150,0,35,0,187,0,0,0,0,0,0,0,0,0,0,0,214,0,111,0,212,0,43,0,168,0,222,0,186,0,153,0,59,0,174,0,86,0,160,0,47,0,96,0,255,0,0,0,137,0,61,0,64,0,209,0,0,0,53,0,173,0,27,0,77,0,205,0,88,0,23,0,4,0,49,0,206,0,25,0,42,0,0,0,51,0,114,0,156,0,94,0,177,0,49,0,172,0,202,0,191,0,98,0,54,0,207,0,48,0,146,0,179,0,0,0,187,0,116,0,134,0,0,0,40,0,190,0,210,0,0,0,99,0,0,0,97,0,0,0,4,0,189,0,230,0,252,0,14,0,34,0,211,0,97,0,205,0,103,0,130,0,224,0,71,0,110,0,245,0,139,0,161,0,234,0,79,0,0,0,6,0,62,0,42,0,0,0,181,0,107,0,134,0,108,0,156,0,246,0,0,0,170,0,0,0,0,0,188,0,0,0,235,0,199,0,165,0,156,0,85,0,236,0,0,0,109,0,137,0,231,0,106,0,3,0,221,0,0,0,62,0,205,0,144,0,215,0,110,0,212,0,71,0,182,0,212,0,161,0,71,0,250,0,51,0,35,0,19,0,249,0,42,0,0,0,143,0,95,0,192,0,47,0,174,0,236,0,0,0,160,0,0,0,120,0,235,0,150,0,0,0,181,0,0,0,191,0,75,0,213,0,182,0,95,0,204,0,197,0,170,0,45,0,86,0,161,0,192,0,246,0,164,0,0,0,61,0,0,0,236,0,114,0,217,0,86,0,17,0,35,0,220,0,55,0,63,0,90,0,154,0,162,0,177,0,86,0,105,0,0,0,0,0,18,0,190,0,95,0,29,0,97,0,195,0,152,0,153,0,65,0,0,0,0,0,161,0,61,0,212,0,214,0,0,0,199,0,246,0,98,0,32,0,0,0,58,0,65,0,127,0,192,0,193,0,184,0,0,0,47,0,0,0,141,0,110,0,0,0,0,0,0,0,232,0,72,0,0,0,51,0,153,0,231,0,158,0,0,0,161,0,45,0,237,0,42,0,169,0,157,0,250,0,25,0,226,0,57,0,120,0,80,0,241,0,140,0,115,0,46,0,124,0,0,0,40,0,92,0,0,0,171,0,209,0,121,0,99,0,158,0,121,0,136,0,0,0,65,0,59,0,37,0,0,0,72,0,72,0,128,0,135,0,0,0,116,0,180,0,0,0,110,0,210,0,113,0,49,0,0,0,166,0,4,0,228,0,47,0,42,0,234,0,194,0,168,0,0,0,250,0,0,0,0,0,128,0,221,0,47,0,148,0,0,0,178,0,0,0,68,0,120,0,0,0,139,0,194,0,141,0,149,0,19,0,6,0,224,0,199,0,138,0,0,0,51,0,0,0,0,0,251,0,129,0,47,0,4,0,29,0,110,0,11,0,183,0,217,0,73,0,27,0,11,0,191,0,0,0,7,0,198,0,83,0,192,0,0,0,0,0,0,0,124,0,172,0,123,0,0,0,148,0,176,0,25,0,214,0,43,0,138,0,0,0,244,0,25,0,0,0,202,0,243,0,0,0,0,0,178,0,0,0,0,0,154,0,115,0,100,0,41,0,80,0,199,0,243,0,0,0,132,0,46,0,214,0,29,0,223,0,57,0,250,0,92,0,148,0,163,0,147,0,182,0,31,0,0,0,0,0,0,0,0,0,194,0,215,0,138,0,202,0,118,0,0,0,112,0,49,0,228,0,120,0,195,0,68,0,0,0,72,0,0,0,103,0,180,0,62,0,188,0,238,0,214,0,109,0,160,0,209,0,97,0,226,0,0,0,151,0,130,0,136,0,218,0,0,0,0,0,82,0,23,0,0,0,154,0,0,0,253,0,189,0,154,0,235,0,131,0,8,0,182,0,0,0,208,0,93,0,212,0,180,0,226,0,179,0,255,0,0,0,47,0,0,0,185,0,17,0,0,0,228,0,142,0,133,0,232,0,193,0,53,0,19,0,27,0,0,0,219,0,154,0,0,0,64,0,184,0,194,0,51,0,209,0,146,0,34,0,0,0,46,0,16,0,185,0,201,0,190,0,211,0,123,0,181,0,242,0,241,0,0,0,75,0,186,0,0,0,0,0,224,0,98,0,197,0,107,0,46,0,107,0,0,0,74,0,71,0,0,0,131,0,16,0,0,0,0,0,0,0,43,0,200,0,173,0,39,0,142,0,132,0,0,0,0,0,0,0,239,0,170,0,209,0,147,0,0,0,0,0,40,0,87,0,206,0,218,0,149,0,0,0,235,0,0,0,0,0,8,0,82,0,39,0,49,0,122,0,0,0,139,0,156,0,0,0,249,0,100,0,247,0,69,0,97,0,201,0,0,0,197,0,10,0,7,0,193,0,61,0,72,0,79,0,112,0,124,0,255,0,80,0,248,0,41,0,110,0,10,0,229,0,1,0,0,0,0,0,0,0,0,0,87,0,0,0,121,0);
signal scenario_full  : scenario_type := (215,31,39,31,141,31,241,31,241,30,193,31,194,31,146,31,146,30,53,31,124,31,209,31,219,31,229,31,102,31,102,30,120,31,54,31,236,31,20,31,132,31,13,31,240,31,162,31,162,30,159,31,106,31,106,30,84,31,84,30,27,31,182,31,207,31,207,30,232,31,45,31,218,31,54,31,219,31,219,30,79,31,79,30,145,31,104,31,14,31,79,31,249,31,179,31,179,30,97,31,97,30,105,31,145,31,255,31,186,31,220,31,176,31,122,31,192,31,128,31,128,30,254,31,100,31,93,31,153,31,153,30,113,31,12,31,12,30,174,31,191,31,96,31,89,31,89,30,89,29,188,31,187,31,43,31,50,31,50,30,50,29,245,31,25,31,109,31,109,30,109,29,147,31,26,31,38,31,32,31,32,30,32,29,151,31,151,30,2,31,25,31,104,31,29,31,42,31,42,30,26,31,40,31,122,31,67,31,226,31,212,31,154,31,119,31,119,30,47,31,47,31,47,30,223,31,64,31,210,31,210,30,140,31,58,31,46,31,78,31,17,31,249,31,34,31,156,31,156,30,159,31,84,31,176,31,81,31,169,31,221,31,98,31,69,31,105,31,118,31,186,31,58,31,200,31,109,31,109,30,19,31,19,30,19,29,207,31,169,31,243,31,243,30,165,31,222,31,239,31,239,30,5,31,241,31,34,31,233,31,178,31,178,30,32,31,100,31,100,30,91,31,91,30,91,29,15,31,183,31,177,31,139,31,221,31,98,31,143,31,201,31,201,30,240,31,234,31,234,30,208,31,116,31,67,31,232,31,19,31,82,31,161,31,148,31,5,31,33,31,50,31,26,31,190,31,190,30,23,31,7,31,136,31,239,31,46,31,87,31,208,31,49,31,49,30,143,31,86,31,36,31,122,31,122,30,5,31,211,31,211,30,36,31,36,30,71,31,85,31,148,31,116,31,211,31,138,31,200,31,219,31,53,31,237,31,140,31,160,31,160,30,28,31,97,31,168,31,235,31,207,31,207,30,207,29,155,31,155,30,194,31,212,31,185,31,61,31,74,31,74,30,56,31,56,30,56,29,247,31,198,31,205,31,7,31,7,30,236,31,236,30,204,31,25,31,123,31,29,31,170,31,244,31,244,30,244,29,156,31,156,30,93,31,93,30,93,29,93,28,223,31,69,31,139,31,114,31,251,31,180,31,62,31,33,31,100,31,143,31,191,31,191,30,199,31,186,31,116,31,230,31,92,31,242,31,199,31,156,31,156,30,89,31,89,30,221,31,221,30,221,29,221,28,210,31,118,31,215,31,50,31,50,30,150,31,35,31,187,31,187,30,187,29,187,28,187,27,187,26,214,31,111,31,212,31,43,31,168,31,222,31,186,31,153,31,59,31,174,31,86,31,160,31,47,31,96,31,255,31,255,30,137,31,61,31,64,31,209,31,209,30,53,31,173,31,27,31,77,31,205,31,88,31,23,31,4,31,49,31,206,31,25,31,42,31,42,30,51,31,114,31,156,31,94,31,177,31,49,31,172,31,202,31,191,31,98,31,54,31,207,31,48,31,146,31,179,31,179,30,187,31,116,31,134,31,134,30,40,31,190,31,210,31,210,30,99,31,99,30,97,31,97,30,4,31,189,31,230,31,252,31,14,31,34,31,211,31,97,31,205,31,103,31,130,31,224,31,71,31,110,31,245,31,139,31,161,31,234,31,79,31,79,30,6,31,62,31,42,31,42,30,181,31,107,31,134,31,108,31,156,31,246,31,246,30,170,31,170,30,170,29,188,31,188,30,235,31,199,31,165,31,156,31,85,31,236,31,236,30,109,31,137,31,231,31,106,31,3,31,221,31,221,30,62,31,205,31,144,31,215,31,110,31,212,31,71,31,182,31,212,31,161,31,71,31,250,31,51,31,35,31,19,31,249,31,42,31,42,30,143,31,95,31,192,31,47,31,174,31,236,31,236,30,160,31,160,30,120,31,235,31,150,31,150,30,181,31,181,30,191,31,75,31,213,31,182,31,95,31,204,31,197,31,170,31,45,31,86,31,161,31,192,31,246,31,164,31,164,30,61,31,61,30,236,31,114,31,217,31,86,31,17,31,35,31,220,31,55,31,63,31,90,31,154,31,162,31,177,31,86,31,105,31,105,30,105,29,18,31,190,31,95,31,29,31,97,31,195,31,152,31,153,31,65,31,65,30,65,29,161,31,61,31,212,31,214,31,214,30,199,31,246,31,98,31,32,31,32,30,58,31,65,31,127,31,192,31,193,31,184,31,184,30,47,31,47,30,141,31,110,31,110,30,110,29,110,28,232,31,72,31,72,30,51,31,153,31,231,31,158,31,158,30,161,31,45,31,237,31,42,31,169,31,157,31,250,31,25,31,226,31,57,31,120,31,80,31,241,31,140,31,115,31,46,31,124,31,124,30,40,31,92,31,92,30,171,31,209,31,121,31,99,31,158,31,121,31,136,31,136,30,65,31,59,31,37,31,37,30,72,31,72,31,128,31,135,31,135,30,116,31,180,31,180,30,110,31,210,31,113,31,49,31,49,30,166,31,4,31,228,31,47,31,42,31,234,31,194,31,168,31,168,30,250,31,250,30,250,29,128,31,221,31,47,31,148,31,148,30,178,31,178,30,68,31,120,31,120,30,139,31,194,31,141,31,149,31,19,31,6,31,224,31,199,31,138,31,138,30,51,31,51,30,51,29,251,31,129,31,47,31,4,31,29,31,110,31,11,31,183,31,217,31,73,31,27,31,11,31,191,31,191,30,7,31,198,31,83,31,192,31,192,30,192,29,192,28,124,31,172,31,123,31,123,30,148,31,176,31,25,31,214,31,43,31,138,31,138,30,244,31,25,31,25,30,202,31,243,31,243,30,243,29,178,31,178,30,178,29,154,31,115,31,100,31,41,31,80,31,199,31,243,31,243,30,132,31,46,31,214,31,29,31,223,31,57,31,250,31,92,31,148,31,163,31,147,31,182,31,31,31,31,30,31,29,31,28,31,27,194,31,215,31,138,31,202,31,118,31,118,30,112,31,49,31,228,31,120,31,195,31,68,31,68,30,72,31,72,30,103,31,180,31,62,31,188,31,238,31,214,31,109,31,160,31,209,31,97,31,226,31,226,30,151,31,130,31,136,31,218,31,218,30,218,29,82,31,23,31,23,30,154,31,154,30,253,31,189,31,154,31,235,31,131,31,8,31,182,31,182,30,208,31,93,31,212,31,180,31,226,31,179,31,255,31,255,30,47,31,47,30,185,31,17,31,17,30,228,31,142,31,133,31,232,31,193,31,53,31,19,31,27,31,27,30,219,31,154,31,154,30,64,31,184,31,194,31,51,31,209,31,146,31,34,31,34,30,46,31,16,31,185,31,201,31,190,31,211,31,123,31,181,31,242,31,241,31,241,30,75,31,186,31,186,30,186,29,224,31,98,31,197,31,107,31,46,31,107,31,107,30,74,31,71,31,71,30,131,31,16,31,16,30,16,29,16,28,43,31,200,31,173,31,39,31,142,31,132,31,132,30,132,29,132,28,239,31,170,31,209,31,147,31,147,30,147,29,40,31,87,31,206,31,218,31,149,31,149,30,235,31,235,30,235,29,8,31,82,31,39,31,49,31,122,31,122,30,139,31,156,31,156,30,249,31,100,31,247,31,69,31,97,31,201,31,201,30,197,31,10,31,7,31,193,31,61,31,72,31,79,31,112,31,124,31,255,31,80,31,248,31,41,31,110,31,10,31,229,31,1,31,1,30,1,29,1,28,1,27,87,31,87,30,121,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
