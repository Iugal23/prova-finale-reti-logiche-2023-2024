-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 746;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (134,0,166,0,88,0,0,0,173,0,50,0,132,0,246,0,52,0,125,0,0,0,192,0,0,0,0,0,64,0,0,0,70,0,153,0,204,0,199,0,0,0,0,0,25,0,185,0,83,0,84,0,193,0,0,0,0,0,65,0,90,0,42,0,85,0,227,0,99,0,235,0,225,0,251,0,53,0,251,0,204,0,139,0,248,0,252,0,235,0,42,0,95,0,196,0,240,0,34,0,42,0,229,0,245,0,250,0,17,0,156,0,128,0,57,0,74,0,255,0,168,0,171,0,95,0,0,0,251,0,206,0,0,0,170,0,0,0,0,0,0,0,112,0,200,0,66,0,237,0,0,0,29,0,41,0,55,0,146,0,218,0,117,0,69,0,0,0,167,0,104,0,48,0,30,0,0,0,0,0,32,0,185,0,0,0,0,0,11,0,133,0,0,0,130,0,25,0,25,0,205,0,142,0,0,0,22,0,56,0,113,0,13,0,31,0,222,0,17,0,162,0,35,0,225,0,99,0,140,0,168,0,151,0,57,0,16,0,0,0,0,0,43,0,83,0,114,0,217,0,166,0,209,0,0,0,183,0,245,0,243,0,0,0,225,0,61,0,243,0,0,0,0,0,116,0,0,0,104,0,89,0,85,0,9,0,67,0,225,0,0,0,158,0,0,0,0,0,143,0,0,0,204,0,13,0,173,0,241,0,0,0,106,0,220,0,0,0,0,0,53,0,70,0,0,0,0,0,0,0,237,0,101,0,250,0,0,0,78,0,212,0,94,0,0,0,153,0,91,0,41,0,63,0,181,0,24,0,61,0,186,0,228,0,26,0,0,0,249,0,63,0,205,0,243,0,142,0,252,0,175,0,149,0,127,0,60,0,91,0,126,0,0,0,188,0,209,0,200,0,113,0,245,0,0,0,156,0,178,0,0,0,234,0,187,0,0,0,1,0,112,0,82,0,182,0,173,0,179,0,155,0,152,0,17,0,169,0,241,0,166,0,30,0,191,0,70,0,177,0,102,0,219,0,210,0,83,0,224,0,129,0,140,0,51,0,80,0,182,0,0,0,88,0,132,0,65,0,40,0,0,0,22,0,197,0,159,0,124,0,28,0,164,0,91,0,14,0,94,0,0,0,205,0,0,0,204,0,96,0,98,0,148,0,0,0,7,0,39,0,156,0,81,0,59,0,212,0,248,0,106,0,82,0,47,0,168,0,186,0,111,0,112,0,185,0,194,0,200,0,135,0,0,0,164,0,214,0,0,0,0,0,195,0,0,0,146,0,44,0,134,0,0,0,231,0,42,0,0,0,161,0,0,0,235,0,0,0,203,0,171,0,79,0,67,0,173,0,246,0,212,0,37,0,155,0,53,0,50,0,0,0,133,0,159,0,0,0,242,0,162,0,170,0,224,0,194,0,126,0,153,0,23,0,0,0,219,0,211,0,254,0,254,0,154,0,136,0,240,0,109,0,0,0,130,0,0,0,82,0,88,0,35,0,95,0,107,0,0,0,22,0,0,0,0,0,248,0,0,0,117,0,151,0,243,0,67,0,207,0,9,0,183,0,229,0,148,0,92,0,129,0,0,0,233,0,154,0,216,0,0,0,234,0,46,0,161,0,0,0,140,0,10,0,110,0,52,0,64,0,237,0,15,0,54,0,176,0,85,0,193,0,0,0,46,0,124,0,89,0,167,0,102,0,93,0,242,0,103,0,207,0,56,0,252,0,0,0,59,0,213,0,35,0,128,0,0,0,154,0,0,0,48,0,153,0,21,0,214,0,120,0,201,0,0,0,179,0,174,0,0,0,143,0,141,0,9,0,111,0,224,0,142,0,251,0,162,0,195,0,127,0,36,0,245,0,51,0,112,0,24,0,124,0,5,0,235,0,183,0,47,0,12,0,167,0,39,0,19,0,40,0,28,0,242,0,0,0,109,0,223,0,151,0,118,0,75,0,43,0,0,0,207,0,35,0,0,0,125,0,204,0,0,0,240,0,0,0,243,0,17,0,225,0,158,0,50,0,51,0,219,0,237,0,163,0,167,0,0,0,181,0,16,0,0,0,44,0,113,0,8,0,0,0,104,0,0,0,96,0,77,0,135,0,105,0,21,0,109,0,0,0,184,0,97,0,152,0,67,0,73,0,239,0,139,0,197,0,103,0,40,0,39,0,253,0,168,0,4,0,190,0,0,0,181,0,0,0,126,0,219,0,184,0,87,0,223,0,96,0,0,0,7,0,0,0,148,0,0,0,212,0,46,0,102,0,9,0,125,0,208,0,114,0,26,0,171,0,128,0,188,0,129,0,231,0,114,0,0,0,144,0,24,0,72,0,253,0,78,0,196,0,239,0,0,0,0,0,92,0,161,0,55,0,35,0,96,0,75,0,0,0,24,0,69,0,67,0,54,0,195,0,0,0,255,0,0,0,62,0,244,0,205,0,0,0,175,0,8,0,254,0,172,0,51,0,141,0,0,0,144,0,204,0,108,0,133,0,51,0,74,0,110,0,131,0,58,0,0,0,0,0,190,0,47,0,39,0,223,0,51,0,114,0,163,0,218,0,204,0,101,0,12,0,120,0,74,0,104,0,95,0,205,0,47,0,50,0,0,0,143,0,151,0,0,0,5,0,128,0,177,0,0,0,87,0,0,0,205,0,223,0,46,0,0,0,165,0,0,0,160,0,115,0,252,0,51,0,126,0,0,0,85,0,0,0,184,0,29,0,255,0,0,0,64,0,118,0,58,0,100,0,0,0,123,0,8,0,0,0,132,0,224,0,153,0,0,0,193,0,244,0,112,0,143,0,150,0,104,0,143,0,240,0,159,0,221,0,156,0,41,0,116,0,128,0,0,0,88,0,204,0,187,0,0,0,72,0,120,0,64,0,39,0,89,0,171,0,119,0,8,0,66,0,178,0,112,0,0,0,10,0,8,0,0,0,100,0,13,0,158,0,0,0,192,0,152,0,221,0,229,0,219,0,92,0,0,0,117,0,212,0,0,0,161,0,150,0,191,0,130,0,190,0,169,0,0,0,137,0,31,0,243,0,152,0,0,0,97,0,0,0,2,0,242,0,112,0,133,0,39,0,246,0,0,0,0,0,104,0,0,0,80,0,83,0,77,0,8,0,19,0,27,0,221,0,192,0,166,0,130,0,73,0,200,0,0,0,77,0,189,0,221,0,126,0,0,0,132,0,47,0,201,0,139,0,0,0,29,0,0,0,0,0,92,0,183,0,235,0,128,0,38,0,0,0,255,0,0,0,132,0,168,0,104,0,251,0,8,0,239,0,185,0,47,0,131,0,188,0,174,0,198,0,0,0,183,0,214,0,0,0,60,0,59,0,215,0,187,0,73,0);
signal scenario_full  : scenario_type := (134,31,166,31,88,31,88,30,173,31,50,31,132,31,246,31,52,31,125,31,125,30,192,31,192,30,192,29,64,31,64,30,70,31,153,31,204,31,199,31,199,30,199,29,25,31,185,31,83,31,84,31,193,31,193,30,193,29,65,31,90,31,42,31,85,31,227,31,99,31,235,31,225,31,251,31,53,31,251,31,204,31,139,31,248,31,252,31,235,31,42,31,95,31,196,31,240,31,34,31,42,31,229,31,245,31,250,31,17,31,156,31,128,31,57,31,74,31,255,31,168,31,171,31,95,31,95,30,251,31,206,31,206,30,170,31,170,30,170,29,170,28,112,31,200,31,66,31,237,31,237,30,29,31,41,31,55,31,146,31,218,31,117,31,69,31,69,30,167,31,104,31,48,31,30,31,30,30,30,29,32,31,185,31,185,30,185,29,11,31,133,31,133,30,130,31,25,31,25,31,205,31,142,31,142,30,22,31,56,31,113,31,13,31,31,31,222,31,17,31,162,31,35,31,225,31,99,31,140,31,168,31,151,31,57,31,16,31,16,30,16,29,43,31,83,31,114,31,217,31,166,31,209,31,209,30,183,31,245,31,243,31,243,30,225,31,61,31,243,31,243,30,243,29,116,31,116,30,104,31,89,31,85,31,9,31,67,31,225,31,225,30,158,31,158,30,158,29,143,31,143,30,204,31,13,31,173,31,241,31,241,30,106,31,220,31,220,30,220,29,53,31,70,31,70,30,70,29,70,28,237,31,101,31,250,31,250,30,78,31,212,31,94,31,94,30,153,31,91,31,41,31,63,31,181,31,24,31,61,31,186,31,228,31,26,31,26,30,249,31,63,31,205,31,243,31,142,31,252,31,175,31,149,31,127,31,60,31,91,31,126,31,126,30,188,31,209,31,200,31,113,31,245,31,245,30,156,31,178,31,178,30,234,31,187,31,187,30,1,31,112,31,82,31,182,31,173,31,179,31,155,31,152,31,17,31,169,31,241,31,166,31,30,31,191,31,70,31,177,31,102,31,219,31,210,31,83,31,224,31,129,31,140,31,51,31,80,31,182,31,182,30,88,31,132,31,65,31,40,31,40,30,22,31,197,31,159,31,124,31,28,31,164,31,91,31,14,31,94,31,94,30,205,31,205,30,204,31,96,31,98,31,148,31,148,30,7,31,39,31,156,31,81,31,59,31,212,31,248,31,106,31,82,31,47,31,168,31,186,31,111,31,112,31,185,31,194,31,200,31,135,31,135,30,164,31,214,31,214,30,214,29,195,31,195,30,146,31,44,31,134,31,134,30,231,31,42,31,42,30,161,31,161,30,235,31,235,30,203,31,171,31,79,31,67,31,173,31,246,31,212,31,37,31,155,31,53,31,50,31,50,30,133,31,159,31,159,30,242,31,162,31,170,31,224,31,194,31,126,31,153,31,23,31,23,30,219,31,211,31,254,31,254,31,154,31,136,31,240,31,109,31,109,30,130,31,130,30,82,31,88,31,35,31,95,31,107,31,107,30,22,31,22,30,22,29,248,31,248,30,117,31,151,31,243,31,67,31,207,31,9,31,183,31,229,31,148,31,92,31,129,31,129,30,233,31,154,31,216,31,216,30,234,31,46,31,161,31,161,30,140,31,10,31,110,31,52,31,64,31,237,31,15,31,54,31,176,31,85,31,193,31,193,30,46,31,124,31,89,31,167,31,102,31,93,31,242,31,103,31,207,31,56,31,252,31,252,30,59,31,213,31,35,31,128,31,128,30,154,31,154,30,48,31,153,31,21,31,214,31,120,31,201,31,201,30,179,31,174,31,174,30,143,31,141,31,9,31,111,31,224,31,142,31,251,31,162,31,195,31,127,31,36,31,245,31,51,31,112,31,24,31,124,31,5,31,235,31,183,31,47,31,12,31,167,31,39,31,19,31,40,31,28,31,242,31,242,30,109,31,223,31,151,31,118,31,75,31,43,31,43,30,207,31,35,31,35,30,125,31,204,31,204,30,240,31,240,30,243,31,17,31,225,31,158,31,50,31,51,31,219,31,237,31,163,31,167,31,167,30,181,31,16,31,16,30,44,31,113,31,8,31,8,30,104,31,104,30,96,31,77,31,135,31,105,31,21,31,109,31,109,30,184,31,97,31,152,31,67,31,73,31,239,31,139,31,197,31,103,31,40,31,39,31,253,31,168,31,4,31,190,31,190,30,181,31,181,30,126,31,219,31,184,31,87,31,223,31,96,31,96,30,7,31,7,30,148,31,148,30,212,31,46,31,102,31,9,31,125,31,208,31,114,31,26,31,171,31,128,31,188,31,129,31,231,31,114,31,114,30,144,31,24,31,72,31,253,31,78,31,196,31,239,31,239,30,239,29,92,31,161,31,55,31,35,31,96,31,75,31,75,30,24,31,69,31,67,31,54,31,195,31,195,30,255,31,255,30,62,31,244,31,205,31,205,30,175,31,8,31,254,31,172,31,51,31,141,31,141,30,144,31,204,31,108,31,133,31,51,31,74,31,110,31,131,31,58,31,58,30,58,29,190,31,47,31,39,31,223,31,51,31,114,31,163,31,218,31,204,31,101,31,12,31,120,31,74,31,104,31,95,31,205,31,47,31,50,31,50,30,143,31,151,31,151,30,5,31,128,31,177,31,177,30,87,31,87,30,205,31,223,31,46,31,46,30,165,31,165,30,160,31,115,31,252,31,51,31,126,31,126,30,85,31,85,30,184,31,29,31,255,31,255,30,64,31,118,31,58,31,100,31,100,30,123,31,8,31,8,30,132,31,224,31,153,31,153,30,193,31,244,31,112,31,143,31,150,31,104,31,143,31,240,31,159,31,221,31,156,31,41,31,116,31,128,31,128,30,88,31,204,31,187,31,187,30,72,31,120,31,64,31,39,31,89,31,171,31,119,31,8,31,66,31,178,31,112,31,112,30,10,31,8,31,8,30,100,31,13,31,158,31,158,30,192,31,152,31,221,31,229,31,219,31,92,31,92,30,117,31,212,31,212,30,161,31,150,31,191,31,130,31,190,31,169,31,169,30,137,31,31,31,243,31,152,31,152,30,97,31,97,30,2,31,242,31,112,31,133,31,39,31,246,31,246,30,246,29,104,31,104,30,80,31,83,31,77,31,8,31,19,31,27,31,221,31,192,31,166,31,130,31,73,31,200,31,200,30,77,31,189,31,221,31,126,31,126,30,132,31,47,31,201,31,139,31,139,30,29,31,29,30,29,29,92,31,183,31,235,31,128,31,38,31,38,30,255,31,255,30,132,31,168,31,104,31,251,31,8,31,239,31,185,31,47,31,131,31,188,31,174,31,198,31,198,30,183,31,214,31,214,30,60,31,59,31,215,31,187,31,73,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
