-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 242;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (26,0,170,0,245,0,159,0,127,0,54,0,254,0,218,0,217,0,170,0,6,0,127,0,149,0,145,0,138,0,0,0,52,0,236,0,149,0,0,0,0,0,44,0,0,0,63,0,142,0,120,0,197,0,245,0,114,0,7,0,0,0,0,0,0,0,120,0,0,0,32,0,120,0,112,0,0,0,40,0,253,0,167,0,152,0,175,0,145,0,32,0,184,0,0,0,0,0,0,0,0,0,32,0,20,0,53,0,160,0,0,0,108,0,183,0,0,0,212,0,109,0,193,0,144,0,114,0,0,0,235,0,0,0,44,0,120,0,152,0,153,0,0,0,191,0,0,0,0,0,127,0,254,0,136,0,148,0,56,0,61,0,240,0,0,0,182,0,202,0,0,0,211,0,0,0,95,0,143,0,221,0,156,0,45,0,47,0,133,0,36,0,17,0,46,0,57,0,31,0,32,0,136,0,0,0,232,0,32,0,218,0,29,0,119,0,6,0,64,0,0,0,0,0,0,0,110,0,45,0,44,0,78,0,86,0,20,0,105,0,90,0,70,0,179,0,28,0,22,0,140,0,201,0,92,0,149,0,88,0,0,0,0,0,0,0,32,0,157,0,151,0,0,0,17,0,81,0,201,0,51,0,0,0,90,0,195,0,164,0,102,0,169,0,70,0,233,0,150,0,0,0,198,0,151,0,165,0,143,0,241,0,0,0,120,0,244,0,199,0,205,0,98,0,221,0,213,0,117,0,0,0,227,0,45,0,97,0,214,0,142,0,133,0,120,0,0,0,118,0,76,0,0,0,0,0,246,0,221,0,15,0,190,0,163,0,36,0,209,0,147,0,89,0,197,0,0,0,245,0,153,0,100,0,146,0,52,0,0,0,212,0,26,0,113,0,55,0,79,0,183,0,214,0,0,0,77,0,170,0,19,0,0,0,167,0,220,0,195,0,128,0,159,0,49,0,236,0,27,0,244,0,149,0,249,0,59,0,0,0,0,0,196,0,155,0,0,0,0,0,0,0,147,0,222,0,221,0,66,0,40,0,219,0,234,0,11,0,9,0,115,0,41,0,213,0,214,0,138,0,202,0,126,0);
signal scenario_full  : scenario_type := (26,31,170,31,245,31,159,31,127,31,54,31,254,31,218,31,217,31,170,31,6,31,127,31,149,31,145,31,138,31,138,30,52,31,236,31,149,31,149,30,149,29,44,31,44,30,63,31,142,31,120,31,197,31,245,31,114,31,7,31,7,30,7,29,7,28,120,31,120,30,32,31,120,31,112,31,112,30,40,31,253,31,167,31,152,31,175,31,145,31,32,31,184,31,184,30,184,29,184,28,184,27,32,31,20,31,53,31,160,31,160,30,108,31,183,31,183,30,212,31,109,31,193,31,144,31,114,31,114,30,235,31,235,30,44,31,120,31,152,31,153,31,153,30,191,31,191,30,191,29,127,31,254,31,136,31,148,31,56,31,61,31,240,31,240,30,182,31,202,31,202,30,211,31,211,30,95,31,143,31,221,31,156,31,45,31,47,31,133,31,36,31,17,31,46,31,57,31,31,31,32,31,136,31,136,30,232,31,32,31,218,31,29,31,119,31,6,31,64,31,64,30,64,29,64,28,110,31,45,31,44,31,78,31,86,31,20,31,105,31,90,31,70,31,179,31,28,31,22,31,140,31,201,31,92,31,149,31,88,31,88,30,88,29,88,28,32,31,157,31,151,31,151,30,17,31,81,31,201,31,51,31,51,30,90,31,195,31,164,31,102,31,169,31,70,31,233,31,150,31,150,30,198,31,151,31,165,31,143,31,241,31,241,30,120,31,244,31,199,31,205,31,98,31,221,31,213,31,117,31,117,30,227,31,45,31,97,31,214,31,142,31,133,31,120,31,120,30,118,31,76,31,76,30,76,29,246,31,221,31,15,31,190,31,163,31,36,31,209,31,147,31,89,31,197,31,197,30,245,31,153,31,100,31,146,31,52,31,52,30,212,31,26,31,113,31,55,31,79,31,183,31,214,31,214,30,77,31,170,31,19,31,19,30,167,31,220,31,195,31,128,31,159,31,49,31,236,31,27,31,244,31,149,31,249,31,59,31,59,30,59,29,196,31,155,31,155,30,155,29,155,28,147,31,222,31,221,31,66,31,40,31,219,31,234,31,11,31,9,31,115,31,41,31,213,31,214,31,138,31,202,31,126,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
