-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 541;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,223,0,81,0,190,0,0,0,136,0,90,0,0,0,213,0,0,0,0,0,4,0,23,0,0,0,165,0,167,0,95,0,93,0,129,0,94,0,221,0,222,0,179,0,0,0,234,0,119,0,134,0,159,0,0,0,36,0,93,0,65,0,51,0,42,0,251,0,13,0,72,0,243,0,0,0,165,0,117,0,195,0,0,0,61,0,77,0,230,0,232,0,195,0,80,0,244,0,107,0,0,0,150,0,240,0,165,0,247,0,17,0,58,0,241,0,71,0,9,0,246,0,0,0,30,0,0,0,68,0,225,0,241,0,219,0,0,0,10,0,164,0,0,0,0,0,77,0,181,0,227,0,0,0,0,0,249,0,0,0,156,0,239,0,230,0,175,0,26,0,203,0,94,0,75,0,173,0,153,0,79,0,213,0,34,0,93,0,103,0,236,0,93,0,232,0,0,0,116,0,144,0,101,0,0,0,87,0,43,0,0,0,63,0,0,0,188,0,116,0,0,0,213,0,0,0,235,0,218,0,74,0,37,0,122,0,118,0,222,0,0,0,131,0,108,0,0,0,0,0,66,0,216,0,196,0,193,0,0,0,0,0,0,0,87,0,218,0,212,0,159,0,25,0,158,0,69,0,5,0,150,0,159,0,241,0,222,0,0,0,170,0,26,0,118,0,0,0,0,0,216,0,105,0,153,0,14,0,0,0,232,0,200,0,188,0,182,0,118,0,58,0,208,0,158,0,0,0,226,0,137,0,54,0,111,0,26,0,88,0,0,0,206,0,198,0,254,0,180,0,152,0,207,0,112,0,32,0,241,0,163,0,124,0,1,0,199,0,122,0,0,0,0,0,0,0,94,0,0,0,0,0,208,0,33,0,145,0,0,0,247,0,110,0,195,0,190,0,253,0,4,0,40,0,180,0,166,0,189,0,244,0,178,0,0,0,115,0,145,0,0,0,37,0,174,0,57,0,178,0,213,0,147,0,14,0,92,0,192,0,42,0,0,0,242,0,0,0,112,0,0,0,222,0,20,0,16,0,0,0,44,0,25,0,5,0,213,0,0,0,23,0,164,0,0,0,104,0,220,0,157,0,8,0,0,0,150,0,137,0,238,0,231,0,12,0,0,0,222,0,32,0,70,0,244,0,0,0,32,0,0,0,202,0,200,0,0,0,18,0,5,0,0,0,84,0,160,0,0,0,253,0,209,0,0,0,1,0,44,0,120,0,161,0,0,0,201,0,221,0,0,0,61,0,186,0,39,0,146,0,0,0,197,0,20,0,20,0,187,0,0,0,60,0,236,0,110,0,199,0,77,0,0,0,54,0,0,0,251,0,29,0,167,0,96,0,108,0,62,0,235,0,32,0,230,0,28,0,133,0,214,0,197,0,78,0,0,0,223,0,234,0,51,0,46,0,223,0,174,0,197,0,192,0,209,0,50,0,135,0,1,0,173,0,131,0,16,0,174,0,226,0,0,0,254,0,162,0,141,0,80,0,0,0,247,0,59,0,102,0,0,0,0,0,141,0,223,0,0,0,69,0,53,0,135,0,157,0,0,0,0,0,79,0,99,0,0,0,71,0,88,0,211,0,79,0,130,0,168,0,8,0,201,0,119,0,253,0,108,0,241,0,238,0,161,0,139,0,149,0,73,0,247,0,84,0,0,0,251,0,250,0,57,0,0,0,155,0,52,0,0,0,2,0,59,0,226,0,188,0,173,0,182,0,228,0,123,0,244,0,92,0,33,0,44,0,37,0,0,0,0,0,0,0,0,0,130,0,0,0,21,0,48,0,0,0,0,0,225,0,238,0,121,0,0,0,173,0,39,0,230,0,80,0,197,0,0,0,221,0,240,0,179,0,0,0,221,0,0,0,228,0,136,0,0,0,18,0,0,0,0,0,44,0,180,0,245,0,148,0,177,0,0,0,169,0,118,0,141,0,163,0,188,0,51,0,147,0,236,0,2,0,23,0,54,0,171,0,242,0,235,0,0,0,251,0,243,0,169,0,157,0,209,0,15,0,34,0,58,0,0,0,31,0,102,0,164,0,72,0,32,0,135,0,0,0,169,0,155,0,12,0,111,0,0,0,158,0,0,0,41,0,165,0,6,0,85,0,196,0,201,0,41,0,193,0,76,0,220,0,24,0,123,0,24,0,169,0,66,0,52,0,218,0,102,0,12,0,136,0,0,0,133,0,0,0,252,0,116,0,237,0,46,0,0,0,28,0,29,0,85,0,138,0,0,0,4,0,0,0,0,0,88,0,56,0,204,0,210,0,254,0,43,0,245,0,11,0,28,0,180,0,0,0,128,0,0,0,246,0,135,0,244,0,99,0,213,0,0,0,0,0,0,0,221,0,0,0,0,0,8,0,177,0,29,0,133,0,0,0,157,0,0,0,82,0,137,0,97,0,92,0,239,0,112,0,77,0,52,0);
signal scenario_full  : scenario_type := (0,0,223,31,81,31,190,31,190,30,136,31,90,31,90,30,213,31,213,30,213,29,4,31,23,31,23,30,165,31,167,31,95,31,93,31,129,31,94,31,221,31,222,31,179,31,179,30,234,31,119,31,134,31,159,31,159,30,36,31,93,31,65,31,51,31,42,31,251,31,13,31,72,31,243,31,243,30,165,31,117,31,195,31,195,30,61,31,77,31,230,31,232,31,195,31,80,31,244,31,107,31,107,30,150,31,240,31,165,31,247,31,17,31,58,31,241,31,71,31,9,31,246,31,246,30,30,31,30,30,68,31,225,31,241,31,219,31,219,30,10,31,164,31,164,30,164,29,77,31,181,31,227,31,227,30,227,29,249,31,249,30,156,31,239,31,230,31,175,31,26,31,203,31,94,31,75,31,173,31,153,31,79,31,213,31,34,31,93,31,103,31,236,31,93,31,232,31,232,30,116,31,144,31,101,31,101,30,87,31,43,31,43,30,63,31,63,30,188,31,116,31,116,30,213,31,213,30,235,31,218,31,74,31,37,31,122,31,118,31,222,31,222,30,131,31,108,31,108,30,108,29,66,31,216,31,196,31,193,31,193,30,193,29,193,28,87,31,218,31,212,31,159,31,25,31,158,31,69,31,5,31,150,31,159,31,241,31,222,31,222,30,170,31,26,31,118,31,118,30,118,29,216,31,105,31,153,31,14,31,14,30,232,31,200,31,188,31,182,31,118,31,58,31,208,31,158,31,158,30,226,31,137,31,54,31,111,31,26,31,88,31,88,30,206,31,198,31,254,31,180,31,152,31,207,31,112,31,32,31,241,31,163,31,124,31,1,31,199,31,122,31,122,30,122,29,122,28,94,31,94,30,94,29,208,31,33,31,145,31,145,30,247,31,110,31,195,31,190,31,253,31,4,31,40,31,180,31,166,31,189,31,244,31,178,31,178,30,115,31,145,31,145,30,37,31,174,31,57,31,178,31,213,31,147,31,14,31,92,31,192,31,42,31,42,30,242,31,242,30,112,31,112,30,222,31,20,31,16,31,16,30,44,31,25,31,5,31,213,31,213,30,23,31,164,31,164,30,104,31,220,31,157,31,8,31,8,30,150,31,137,31,238,31,231,31,12,31,12,30,222,31,32,31,70,31,244,31,244,30,32,31,32,30,202,31,200,31,200,30,18,31,5,31,5,30,84,31,160,31,160,30,253,31,209,31,209,30,1,31,44,31,120,31,161,31,161,30,201,31,221,31,221,30,61,31,186,31,39,31,146,31,146,30,197,31,20,31,20,31,187,31,187,30,60,31,236,31,110,31,199,31,77,31,77,30,54,31,54,30,251,31,29,31,167,31,96,31,108,31,62,31,235,31,32,31,230,31,28,31,133,31,214,31,197,31,78,31,78,30,223,31,234,31,51,31,46,31,223,31,174,31,197,31,192,31,209,31,50,31,135,31,1,31,173,31,131,31,16,31,174,31,226,31,226,30,254,31,162,31,141,31,80,31,80,30,247,31,59,31,102,31,102,30,102,29,141,31,223,31,223,30,69,31,53,31,135,31,157,31,157,30,157,29,79,31,99,31,99,30,71,31,88,31,211,31,79,31,130,31,168,31,8,31,201,31,119,31,253,31,108,31,241,31,238,31,161,31,139,31,149,31,73,31,247,31,84,31,84,30,251,31,250,31,57,31,57,30,155,31,52,31,52,30,2,31,59,31,226,31,188,31,173,31,182,31,228,31,123,31,244,31,92,31,33,31,44,31,37,31,37,30,37,29,37,28,37,27,130,31,130,30,21,31,48,31,48,30,48,29,225,31,238,31,121,31,121,30,173,31,39,31,230,31,80,31,197,31,197,30,221,31,240,31,179,31,179,30,221,31,221,30,228,31,136,31,136,30,18,31,18,30,18,29,44,31,180,31,245,31,148,31,177,31,177,30,169,31,118,31,141,31,163,31,188,31,51,31,147,31,236,31,2,31,23,31,54,31,171,31,242,31,235,31,235,30,251,31,243,31,169,31,157,31,209,31,15,31,34,31,58,31,58,30,31,31,102,31,164,31,72,31,32,31,135,31,135,30,169,31,155,31,12,31,111,31,111,30,158,31,158,30,41,31,165,31,6,31,85,31,196,31,201,31,41,31,193,31,76,31,220,31,24,31,123,31,24,31,169,31,66,31,52,31,218,31,102,31,12,31,136,31,136,30,133,31,133,30,252,31,116,31,237,31,46,31,46,30,28,31,29,31,85,31,138,31,138,30,4,31,4,30,4,29,88,31,56,31,204,31,210,31,254,31,43,31,245,31,11,31,28,31,180,31,180,30,128,31,128,30,246,31,135,31,244,31,99,31,213,31,213,30,213,29,213,28,221,31,221,30,221,29,8,31,177,31,29,31,133,31,133,30,157,31,157,30,82,31,137,31,97,31,92,31,239,31,112,31,77,31,52,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
