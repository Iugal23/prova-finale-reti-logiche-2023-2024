-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_589 is
end project_tb_589;

architecture project_tb_arch_589 of project_tb_589 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 695;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (106,0,0,0,249,0,177,0,0,0,53,0,171,0,79,0,64,0,106,0,112,0,21,0,143,0,16,0,253,0,6,0,0,0,0,0,81,0,236,0,207,0,151,0,0,0,198,0,117,0,79,0,94,0,1,0,0,0,0,0,86,0,222,0,131,0,0,0,0,0,81,0,235,0,221,0,141,0,0,0,117,0,250,0,0,0,76,0,0,0,217,0,52,0,148,0,83,0,53,0,227,0,0,0,63,0,3,0,222,0,0,0,132,0,114,0,0,0,0,0,58,0,112,0,16,0,71,0,76,0,172,0,229,0,16,0,246,0,242,0,82,0,0,0,0,0,200,0,77,0,92,0,43,0,32,0,19,0,0,0,185,0,18,0,217,0,59,0,13,0,35,0,255,0,204,0,235,0,27,0,0,0,208,0,211,0,200,0,164,0,158,0,205,0,0,0,140,0,0,0,204,0,216,0,0,0,171,0,194,0,21,0,232,0,232,0,246,0,112,0,160,0,5,0,0,0,246,0,73,0,0,0,26,0,106,0,224,0,57,0,148,0,54,0,0,0,35,0,136,0,0,0,222,0,243,0,0,0,120,0,238,0,182,0,83,0,5,0,177,0,154,0,55,0,73,0,225,0,43,0,218,0,0,0,189,0,90,0,4,0,0,0,23,0,86,0,252,0,207,0,90,0,168,0,36,0,0,0,123,0,254,0,232,0,49,0,0,0,0,0,158,0,30,0,162,0,155,0,168,0,0,0,0,0,212,0,0,0,60,0,125,0,164,0,198,0,1,0,114,0,0,0,249,0,78,0,111,0,6,0,3,0,203,0,216,0,0,0,64,0,178,0,52,0,192,0,213,0,52,0,182,0,0,0,190,0,208,0,248,0,0,0,0,0,0,0,2,0,63,0,234,0,2,0,20,0,146,0,103,0,194,0,0,0,12,0,0,0,14,0,0,0,248,0,72,0,182,0,245,0,60,0,98,0,78,0,0,0,138,0,172,0,241,0,244,0,228,0,101,0,0,0,18,0,215,0,38,0,111,0,67,0,154,0,144,0,239,0,120,0,0,0,56,0,187,0,0,0,218,0,18,0,0,0,82,0,0,0,182,0,123,0,130,0,77,0,134,0,0,0,0,0,36,0,0,0,0,0,43,0,231,0,25,0,230,0,0,0,230,0,18,0,191,0,109,0,241,0,0,0,89,0,231,0,127,0,130,0,109,0,0,0,176,0,6,0,89,0,0,0,181,0,213,0,251,0,50,0,220,0,7,0,61,0,226,0,102,0,176,0,163,0,0,0,97,0,47,0,0,0,118,0,0,0,116,0,48,0,37,0,179,0,26,0,63,0,239,0,0,0,131,0,129,0,0,0,0,0,112,0,101,0,169,0,60,0,55,0,59,0,77,0,160,0,235,0,16,0,196,0,0,0,198,0,199,0,251,0,86,0,0,0,0,0,197,0,28,0,197,0,9,0,185,0,0,0,249,0,238,0,41,0,0,0,0,0,102,0,231,0,0,0,0,0,67,0,66,0,9,0,139,0,213,0,197,0,9,0,100,0,12,0,0,0,124,0,0,0,108,0,109,0,45,0,0,0,0,0,160,0,0,0,170,0,95,0,0,0,37,0,221,0,0,0,13,0,142,0,91,0,0,0,130,0,70,0,0,0,0,0,190,0,20,0,159,0,127,0,231,0,59,0,0,0,172,0,0,0,0,0,0,0,19,0,38,0,231,0,105,0,0,0,228,0,113,0,0,0,242,0,135,0,230,0,65,0,105,0,62,0,181,0,43,0,113,0,135,0,187,0,254,0,149,0,0,0,244,0,52,0,183,0,113,0,167,0,0,0,247,0,0,0,0,0,160,0,30,0,0,0,147,0,184,0,0,0,117,0,92,0,211,0,211,0,68,0,33,0,55,0,0,0,0,0,166,0,0,0,99,0,42,0,74,0,132,0,0,0,187,0,227,0,126,0,208,0,0,0,154,0,26,0,166,0,27,0,237,0,39,0,49,0,251,0,34,0,0,0,118,0,33,0,0,0,255,0,0,0,149,0,109,0,0,0,215,0,80,0,248,0,94,0,77,0,81,0,125,0,243,0,138,0,129,0,224,0,81,0,160,0,0,0,248,0,58,0,138,0,0,0,167,0,76,0,0,0,0,0,63,0,255,0,0,0,219,0,52,0,174,0,173,0,36,0,126,0,3,0,18,0,59,0,182,0,13,0,43,0,7,0,0,0,107,0,226,0,129,0,224,0,120,0,195,0,178,0,225,0,0,0,177,0,190,0,160,0,0,0,221,0,14,0,47,0,172,0,0,0,185,0,1,0,78,0,118,0,104,0,223,0,215,0,214,0,83,0,188,0,158,0,49,0,125,0,163,0,155,0,123,0,0,0,198,0,81,0,38,0,208,0,85,0,223,0,0,0,24,0,0,0,171,0,38,0,191,0,241,0,96,0,129,0,232,0,247,0,0,0,217,0,105,0,12,0,0,0,93,0,1,0,7,0,8,0,69,0,112,0,127,0,23,0,247,0,134,0,173,0,38,0,18,0,0,0,0,0,77,0,80,0,13,0,0,0,144,0,0,0,0,0,144,0,184,0,74,0,97,0,225,0,0,0,35,0,72,0,89,0,0,0,222,0,0,0,144,0,19,0,108,0,0,0,0,0,143,0,0,0,33,0,223,0,175,0,134,0,138,0,224,0,57,0,0,0,48,0,25,0,0,0,90,0,31,0,225,0,75,0,71,0,231,0,235,0,108,0,248,0,0,0,0,0,0,0,87,0,0,0,41,0,59,0,222,0,191,0,158,0,0,0,69,0,0,0,36,0,112,0,201,0,89,0,0,0,1,0,239,0,33,0,111,0,132,0,19,0,128,0,0,0,35,0,66,0,209,0,200,0,105,0,148,0,234,0,99,0,194,0,0,0,207,0,140,0,0,0,189,0,27,0,160,0,230,0,96,0,226,0,19,0,228,0,56,0,230,0,48,0,182,0,216,0,214,0,199,0,131,0,118,0,39,0,177,0,110,0,11,0,106,0,121,0,3,0,172,0,69,0,144,0,0,0,200,0,253,0,139,0,196,0,0,0,172,0,45,0,191,0,142,0,243,0,84,0,96,0,0,0,0,0);
signal scenario_full  : scenario_type := (106,31,106,30,249,31,177,31,177,30,53,31,171,31,79,31,64,31,106,31,112,31,21,31,143,31,16,31,253,31,6,31,6,30,6,29,81,31,236,31,207,31,151,31,151,30,198,31,117,31,79,31,94,31,1,31,1,30,1,29,86,31,222,31,131,31,131,30,131,29,81,31,235,31,221,31,141,31,141,30,117,31,250,31,250,30,76,31,76,30,217,31,52,31,148,31,83,31,53,31,227,31,227,30,63,31,3,31,222,31,222,30,132,31,114,31,114,30,114,29,58,31,112,31,16,31,71,31,76,31,172,31,229,31,16,31,246,31,242,31,82,31,82,30,82,29,200,31,77,31,92,31,43,31,32,31,19,31,19,30,185,31,18,31,217,31,59,31,13,31,35,31,255,31,204,31,235,31,27,31,27,30,208,31,211,31,200,31,164,31,158,31,205,31,205,30,140,31,140,30,204,31,216,31,216,30,171,31,194,31,21,31,232,31,232,31,246,31,112,31,160,31,5,31,5,30,246,31,73,31,73,30,26,31,106,31,224,31,57,31,148,31,54,31,54,30,35,31,136,31,136,30,222,31,243,31,243,30,120,31,238,31,182,31,83,31,5,31,177,31,154,31,55,31,73,31,225,31,43,31,218,31,218,30,189,31,90,31,4,31,4,30,23,31,86,31,252,31,207,31,90,31,168,31,36,31,36,30,123,31,254,31,232,31,49,31,49,30,49,29,158,31,30,31,162,31,155,31,168,31,168,30,168,29,212,31,212,30,60,31,125,31,164,31,198,31,1,31,114,31,114,30,249,31,78,31,111,31,6,31,3,31,203,31,216,31,216,30,64,31,178,31,52,31,192,31,213,31,52,31,182,31,182,30,190,31,208,31,248,31,248,30,248,29,248,28,2,31,63,31,234,31,2,31,20,31,146,31,103,31,194,31,194,30,12,31,12,30,14,31,14,30,248,31,72,31,182,31,245,31,60,31,98,31,78,31,78,30,138,31,172,31,241,31,244,31,228,31,101,31,101,30,18,31,215,31,38,31,111,31,67,31,154,31,144,31,239,31,120,31,120,30,56,31,187,31,187,30,218,31,18,31,18,30,82,31,82,30,182,31,123,31,130,31,77,31,134,31,134,30,134,29,36,31,36,30,36,29,43,31,231,31,25,31,230,31,230,30,230,31,18,31,191,31,109,31,241,31,241,30,89,31,231,31,127,31,130,31,109,31,109,30,176,31,6,31,89,31,89,30,181,31,213,31,251,31,50,31,220,31,7,31,61,31,226,31,102,31,176,31,163,31,163,30,97,31,47,31,47,30,118,31,118,30,116,31,48,31,37,31,179,31,26,31,63,31,239,31,239,30,131,31,129,31,129,30,129,29,112,31,101,31,169,31,60,31,55,31,59,31,77,31,160,31,235,31,16,31,196,31,196,30,198,31,199,31,251,31,86,31,86,30,86,29,197,31,28,31,197,31,9,31,185,31,185,30,249,31,238,31,41,31,41,30,41,29,102,31,231,31,231,30,231,29,67,31,66,31,9,31,139,31,213,31,197,31,9,31,100,31,12,31,12,30,124,31,124,30,108,31,109,31,45,31,45,30,45,29,160,31,160,30,170,31,95,31,95,30,37,31,221,31,221,30,13,31,142,31,91,31,91,30,130,31,70,31,70,30,70,29,190,31,20,31,159,31,127,31,231,31,59,31,59,30,172,31,172,30,172,29,172,28,19,31,38,31,231,31,105,31,105,30,228,31,113,31,113,30,242,31,135,31,230,31,65,31,105,31,62,31,181,31,43,31,113,31,135,31,187,31,254,31,149,31,149,30,244,31,52,31,183,31,113,31,167,31,167,30,247,31,247,30,247,29,160,31,30,31,30,30,147,31,184,31,184,30,117,31,92,31,211,31,211,31,68,31,33,31,55,31,55,30,55,29,166,31,166,30,99,31,42,31,74,31,132,31,132,30,187,31,227,31,126,31,208,31,208,30,154,31,26,31,166,31,27,31,237,31,39,31,49,31,251,31,34,31,34,30,118,31,33,31,33,30,255,31,255,30,149,31,109,31,109,30,215,31,80,31,248,31,94,31,77,31,81,31,125,31,243,31,138,31,129,31,224,31,81,31,160,31,160,30,248,31,58,31,138,31,138,30,167,31,76,31,76,30,76,29,63,31,255,31,255,30,219,31,52,31,174,31,173,31,36,31,126,31,3,31,18,31,59,31,182,31,13,31,43,31,7,31,7,30,107,31,226,31,129,31,224,31,120,31,195,31,178,31,225,31,225,30,177,31,190,31,160,31,160,30,221,31,14,31,47,31,172,31,172,30,185,31,1,31,78,31,118,31,104,31,223,31,215,31,214,31,83,31,188,31,158,31,49,31,125,31,163,31,155,31,123,31,123,30,198,31,81,31,38,31,208,31,85,31,223,31,223,30,24,31,24,30,171,31,38,31,191,31,241,31,96,31,129,31,232,31,247,31,247,30,217,31,105,31,12,31,12,30,93,31,1,31,7,31,8,31,69,31,112,31,127,31,23,31,247,31,134,31,173,31,38,31,18,31,18,30,18,29,77,31,80,31,13,31,13,30,144,31,144,30,144,29,144,31,184,31,74,31,97,31,225,31,225,30,35,31,72,31,89,31,89,30,222,31,222,30,144,31,19,31,108,31,108,30,108,29,143,31,143,30,33,31,223,31,175,31,134,31,138,31,224,31,57,31,57,30,48,31,25,31,25,30,90,31,31,31,225,31,75,31,71,31,231,31,235,31,108,31,248,31,248,30,248,29,248,28,87,31,87,30,41,31,59,31,222,31,191,31,158,31,158,30,69,31,69,30,36,31,112,31,201,31,89,31,89,30,1,31,239,31,33,31,111,31,132,31,19,31,128,31,128,30,35,31,66,31,209,31,200,31,105,31,148,31,234,31,99,31,194,31,194,30,207,31,140,31,140,30,189,31,27,31,160,31,230,31,96,31,226,31,19,31,228,31,56,31,230,31,48,31,182,31,216,31,214,31,199,31,131,31,118,31,39,31,177,31,110,31,11,31,106,31,121,31,3,31,172,31,69,31,144,31,144,30,200,31,253,31,139,31,196,31,196,30,172,31,45,31,191,31,142,31,243,31,84,31,96,31,96,30,96,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
