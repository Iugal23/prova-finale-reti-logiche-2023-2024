-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_294 is
end project_tb_294;

architecture project_tb_arch_294 of project_tb_294 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 536;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (157,0,94,0,223,0,0,0,243,0,235,0,92,0,0,0,11,0,135,0,7,0,227,0,50,0,0,0,243,0,156,0,0,0,0,0,69,0,215,0,0,0,86,0,8,0,100,0,128,0,248,0,214,0,216,0,116,0,117,0,149,0,255,0,201,0,0,0,150,0,48,0,78,0,173,0,12,0,0,0,167,0,36,0,217,0,140,0,0,0,142,0,207,0,0,0,204,0,61,0,50,0,241,0,75,0,131,0,0,0,119,0,52,0,48,0,18,0,188,0,0,0,84,0,130,0,125,0,56,0,254,0,221,0,0,0,163,0,21,0,140,0,159,0,122,0,43,0,0,0,30,0,233,0,226,0,0,0,137,0,169,0,6,0,44,0,253,0,204,0,113,0,202,0,45,0,166,0,172,0,0,0,125,0,0,0,0,0,228,0,137,0,242,0,12,0,220,0,159,0,149,0,11,0,195,0,0,0,1,0,228,0,211,0,43,0,0,0,0,0,154,0,57,0,0,0,0,0,202,0,19,0,10,0,211,0,109,0,67,0,0,0,63,0,145,0,1,0,152,0,82,0,224,0,87,0,115,0,71,0,53,0,54,0,92,0,201,0,100,0,101,0,171,0,180,0,111,0,201,0,238,0,131,0,84,0,88,0,153,0,14,0,93,0,70,0,70,0,10,0,194,0,0,0,125,0,174,0,127,0,123,0,177,0,0,0,39,0,23,0,225,0,233,0,86,0,0,0,0,0,118,0,42,0,48,0,20,0,32,0,145,0,0,0,21,0,151,0,245,0,209,0,231,0,178,0,160,0,154,0,181,0,172,0,0,0,0,0,193,0,76,0,112,0,193,0,0,0,0,0,97,0,191,0,113,0,11,0,85,0,3,0,194,0,235,0,218,0,218,0,175,0,0,0,182,0,64,0,24,0,202,0,119,0,64,0,57,0,0,0,181,0,242,0,123,0,232,0,163,0,230,0,0,0,0,0,69,0,26,0,199,0,0,0,68,0,101,0,177,0,1,0,64,0,194,0,11,0,0,0,79,0,0,0,112,0,113,0,229,0,190,0,127,0,241,0,170,0,152,0,23,0,191,0,0,0,56,0,95,0,84,0,61,0,32,0,0,0,179,0,210,0,44,0,0,0,248,0,0,0,21,0,158,0,226,0,0,0,16,0,0,0,141,0,242,0,0,0,198,0,166,0,158,0,53,0,192,0,0,0,40,0,199,0,41,0,28,0,0,0,61,0,123,0,0,0,183,0,0,0,0,0,238,0,44,0,0,0,169,0,0,0,41,0,221,0,235,0,140,0,20,0,46,0,66,0,0,0,39,0,145,0,3,0,36,0,200,0,151,0,80,0,85,0,0,0,0,0,137,0,0,0,152,0,76,0,164,0,0,0,40,0,130,0,224,0,0,0,201,0,107,0,185,0,78,0,249,0,124,0,38,0,0,0,50,0,0,0,243,0,162,0,0,0,57,0,209,0,230,0,231,0,29,0,122,0,183,0,129,0,0,0,74,0,0,0,187,0,0,0,56,0,129,0,2,0,143,0,0,0,158,0,236,0,197,0,228,0,130,0,150,0,148,0,49,0,38,0,35,0,0,0,144,0,221,0,22,0,37,0,63,0,246,0,117,0,200,0,123,0,163,0,228,0,173,0,186,0,168,0,230,0,157,0,199,0,228,0,203,0,200,0,0,0,208,0,16,0,140,0,74,0,244,0,0,0,227,0,202,0,103,0,0,0,160,0,110,0,167,0,203,0,38,0,242,0,0,0,120,0,102,0,221,0,0,0,149,0,248,0,133,0,0,0,143,0,101,0,68,0,45,0,191,0,0,0,164,0,69,0,0,0,65,0,0,0,37,0,96,0,153,0,147,0,10,0,125,0,172,0,105,0,0,0,71,0,143,0,47,0,175,0,232,0,197,0,0,0,233,0,157,0,0,0,195,0,142,0,227,0,27,0,68,0,111,0,59,0,142,0,68,0,23,0,28,0,0,0,144,0,149,0,1,0,72,0,0,0,0,0,0,0,130,0,0,0,179,0,120,0,200,0,80,0,191,0,0,0,187,0,250,0,0,0,136,0,11,0,164,0,27,0,138,0,248,0,58,0,44,0,58,0,116,0,174,0,245,0,136,0,54,0,147,0,0,0,13,0,194,0,26,0,104,0,112,0,172,0,0,0,38,0,23,0,0,0,229,0,0,0,198,0,38,0,0,0,79,0,244,0,0,0,92,0,32,0,227,0,0,0,139,0,45,0,138,0,177,0,187,0,33,0,17,0,26,0,4,0,131,0,181,0,188,0,0,0,0,0,170,0,13,0,136,0,109,0,131,0,225,0,243,0,108,0,16,0,73,0,29,0,93,0,178,0,102,0,0,0,234,0,0,0,175,0,233,0,84,0,0,0,223,0);
signal scenario_full  : scenario_type := (157,31,94,31,223,31,223,30,243,31,235,31,92,31,92,30,11,31,135,31,7,31,227,31,50,31,50,30,243,31,156,31,156,30,156,29,69,31,215,31,215,30,86,31,8,31,100,31,128,31,248,31,214,31,216,31,116,31,117,31,149,31,255,31,201,31,201,30,150,31,48,31,78,31,173,31,12,31,12,30,167,31,36,31,217,31,140,31,140,30,142,31,207,31,207,30,204,31,61,31,50,31,241,31,75,31,131,31,131,30,119,31,52,31,48,31,18,31,188,31,188,30,84,31,130,31,125,31,56,31,254,31,221,31,221,30,163,31,21,31,140,31,159,31,122,31,43,31,43,30,30,31,233,31,226,31,226,30,137,31,169,31,6,31,44,31,253,31,204,31,113,31,202,31,45,31,166,31,172,31,172,30,125,31,125,30,125,29,228,31,137,31,242,31,12,31,220,31,159,31,149,31,11,31,195,31,195,30,1,31,228,31,211,31,43,31,43,30,43,29,154,31,57,31,57,30,57,29,202,31,19,31,10,31,211,31,109,31,67,31,67,30,63,31,145,31,1,31,152,31,82,31,224,31,87,31,115,31,71,31,53,31,54,31,92,31,201,31,100,31,101,31,171,31,180,31,111,31,201,31,238,31,131,31,84,31,88,31,153,31,14,31,93,31,70,31,70,31,10,31,194,31,194,30,125,31,174,31,127,31,123,31,177,31,177,30,39,31,23,31,225,31,233,31,86,31,86,30,86,29,118,31,42,31,48,31,20,31,32,31,145,31,145,30,21,31,151,31,245,31,209,31,231,31,178,31,160,31,154,31,181,31,172,31,172,30,172,29,193,31,76,31,112,31,193,31,193,30,193,29,97,31,191,31,113,31,11,31,85,31,3,31,194,31,235,31,218,31,218,31,175,31,175,30,182,31,64,31,24,31,202,31,119,31,64,31,57,31,57,30,181,31,242,31,123,31,232,31,163,31,230,31,230,30,230,29,69,31,26,31,199,31,199,30,68,31,101,31,177,31,1,31,64,31,194,31,11,31,11,30,79,31,79,30,112,31,113,31,229,31,190,31,127,31,241,31,170,31,152,31,23,31,191,31,191,30,56,31,95,31,84,31,61,31,32,31,32,30,179,31,210,31,44,31,44,30,248,31,248,30,21,31,158,31,226,31,226,30,16,31,16,30,141,31,242,31,242,30,198,31,166,31,158,31,53,31,192,31,192,30,40,31,199,31,41,31,28,31,28,30,61,31,123,31,123,30,183,31,183,30,183,29,238,31,44,31,44,30,169,31,169,30,41,31,221,31,235,31,140,31,20,31,46,31,66,31,66,30,39,31,145,31,3,31,36,31,200,31,151,31,80,31,85,31,85,30,85,29,137,31,137,30,152,31,76,31,164,31,164,30,40,31,130,31,224,31,224,30,201,31,107,31,185,31,78,31,249,31,124,31,38,31,38,30,50,31,50,30,243,31,162,31,162,30,57,31,209,31,230,31,231,31,29,31,122,31,183,31,129,31,129,30,74,31,74,30,187,31,187,30,56,31,129,31,2,31,143,31,143,30,158,31,236,31,197,31,228,31,130,31,150,31,148,31,49,31,38,31,35,31,35,30,144,31,221,31,22,31,37,31,63,31,246,31,117,31,200,31,123,31,163,31,228,31,173,31,186,31,168,31,230,31,157,31,199,31,228,31,203,31,200,31,200,30,208,31,16,31,140,31,74,31,244,31,244,30,227,31,202,31,103,31,103,30,160,31,110,31,167,31,203,31,38,31,242,31,242,30,120,31,102,31,221,31,221,30,149,31,248,31,133,31,133,30,143,31,101,31,68,31,45,31,191,31,191,30,164,31,69,31,69,30,65,31,65,30,37,31,96,31,153,31,147,31,10,31,125,31,172,31,105,31,105,30,71,31,143,31,47,31,175,31,232,31,197,31,197,30,233,31,157,31,157,30,195,31,142,31,227,31,27,31,68,31,111,31,59,31,142,31,68,31,23,31,28,31,28,30,144,31,149,31,1,31,72,31,72,30,72,29,72,28,130,31,130,30,179,31,120,31,200,31,80,31,191,31,191,30,187,31,250,31,250,30,136,31,11,31,164,31,27,31,138,31,248,31,58,31,44,31,58,31,116,31,174,31,245,31,136,31,54,31,147,31,147,30,13,31,194,31,26,31,104,31,112,31,172,31,172,30,38,31,23,31,23,30,229,31,229,30,198,31,38,31,38,30,79,31,244,31,244,30,92,31,32,31,227,31,227,30,139,31,45,31,138,31,177,31,187,31,33,31,17,31,26,31,4,31,131,31,181,31,188,31,188,30,188,29,170,31,13,31,136,31,109,31,131,31,225,31,243,31,108,31,16,31,73,31,29,31,93,31,178,31,102,31,102,30,234,31,234,30,175,31,233,31,84,31,84,30,223,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
