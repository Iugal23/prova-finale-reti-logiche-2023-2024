-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_146 is
end project_tb_146;

architecture project_tb_arch_146 of project_tb_146 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 623;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (248,0,97,0,245,0,114,0,0,0,70,0,117,0,100,0,201,0,217,0,0,0,126,0,86,0,174,0,44,0,82,0,248,0,183,0,138,0,241,0,0,0,0,0,223,0,48,0,26,0,0,0,138,0,47,0,196,0,238,0,240,0,183,0,179,0,58,0,240,0,152,0,141,0,0,0,0,0,61,0,0,0,0,0,0,0,0,0,213,0,157,0,113,0,160,0,157,0,0,0,70,0,181,0,0,0,168,0,212,0,57,0,147,0,0,0,88,0,141,0,186,0,0,0,39,0,30,0,0,0,0,0,58,0,247,0,224,0,81,0,217,0,121,0,0,0,5,0,224,0,47,0,0,0,212,0,145,0,0,0,87,0,64,0,153,0,111,0,239,0,0,0,121,0,179,0,151,0,0,0,17,0,180,0,72,0,116,0,0,0,92,0,249,0,247,0,182,0,38,0,5,0,0,0,61,0,108,0,50,0,254,0,0,0,86,0,176,0,36,0,0,0,161,0,0,0,251,0,0,0,74,0,195,0,0,0,6,0,186,0,0,0,0,0,157,0,160,0,23,0,190,0,223,0,141,0,0,0,224,0,0,0,54,0,245,0,0,0,62,0,225,0,0,0,0,0,30,0,0,0,207,0,84,0,145,0,154,0,233,0,18,0,116,0,0,0,207,0,139,0,0,0,22,0,164,0,126,0,82,0,176,0,153,0,147,0,134,0,0,0,192,0,229,0,9,0,124,0,40,0,105,0,231,0,190,0,118,0,0,0,30,0,239,0,148,0,0,0,248,0,137,0,0,0,209,0,0,0,116,0,66,0,200,0,178,0,0,0,255,0,28,0,224,0,107,0,85,0,24,0,8,0,0,0,201,0,169,0,0,0,130,0,209,0,211,0,135,0,0,0,0,0,4,0,156,0,0,0,77,0,88,0,185,0,153,0,196,0,146,0,128,0,146,0,0,0,0,0,246,0,182,0,225,0,213,0,102,0,52,0,138,0,0,0,194,0,82,0,48,0,0,0,182,0,150,0,28,0,243,0,0,0,180,0,222,0,102,0,0,0,0,0,10,0,223,0,210,0,68,0,199,0,171,0,102,0,211,0,183,0,170,0,210,0,142,0,18,0,231,0,107,0,1,0,38,0,0,0,0,0,0,0,121,0,73,0,0,0,183,0,0,0,227,0,133,0,117,0,77,0,87,0,0,0,0,0,0,0,133,0,189,0,242,0,7,0,101,0,0,0,0,0,25,0,53,0,215,0,205,0,212,0,49,0,225,0,249,0,226,0,244,0,12,0,94,0,137,0,229,0,20,0,132,0,216,0,0,0,72,0,231,0,69,0,0,0,0,0,11,0,202,0,115,0,208,0,200,0,135,0,202,0,0,0,83,0,154,0,248,0,177,0,0,0,45,0,40,0,218,0,0,0,106,0,0,0,115,0,78,0,0,0,0,0,208,0,231,0,217,0,84,0,182,0,192,0,11,0,9,0,244,0,63,0,71,0,186,0,191,0,83,0,12,0,43,0,0,0,7,0,3,0,141,0,148,0,37,0,0,0,23,0,253,0,114,0,0,0,55,0,84,0,0,0,208,0,121,0,233,0,0,0,205,0,17,0,22,0,8,0,0,0,70,0,187,0,183,0,19,0,0,0,77,0,0,0,220,0,0,0,224,0,113,0,76,0,1,0,0,0,0,0,228,0,154,0,248,0,0,0,79,0,249,0,131,0,130,0,86,0,11,0,215,0,20,0,50,0,0,0,240,0,15,0,146,0,241,0,229,0,185,0,0,0,217,0,67,0,144,0,99,0,0,0,0,0,29,0,13,0,42,0,252,0,118,0,44,0,210,0,0,0,0,0,69,0,122,0,84,0,52,0,113,0,148,0,177,0,165,0,0,0,254,0,0,0,136,0,154,0,0,0,164,0,30,0,231,0,118,0,0,0,0,0,25,0,85,0,70,0,151,0,70,0,107,0,0,0,134,0,64,0,0,0,24,0,38,0,79,0,200,0,82,0,66,0,95,0,202,0,0,0,6,0,62,0,95,0,149,0,137,0,174,0,25,0,162,0,0,0,209,0,0,0,111,0,221,0,35,0,220,0,119,0,68,0,10,0,21,0,19,0,159,0,78,0,208,0,221,0,239,0,172,0,34,0,121,0,45,0,133,0,98,0,95,0,39,0,206,0,0,0,232,0,8,0,199,0,243,0,41,0,0,0,212,0,0,0,0,0,201,0,130,0,114,0,231,0,0,0,39,0,0,0,191,0,0,0,37,0,184,0,103,0,197,0,59,0,32,0,0,0,173,0,47,0,49,0,225,0,27,0,70,0,49,0,227,0,185,0,107,0,89,0,119,0,159,0,0,0,20,0,110,0,131,0,135,0,156,0,112,0,177,0,187,0,84,0,234,0,50,0,202,0,0,0,195,0,237,0,0,0,0,0,213,0,109,0,54,0,217,0,0,0,206,0,116,0,5,0,182,0,25,0,166,0,106,0,95,0,0,0,0,0,44,0,0,0,153,0,252,0,0,0,20,0,0,0,56,0,110,0,87,0,128,0,179,0,147,0,0,0,93,0,221,0,232,0,209,0,41,0,9,0,176,0,168,0,82,0,101,0,11,0,156,0,0,0,196,0,252,0,167,0,126,0,24,0,143,0,189,0,50,0,131,0,0,0,102,0,132,0,91,0,88,0,101,0,220,0,223,0,0,0,206,0,103,0,204,0,0,0,222,0,245,0,223,0,202,0,150,0,0,0,0,0,0,0,63,0,159,0,121,0,24,0,0,0,206,0,222,0,95,0,150,0);
signal scenario_full  : scenario_type := (248,31,97,31,245,31,114,31,114,30,70,31,117,31,100,31,201,31,217,31,217,30,126,31,86,31,174,31,44,31,82,31,248,31,183,31,138,31,241,31,241,30,241,29,223,31,48,31,26,31,26,30,138,31,47,31,196,31,238,31,240,31,183,31,179,31,58,31,240,31,152,31,141,31,141,30,141,29,61,31,61,30,61,29,61,28,61,27,213,31,157,31,113,31,160,31,157,31,157,30,70,31,181,31,181,30,168,31,212,31,57,31,147,31,147,30,88,31,141,31,186,31,186,30,39,31,30,31,30,30,30,29,58,31,247,31,224,31,81,31,217,31,121,31,121,30,5,31,224,31,47,31,47,30,212,31,145,31,145,30,87,31,64,31,153,31,111,31,239,31,239,30,121,31,179,31,151,31,151,30,17,31,180,31,72,31,116,31,116,30,92,31,249,31,247,31,182,31,38,31,5,31,5,30,61,31,108,31,50,31,254,31,254,30,86,31,176,31,36,31,36,30,161,31,161,30,251,31,251,30,74,31,195,31,195,30,6,31,186,31,186,30,186,29,157,31,160,31,23,31,190,31,223,31,141,31,141,30,224,31,224,30,54,31,245,31,245,30,62,31,225,31,225,30,225,29,30,31,30,30,207,31,84,31,145,31,154,31,233,31,18,31,116,31,116,30,207,31,139,31,139,30,22,31,164,31,126,31,82,31,176,31,153,31,147,31,134,31,134,30,192,31,229,31,9,31,124,31,40,31,105,31,231,31,190,31,118,31,118,30,30,31,239,31,148,31,148,30,248,31,137,31,137,30,209,31,209,30,116,31,66,31,200,31,178,31,178,30,255,31,28,31,224,31,107,31,85,31,24,31,8,31,8,30,201,31,169,31,169,30,130,31,209,31,211,31,135,31,135,30,135,29,4,31,156,31,156,30,77,31,88,31,185,31,153,31,196,31,146,31,128,31,146,31,146,30,146,29,246,31,182,31,225,31,213,31,102,31,52,31,138,31,138,30,194,31,82,31,48,31,48,30,182,31,150,31,28,31,243,31,243,30,180,31,222,31,102,31,102,30,102,29,10,31,223,31,210,31,68,31,199,31,171,31,102,31,211,31,183,31,170,31,210,31,142,31,18,31,231,31,107,31,1,31,38,31,38,30,38,29,38,28,121,31,73,31,73,30,183,31,183,30,227,31,133,31,117,31,77,31,87,31,87,30,87,29,87,28,133,31,189,31,242,31,7,31,101,31,101,30,101,29,25,31,53,31,215,31,205,31,212,31,49,31,225,31,249,31,226,31,244,31,12,31,94,31,137,31,229,31,20,31,132,31,216,31,216,30,72,31,231,31,69,31,69,30,69,29,11,31,202,31,115,31,208,31,200,31,135,31,202,31,202,30,83,31,154,31,248,31,177,31,177,30,45,31,40,31,218,31,218,30,106,31,106,30,115,31,78,31,78,30,78,29,208,31,231,31,217,31,84,31,182,31,192,31,11,31,9,31,244,31,63,31,71,31,186,31,191,31,83,31,12,31,43,31,43,30,7,31,3,31,141,31,148,31,37,31,37,30,23,31,253,31,114,31,114,30,55,31,84,31,84,30,208,31,121,31,233,31,233,30,205,31,17,31,22,31,8,31,8,30,70,31,187,31,183,31,19,31,19,30,77,31,77,30,220,31,220,30,224,31,113,31,76,31,1,31,1,30,1,29,228,31,154,31,248,31,248,30,79,31,249,31,131,31,130,31,86,31,11,31,215,31,20,31,50,31,50,30,240,31,15,31,146,31,241,31,229,31,185,31,185,30,217,31,67,31,144,31,99,31,99,30,99,29,29,31,13,31,42,31,252,31,118,31,44,31,210,31,210,30,210,29,69,31,122,31,84,31,52,31,113,31,148,31,177,31,165,31,165,30,254,31,254,30,136,31,154,31,154,30,164,31,30,31,231,31,118,31,118,30,118,29,25,31,85,31,70,31,151,31,70,31,107,31,107,30,134,31,64,31,64,30,24,31,38,31,79,31,200,31,82,31,66,31,95,31,202,31,202,30,6,31,62,31,95,31,149,31,137,31,174,31,25,31,162,31,162,30,209,31,209,30,111,31,221,31,35,31,220,31,119,31,68,31,10,31,21,31,19,31,159,31,78,31,208,31,221,31,239,31,172,31,34,31,121,31,45,31,133,31,98,31,95,31,39,31,206,31,206,30,232,31,8,31,199,31,243,31,41,31,41,30,212,31,212,30,212,29,201,31,130,31,114,31,231,31,231,30,39,31,39,30,191,31,191,30,37,31,184,31,103,31,197,31,59,31,32,31,32,30,173,31,47,31,49,31,225,31,27,31,70,31,49,31,227,31,185,31,107,31,89,31,119,31,159,31,159,30,20,31,110,31,131,31,135,31,156,31,112,31,177,31,187,31,84,31,234,31,50,31,202,31,202,30,195,31,237,31,237,30,237,29,213,31,109,31,54,31,217,31,217,30,206,31,116,31,5,31,182,31,25,31,166,31,106,31,95,31,95,30,95,29,44,31,44,30,153,31,252,31,252,30,20,31,20,30,56,31,110,31,87,31,128,31,179,31,147,31,147,30,93,31,221,31,232,31,209,31,41,31,9,31,176,31,168,31,82,31,101,31,11,31,156,31,156,30,196,31,252,31,167,31,126,31,24,31,143,31,189,31,50,31,131,31,131,30,102,31,132,31,91,31,88,31,101,31,220,31,223,31,223,30,206,31,103,31,204,31,204,30,222,31,245,31,223,31,202,31,150,31,150,30,150,29,150,28,63,31,159,31,121,31,24,31,24,30,206,31,222,31,95,31,150,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
