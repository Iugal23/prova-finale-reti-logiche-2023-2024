-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 826;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (50,0,251,0,147,0,160,0,98,0,8,0,96,0,53,0,213,0,148,0,181,0,136,0,0,0,185,0,124,0,240,0,198,0,0,0,0,0,193,0,90,0,32,0,55,0,51,0,0,0,84,0,0,0,244,0,0,0,0,0,102,0,115,0,142,0,0,0,93,0,77,0,21,0,247,0,170,0,143,0,23,0,245,0,0,0,0,0,207,0,27,0,18,0,28,0,67,0,0,0,63,0,21,0,102,0,0,0,0,0,96,0,201,0,204,0,85,0,0,0,80,0,0,0,173,0,232,0,248,0,166,0,0,0,0,0,209,0,156,0,225,0,92,0,52,0,100,0,103,0,248,0,237,0,89,0,45,0,204,0,191,0,190,0,208,0,249,0,0,0,0,0,89,0,0,0,135,0,136,0,110,0,241,0,140,0,194,0,148,0,77,0,154,0,86,0,0,0,152,0,28,0,90,0,79,0,0,0,250,0,0,0,0,0,125,0,152,0,0,0,0,0,58,0,59,0,255,0,0,0,35,0,0,0,44,0,175,0,0,0,0,0,0,0,207,0,1,0,201,0,110,0,38,0,109,0,80,0,11,0,120,0,0,0,0,0,0,0,63,0,0,0,0,0,157,0,251,0,23,0,203,0,160,0,177,0,0,0,23,0,31,0,0,0,0,0,0,0,133,0,27,0,41,0,100,0,0,0,1,0,98,0,38,0,164,0,210,0,49,0,110,0,130,0,224,0,200,0,225,0,0,0,90,0,120,0,65,0,101,0,240,0,180,0,161,0,254,0,172,0,0,0,26,0,238,0,102,0,21,0,0,0,12,0,40,0,0,0,223,0,173,0,73,0,44,0,0,0,0,0,0,0,155,0,176,0,228,0,98,0,33,0,135,0,172,0,124,0,180,0,90,0,87,0,0,0,42,0,185,0,0,0,2,0,133,0,21,0,131,0,92,0,115,0,0,0,0,0,51,0,157,0,224,0,243,0,216,0,209,0,108,0,148,0,152,0,236,0,0,0,167,0,69,0,47,0,102,0,64,0,73,0,0,0,205,0,86,0,135,0,247,0,24,0,0,0,0,0,68,0,247,0,60,0,0,0,0,0,0,0,184,0,172,0,0,0,12,0,0,0,224,0,250,0,251,0,18,0,34,0,17,0,206,0,163,0,221,0,0,0,0,0,141,0,94,0,216,0,38,0,138,0,171,0,0,0,226,0,191,0,62,0,0,0,0,0,102,0,14,0,132,0,54,0,162,0,229,0,14,0,15,0,169,0,0,0,12,0,69,0,75,0,52,0,240,0,154,0,183,0,202,0,77,0,125,0,61,0,231,0,26,0,116,0,199,0,0,0,48,0,0,0,60,0,0,0,96,0,64,0,78,0,214,0,0,0,3,0,183,0,0,0,253,0,34,0,160,0,70,0,242,0,140,0,144,0,227,0,173,0,246,0,166,0,206,0,92,0,8,0,197,0,192,0,131,0,0,0,151,0,123,0,126,0,79,0,13,0,0,0,0,0,19,0,65,0,246,0,47,0,138,0,245,0,163,0,25,0,0,0,214,0,81,0,45,0,148,0,95,0,126,0,240,0,35,0,169,0,87,0,191,0,191,0,55,0,129,0,187,0,61,0,235,0,214,0,0,0,143,0,18,0,208,0,1,0,203,0,94,0,105,0,239,0,203,0,128,0,131,0,197,0,107,0,107,0,75,0,0,0,198,0,0,0,0,0,84,0,108,0,0,0,187,0,16,0,228,0,244,0,17,0,50,0,77,0,177,0,10,0,79,0,205,0,215,0,39,0,83,0,205,0,117,0,149,0,14,0,210,0,35,0,64,0,0,0,59,0,81,0,0,0,124,0,12,0,0,0,0,0,218,0,22,0,0,0,0,0,216,0,156,0,93,0,101,0,246,0,229,0,0,0,0,0,40,0,224,0,116,0,184,0,42,0,11,0,0,0,80,0,0,0,151,0,179,0,237,0,33,0,120,0,142,0,62,0,0,0,161,0,86,0,232,0,0,0,190,0,209,0,253,0,0,0,74,0,9,0,111,0,0,0,18,0,0,0,250,0,0,0,213,0,134,0,164,0,0,0,110,0,165,0,223,0,0,0,23,0,204,0,161,0,0,0,61,0,118,0,194,0,0,0,138,0,87,0,36,0,51,0,187,0,97,0,229,0,229,0,0,0,0,0,0,0,103,0,0,0,245,0,0,0,0,0,0,0,162,0,113,0,209,0,0,0,232,0,0,0,0,0,214,0,253,0,249,0,0,0,0,0,21,0,40,0,58,0,227,0,133,0,193,0,125,0,218,0,101,0,146,0,0,0,0,0,50,0,0,0,54,0,0,0,0,0,0,0,10,0,0,0,200,0,0,0,0,0,49,0,106,0,0,0,249,0,16,0,177,0,236,0,14,0,242,0,119,0,0,0,0,0,0,0,85,0,213,0,6,0,145,0,0,0,31,0,133,0,192,0,0,0,241,0,120,0,0,0,170,0,13,0,123,0,196,0,135,0,154,0,238,0,139,0,185,0,129,0,170,0,145,0,223,0,0,0,79,0,7,0,154,0,33,0,0,0,0,0,79,0,121,0,62,0,0,0,0,0,234,0,68,0,15,0,112,0,82,0,130,0,0,0,189,0,227,0,154,0,141,0,19,0,0,0,232,0,2,0,0,0,103,0,147,0,98,0,0,0,19,0,0,0,33,0,82,0,142,0,91,0,0,0,192,0,46,0,48,0,0,0,196,0,169,0,29,0,195,0,87,0,206,0,0,0,4,0,228,0,231,0,213,0,160,0,142,0,4,0,0,0,12,0,0,0,55,0,0,0,154,0,142,0,153,0,248,0,107,0,100,0,161,0,128,0,0,0,160,0,222,0,0,0,161,0,69,0,58,0,199,0,2,0,0,0,191,0,196,0,0,0,227,0,194,0,73,0,156,0,174,0,28,0,69,0,60,0,229,0,65,0,155,0,0,0,182,0,104,0,0,0,105,0,213,0,32,0,44,0,0,0,65,0,147,0,117,0,23,0,242,0,0,0,71,0,5,0,83,0,241,0,185,0,0,0,150,0,59,0,10,0,235,0,0,0,28,0,176,0,0,0,0,0,208,0,53,0,11,0,13,0,85,0,0,0,136,0,103,0,246,0,198,0,124,0,233,0,135,0,112,0,43,0,139,0,143,0,0,0,199,0,161,0,50,0,0,0,49,0,148,0,126,0,118,0,93,0,117,0,0,0,239,0,0,0,35,0,189,0,163,0,144,0,159,0,195,0,0,0,183,0,104,0,127,0,0,0,74,0,252,0,123,0,0,0,0,0,6,0,228,0,225,0,217,0,0,0,155,0,102,0,202,0,163,0,83,0,142,0,0,0,169,0,255,0,10,0,42,0,151,0,0,0,0,0,85,0,147,0,178,0,47,0,66,0,94,0,0,0,235,0,144,0,0,0,65,0,160,0,238,0,135,0,0,0,27,0,241,0,24,0,142,0,20,0,0,0,0,0,0,0,135,0,207,0,0,0,193,0,145,0,151,0,0,0,191,0,0,0,46,0,178,0,0,0,252,0,213,0,85,0,184,0,81,0,0,0,0,0,76,0,168,0,158,0,221,0,0,0,226,0,92,0,155,0,223,0,0,0,213,0,159,0,0,0,82,0,69,0,0,0,88,0,0,0,188,0,125,0,204,0,12,0,254,0,140,0,199,0,6,0,207,0,55,0);
signal scenario_full  : scenario_type := (50,31,251,31,147,31,160,31,98,31,8,31,96,31,53,31,213,31,148,31,181,31,136,31,136,30,185,31,124,31,240,31,198,31,198,30,198,29,193,31,90,31,32,31,55,31,51,31,51,30,84,31,84,30,244,31,244,30,244,29,102,31,115,31,142,31,142,30,93,31,77,31,21,31,247,31,170,31,143,31,23,31,245,31,245,30,245,29,207,31,27,31,18,31,28,31,67,31,67,30,63,31,21,31,102,31,102,30,102,29,96,31,201,31,204,31,85,31,85,30,80,31,80,30,173,31,232,31,248,31,166,31,166,30,166,29,209,31,156,31,225,31,92,31,52,31,100,31,103,31,248,31,237,31,89,31,45,31,204,31,191,31,190,31,208,31,249,31,249,30,249,29,89,31,89,30,135,31,136,31,110,31,241,31,140,31,194,31,148,31,77,31,154,31,86,31,86,30,152,31,28,31,90,31,79,31,79,30,250,31,250,30,250,29,125,31,152,31,152,30,152,29,58,31,59,31,255,31,255,30,35,31,35,30,44,31,175,31,175,30,175,29,175,28,207,31,1,31,201,31,110,31,38,31,109,31,80,31,11,31,120,31,120,30,120,29,120,28,63,31,63,30,63,29,157,31,251,31,23,31,203,31,160,31,177,31,177,30,23,31,31,31,31,30,31,29,31,28,133,31,27,31,41,31,100,31,100,30,1,31,98,31,38,31,164,31,210,31,49,31,110,31,130,31,224,31,200,31,225,31,225,30,90,31,120,31,65,31,101,31,240,31,180,31,161,31,254,31,172,31,172,30,26,31,238,31,102,31,21,31,21,30,12,31,40,31,40,30,223,31,173,31,73,31,44,31,44,30,44,29,44,28,155,31,176,31,228,31,98,31,33,31,135,31,172,31,124,31,180,31,90,31,87,31,87,30,42,31,185,31,185,30,2,31,133,31,21,31,131,31,92,31,115,31,115,30,115,29,51,31,157,31,224,31,243,31,216,31,209,31,108,31,148,31,152,31,236,31,236,30,167,31,69,31,47,31,102,31,64,31,73,31,73,30,205,31,86,31,135,31,247,31,24,31,24,30,24,29,68,31,247,31,60,31,60,30,60,29,60,28,184,31,172,31,172,30,12,31,12,30,224,31,250,31,251,31,18,31,34,31,17,31,206,31,163,31,221,31,221,30,221,29,141,31,94,31,216,31,38,31,138,31,171,31,171,30,226,31,191,31,62,31,62,30,62,29,102,31,14,31,132,31,54,31,162,31,229,31,14,31,15,31,169,31,169,30,12,31,69,31,75,31,52,31,240,31,154,31,183,31,202,31,77,31,125,31,61,31,231,31,26,31,116,31,199,31,199,30,48,31,48,30,60,31,60,30,96,31,64,31,78,31,214,31,214,30,3,31,183,31,183,30,253,31,34,31,160,31,70,31,242,31,140,31,144,31,227,31,173,31,246,31,166,31,206,31,92,31,8,31,197,31,192,31,131,31,131,30,151,31,123,31,126,31,79,31,13,31,13,30,13,29,19,31,65,31,246,31,47,31,138,31,245,31,163,31,25,31,25,30,214,31,81,31,45,31,148,31,95,31,126,31,240,31,35,31,169,31,87,31,191,31,191,31,55,31,129,31,187,31,61,31,235,31,214,31,214,30,143,31,18,31,208,31,1,31,203,31,94,31,105,31,239,31,203,31,128,31,131,31,197,31,107,31,107,31,75,31,75,30,198,31,198,30,198,29,84,31,108,31,108,30,187,31,16,31,228,31,244,31,17,31,50,31,77,31,177,31,10,31,79,31,205,31,215,31,39,31,83,31,205,31,117,31,149,31,14,31,210,31,35,31,64,31,64,30,59,31,81,31,81,30,124,31,12,31,12,30,12,29,218,31,22,31,22,30,22,29,216,31,156,31,93,31,101,31,246,31,229,31,229,30,229,29,40,31,224,31,116,31,184,31,42,31,11,31,11,30,80,31,80,30,151,31,179,31,237,31,33,31,120,31,142,31,62,31,62,30,161,31,86,31,232,31,232,30,190,31,209,31,253,31,253,30,74,31,9,31,111,31,111,30,18,31,18,30,250,31,250,30,213,31,134,31,164,31,164,30,110,31,165,31,223,31,223,30,23,31,204,31,161,31,161,30,61,31,118,31,194,31,194,30,138,31,87,31,36,31,51,31,187,31,97,31,229,31,229,31,229,30,229,29,229,28,103,31,103,30,245,31,245,30,245,29,245,28,162,31,113,31,209,31,209,30,232,31,232,30,232,29,214,31,253,31,249,31,249,30,249,29,21,31,40,31,58,31,227,31,133,31,193,31,125,31,218,31,101,31,146,31,146,30,146,29,50,31,50,30,54,31,54,30,54,29,54,28,10,31,10,30,200,31,200,30,200,29,49,31,106,31,106,30,249,31,16,31,177,31,236,31,14,31,242,31,119,31,119,30,119,29,119,28,85,31,213,31,6,31,145,31,145,30,31,31,133,31,192,31,192,30,241,31,120,31,120,30,170,31,13,31,123,31,196,31,135,31,154,31,238,31,139,31,185,31,129,31,170,31,145,31,223,31,223,30,79,31,7,31,154,31,33,31,33,30,33,29,79,31,121,31,62,31,62,30,62,29,234,31,68,31,15,31,112,31,82,31,130,31,130,30,189,31,227,31,154,31,141,31,19,31,19,30,232,31,2,31,2,30,103,31,147,31,98,31,98,30,19,31,19,30,33,31,82,31,142,31,91,31,91,30,192,31,46,31,48,31,48,30,196,31,169,31,29,31,195,31,87,31,206,31,206,30,4,31,228,31,231,31,213,31,160,31,142,31,4,31,4,30,12,31,12,30,55,31,55,30,154,31,142,31,153,31,248,31,107,31,100,31,161,31,128,31,128,30,160,31,222,31,222,30,161,31,69,31,58,31,199,31,2,31,2,30,191,31,196,31,196,30,227,31,194,31,73,31,156,31,174,31,28,31,69,31,60,31,229,31,65,31,155,31,155,30,182,31,104,31,104,30,105,31,213,31,32,31,44,31,44,30,65,31,147,31,117,31,23,31,242,31,242,30,71,31,5,31,83,31,241,31,185,31,185,30,150,31,59,31,10,31,235,31,235,30,28,31,176,31,176,30,176,29,208,31,53,31,11,31,13,31,85,31,85,30,136,31,103,31,246,31,198,31,124,31,233,31,135,31,112,31,43,31,139,31,143,31,143,30,199,31,161,31,50,31,50,30,49,31,148,31,126,31,118,31,93,31,117,31,117,30,239,31,239,30,35,31,189,31,163,31,144,31,159,31,195,31,195,30,183,31,104,31,127,31,127,30,74,31,252,31,123,31,123,30,123,29,6,31,228,31,225,31,217,31,217,30,155,31,102,31,202,31,163,31,83,31,142,31,142,30,169,31,255,31,10,31,42,31,151,31,151,30,151,29,85,31,147,31,178,31,47,31,66,31,94,31,94,30,235,31,144,31,144,30,65,31,160,31,238,31,135,31,135,30,27,31,241,31,24,31,142,31,20,31,20,30,20,29,20,28,135,31,207,31,207,30,193,31,145,31,151,31,151,30,191,31,191,30,46,31,178,31,178,30,252,31,213,31,85,31,184,31,81,31,81,30,81,29,76,31,168,31,158,31,221,31,221,30,226,31,92,31,155,31,223,31,223,30,213,31,159,31,159,30,82,31,69,31,69,30,88,31,88,30,188,31,125,31,204,31,12,31,254,31,140,31,199,31,6,31,207,31,55,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
