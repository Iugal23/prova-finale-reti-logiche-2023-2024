-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_253 is
end project_tb_253;

architecture project_tb_arch_253 of project_tb_253 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 724;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (195,0,166,0,63,0,73,0,174,0,0,0,240,0,0,0,44,0,116,0,70,0,241,0,187,0,0,0,62,0,116,0,0,0,40,0,111,0,72,0,141,0,8,0,244,0,42,0,92,0,48,0,52,0,172,0,19,0,213,0,208,0,212,0,0,0,217,0,90,0,165,0,103,0,0,0,137,0,0,0,168,0,89,0,0,0,84,0,215,0,192,0,185,0,79,0,113,0,200,0,175,0,13,0,159,0,182,0,141,0,32,0,110,0,110,0,78,0,134,0,83,0,185,0,117,0,59,0,111,0,197,0,174,0,246,0,225,0,27,0,0,0,206,0,22,0,221,0,170,0,119,0,159,0,58,0,107,0,219,0,63,0,168,0,158,0,233,0,36,0,31,0,58,0,33,0,0,0,111,0,60,0,131,0,79,0,10,0,65,0,0,0,120,0,239,0,20,0,0,0,202,0,121,0,240,0,139,0,0,0,176,0,168,0,246,0,0,0,63,0,128,0,249,0,71,0,119,0,101,0,20,0,236,0,26,0,231,0,193,0,178,0,80,0,196,0,0,0,63,0,13,0,0,0,0,0,3,0,184,0,42,0,59,0,159,0,0,0,0,0,231,0,234,0,0,0,39,0,215,0,128,0,41,0,0,0,160,0,204,0,0,0,78,0,73,0,29,0,8,0,41,0,115,0,249,0,33,0,94,0,9,0,16,0,143,0,0,0,136,0,137,0,69,0,187,0,236,0,130,0,36,0,0,0,0,0,206,0,132,0,149,0,14,0,207,0,31,0,166,0,148,0,196,0,52,0,235,0,0,0,163,0,78,0,9,0,0,0,89,0,213,0,0,0,4,0,220,0,91,0,138,0,0,0,72,0,114,0,107,0,42,0,40,0,0,0,157,0,185,0,228,0,247,0,251,0,160,0,105,0,123,0,81,0,250,0,134,0,0,0,230,0,107,0,79,0,195,0,27,0,93,0,91,0,0,0,166,0,252,0,170,0,12,0,62,0,118,0,0,0,249,0,77,0,182,0,142,0,225,0,181,0,48,0,80,0,234,0,214,0,16,0,1,0,202,0,0,0,0,0,50,0,95,0,160,0,115,0,76,0,113,0,229,0,43,0,245,0,219,0,55,0,41,0,126,0,0,0,83,0,0,0,189,0,128,0,142,0,241,0,0,0,0,0,102,0,248,0,162,0,96,0,0,0,96,0,41,0,241,0,150,0,0,0,205,0,138,0,112,0,132,0,0,0,135,0,182,0,63,0,237,0,226,0,195,0,42,0,155,0,234,0,84,0,189,0,207,0,235,0,175,0,252,0,160,0,0,0,138,0,0,0,0,0,86,0,195,0,0,0,89,0,0,0,0,0,187,0,116,0,30,0,69,0,50,0,28,0,242,0,53,0,131,0,5,0,149,0,91,0,47,0,0,0,189,0,64,0,139,0,152,0,186,0,225,0,98,0,113,0,30,0,201,0,3,0,29,0,0,0,154,0,78,0,0,0,133,0,202,0,0,0,189,0,195,0,248,0,101,0,70,0,1,0,0,0,89,0,31,0,0,0,63,0,50,0,75,0,173,0,189,0,214,0,167,0,184,0,6,0,16,0,242,0,214,0,28,0,236,0,71,0,34,0,192,0,123,0,0,0,115,0,226,0,223,0,62,0,3,0,181,0,0,0,206,0,0,0,0,0,63,0,29,0,36,0,185,0,100,0,98,0,81,0,64,0,0,0,106,0,22,0,181,0,12,0,162,0,0,0,86,0,79,0,16,0,232,0,7,0,211,0,104,0,89,0,69,0,0,0,143,0,150,0,0,0,46,0,37,0,7,0,0,0,181,0,196,0,218,0,135,0,0,0,236,0,64,0,134,0,179,0,49,0,238,0,121,0,237,0,234,0,0,0,74,0,122,0,201,0,0,0,208,0,245,0,0,0,71,0,206,0,214,0,0,0,0,0,227,0,0,0,79,0,160,0,108,0,67,0,14,0,0,0,247,0,242,0,239,0,189,0,245,0,235,0,146,0,134,0,174,0,33,0,41,0,96,0,38,0,0,0,148,0,0,0,0,0,206,0,177,0,7,0,0,0,72,0,3,0,110,0,7,0,0,0,112,0,200,0,0,0,0,0,0,0,225,0,217,0,236,0,46,0,189,0,0,0,113,0,21,0,255,0,65,0,73,0,20,0,60,0,213,0,242,0,203,0,129,0,200,0,18,0,142,0,141,0,120,0,179,0,170,0,6,0,62,0,252,0,204,0,217,0,6,0,26,0,150,0,251,0,27,0,60,0,222,0,213,0,0,0,47,0,65,0,249,0,135,0,0,0,0,0,0,0,23,0,0,0,254,0,223,0,174,0,0,0,134,0,0,0,32,0,97,0,244,0,166,0,88,0,0,0,0,0,226,0,136,0,206,0,218,0,22,0,155,0,236,0,156,0,0,0,51,0,106,0,142,0,187,0,21,0,52,0,3,0,26,0,0,0,97,0,74,0,204,0,0,0,245,0,97,0,123,0,64,0,231,0,140,0,0,0,39,0,53,0,123,0,0,0,208,0,44,0,211,0,222,0,0,0,0,0,0,0,30,0,33,0,59,0,0,0,36,0,145,0,217,0,174,0,114,0,23,0,239,0,57,0,145,0,246,0,60,0,108,0,0,0,214,0,74,0,82,0,30,0,198,0,221,0,0,0,140,0,202,0,19,0,87,0,100,0,18,0,0,0,244,0,188,0,60,0,75,0,0,0,99,0,172,0,0,0,231,0,66,0,7,0,102,0,99,0,139,0,134,0,0,0,248,0,206,0,218,0,45,0,179,0,43,0,42,0,209,0,141,0,0,0,131,0,29,0,192,0,124,0,184,0,196,0,0,0,191,0,175,0,0,0,2,0,0,0,65,0,157,0,7,0,143,0,9,0,198,0,26,0,106,0,206,0,0,0,81,0,0,0,50,0,0,0,0,0,92,0,37,0,142,0,66,0,91,0,78,0,126,0,67,0,181,0,8,0,223,0,188,0,231,0,213,0,127,0,189,0,252,0,203,0,121,0,75,0,223,0,15,0,89,0,242,0,36,0,53,0,242,0,0,0,36,0,44,0,0,0,0,0,8,0,13,0,0,0,143,0,49,0,164,0,227,0,166,0,80,0,223,0,34,0,252,0,125,0,220,0,62,0,101,0,10,0,0,0,14,0,17,0,0,0,173,0,197,0,0,0,100,0,7,0,170,0,0,0,0,0,91,0,0,0,36,0,0,0,0,0,4,0);
signal scenario_full  : scenario_type := (195,31,166,31,63,31,73,31,174,31,174,30,240,31,240,30,44,31,116,31,70,31,241,31,187,31,187,30,62,31,116,31,116,30,40,31,111,31,72,31,141,31,8,31,244,31,42,31,92,31,48,31,52,31,172,31,19,31,213,31,208,31,212,31,212,30,217,31,90,31,165,31,103,31,103,30,137,31,137,30,168,31,89,31,89,30,84,31,215,31,192,31,185,31,79,31,113,31,200,31,175,31,13,31,159,31,182,31,141,31,32,31,110,31,110,31,78,31,134,31,83,31,185,31,117,31,59,31,111,31,197,31,174,31,246,31,225,31,27,31,27,30,206,31,22,31,221,31,170,31,119,31,159,31,58,31,107,31,219,31,63,31,168,31,158,31,233,31,36,31,31,31,58,31,33,31,33,30,111,31,60,31,131,31,79,31,10,31,65,31,65,30,120,31,239,31,20,31,20,30,202,31,121,31,240,31,139,31,139,30,176,31,168,31,246,31,246,30,63,31,128,31,249,31,71,31,119,31,101,31,20,31,236,31,26,31,231,31,193,31,178,31,80,31,196,31,196,30,63,31,13,31,13,30,13,29,3,31,184,31,42,31,59,31,159,31,159,30,159,29,231,31,234,31,234,30,39,31,215,31,128,31,41,31,41,30,160,31,204,31,204,30,78,31,73,31,29,31,8,31,41,31,115,31,249,31,33,31,94,31,9,31,16,31,143,31,143,30,136,31,137,31,69,31,187,31,236,31,130,31,36,31,36,30,36,29,206,31,132,31,149,31,14,31,207,31,31,31,166,31,148,31,196,31,52,31,235,31,235,30,163,31,78,31,9,31,9,30,89,31,213,31,213,30,4,31,220,31,91,31,138,31,138,30,72,31,114,31,107,31,42,31,40,31,40,30,157,31,185,31,228,31,247,31,251,31,160,31,105,31,123,31,81,31,250,31,134,31,134,30,230,31,107,31,79,31,195,31,27,31,93,31,91,31,91,30,166,31,252,31,170,31,12,31,62,31,118,31,118,30,249,31,77,31,182,31,142,31,225,31,181,31,48,31,80,31,234,31,214,31,16,31,1,31,202,31,202,30,202,29,50,31,95,31,160,31,115,31,76,31,113,31,229,31,43,31,245,31,219,31,55,31,41,31,126,31,126,30,83,31,83,30,189,31,128,31,142,31,241,31,241,30,241,29,102,31,248,31,162,31,96,31,96,30,96,31,41,31,241,31,150,31,150,30,205,31,138,31,112,31,132,31,132,30,135,31,182,31,63,31,237,31,226,31,195,31,42,31,155,31,234,31,84,31,189,31,207,31,235,31,175,31,252,31,160,31,160,30,138,31,138,30,138,29,86,31,195,31,195,30,89,31,89,30,89,29,187,31,116,31,30,31,69,31,50,31,28,31,242,31,53,31,131,31,5,31,149,31,91,31,47,31,47,30,189,31,64,31,139,31,152,31,186,31,225,31,98,31,113,31,30,31,201,31,3,31,29,31,29,30,154,31,78,31,78,30,133,31,202,31,202,30,189,31,195,31,248,31,101,31,70,31,1,31,1,30,89,31,31,31,31,30,63,31,50,31,75,31,173,31,189,31,214,31,167,31,184,31,6,31,16,31,242,31,214,31,28,31,236,31,71,31,34,31,192,31,123,31,123,30,115,31,226,31,223,31,62,31,3,31,181,31,181,30,206,31,206,30,206,29,63,31,29,31,36,31,185,31,100,31,98,31,81,31,64,31,64,30,106,31,22,31,181,31,12,31,162,31,162,30,86,31,79,31,16,31,232,31,7,31,211,31,104,31,89,31,69,31,69,30,143,31,150,31,150,30,46,31,37,31,7,31,7,30,181,31,196,31,218,31,135,31,135,30,236,31,64,31,134,31,179,31,49,31,238,31,121,31,237,31,234,31,234,30,74,31,122,31,201,31,201,30,208,31,245,31,245,30,71,31,206,31,214,31,214,30,214,29,227,31,227,30,79,31,160,31,108,31,67,31,14,31,14,30,247,31,242,31,239,31,189,31,245,31,235,31,146,31,134,31,174,31,33,31,41,31,96,31,38,31,38,30,148,31,148,30,148,29,206,31,177,31,7,31,7,30,72,31,3,31,110,31,7,31,7,30,112,31,200,31,200,30,200,29,200,28,225,31,217,31,236,31,46,31,189,31,189,30,113,31,21,31,255,31,65,31,73,31,20,31,60,31,213,31,242,31,203,31,129,31,200,31,18,31,142,31,141,31,120,31,179,31,170,31,6,31,62,31,252,31,204,31,217,31,6,31,26,31,150,31,251,31,27,31,60,31,222,31,213,31,213,30,47,31,65,31,249,31,135,31,135,30,135,29,135,28,23,31,23,30,254,31,223,31,174,31,174,30,134,31,134,30,32,31,97,31,244,31,166,31,88,31,88,30,88,29,226,31,136,31,206,31,218,31,22,31,155,31,236,31,156,31,156,30,51,31,106,31,142,31,187,31,21,31,52,31,3,31,26,31,26,30,97,31,74,31,204,31,204,30,245,31,97,31,123,31,64,31,231,31,140,31,140,30,39,31,53,31,123,31,123,30,208,31,44,31,211,31,222,31,222,30,222,29,222,28,30,31,33,31,59,31,59,30,36,31,145,31,217,31,174,31,114,31,23,31,239,31,57,31,145,31,246,31,60,31,108,31,108,30,214,31,74,31,82,31,30,31,198,31,221,31,221,30,140,31,202,31,19,31,87,31,100,31,18,31,18,30,244,31,188,31,60,31,75,31,75,30,99,31,172,31,172,30,231,31,66,31,7,31,102,31,99,31,139,31,134,31,134,30,248,31,206,31,218,31,45,31,179,31,43,31,42,31,209,31,141,31,141,30,131,31,29,31,192,31,124,31,184,31,196,31,196,30,191,31,175,31,175,30,2,31,2,30,65,31,157,31,7,31,143,31,9,31,198,31,26,31,106,31,206,31,206,30,81,31,81,30,50,31,50,30,50,29,92,31,37,31,142,31,66,31,91,31,78,31,126,31,67,31,181,31,8,31,223,31,188,31,231,31,213,31,127,31,189,31,252,31,203,31,121,31,75,31,223,31,15,31,89,31,242,31,36,31,53,31,242,31,242,30,36,31,44,31,44,30,44,29,8,31,13,31,13,30,143,31,49,31,164,31,227,31,166,31,80,31,223,31,34,31,252,31,125,31,220,31,62,31,101,31,10,31,10,30,14,31,17,31,17,30,173,31,197,31,197,30,100,31,7,31,170,31,170,30,170,29,91,31,91,30,36,31,36,30,36,29,4,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
