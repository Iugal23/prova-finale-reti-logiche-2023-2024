-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_400 is
end project_tb_400;

architecture project_tb_arch_400 of project_tb_400 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 773;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (193,0,60,0,41,0,242,0,120,0,183,0,0,0,0,0,138,0,53,0,1,0,180,0,0,0,0,0,144,0,34,0,120,0,192,0,235,0,45,0,39,0,142,0,0,0,131,0,24,0,251,0,49,0,135,0,154,0,108,0,0,0,235,0,0,0,89,0,50,0,142,0,49,0,66,0,77,0,105,0,100,0,127,0,34,0,191,0,54,0,14,0,162,0,203,0,0,0,178,0,178,0,81,0,69,0,1,0,15,0,123,0,185,0,250,0,48,0,0,0,80,0,57,0,205,0,109,0,0,0,190,0,0,0,51,0,82,0,133,0,200,0,195,0,196,0,168,0,0,0,165,0,45,0,84,0,74,0,38,0,0,0,87,0,174,0,175,0,129,0,86,0,40,0,0,0,26,0,0,0,1,0,22,0,0,0,215,0,33,0,0,0,99,0,12,0,29,0,0,0,0,0,18,0,40,0,254,0,0,0,132,0,185,0,155,0,0,0,17,0,21,0,0,0,146,0,130,0,0,0,164,0,247,0,248,0,116,0,39,0,47,0,0,0,218,0,221,0,221,0,32,0,212,0,0,0,76,0,223,0,227,0,0,0,217,0,181,0,234,0,3,0,133,0,87,0,0,0,98,0,88,0,10,0,108,0,126,0,108,0,185,0,24,0,134,0,85,0,125,0,0,0,69,0,0,0,205,0,247,0,0,0,225,0,1,0,228,0,14,0,204,0,219,0,229,0,2,0,144,0,188,0,0,0,150,0,200,0,195,0,113,0,0,0,77,0,118,0,0,0,169,0,0,0,0,0,189,0,0,0,162,0,33,0,224,0,0,0,10,0,105,0,125,0,82,0,0,0,100,0,0,0,53,0,0,0,36,0,0,0,238,0,25,0,152,0,0,0,243,0,91,0,177,0,0,0,51,0,0,0,229,0,0,0,197,0,123,0,26,0,201,0,127,0,92,0,95,0,218,0,0,0,174,0,34,0,63,0,0,0,228,0,116,0,0,0,105,0,177,0,0,0,184,0,65,0,200,0,88,0,129,0,81,0,252,0,21,0,195,0,0,0,91,0,0,0,31,0,235,0,234,0,242,0,0,0,219,0,130,0,0,0,99,0,57,0,0,0,175,0,0,0,163,0,247,0,210,0,0,0,251,0,0,0,77,0,233,0,221,0,6,0,0,0,0,0,9,0,0,0,106,0,138,0,0,0,19,0,34,0,0,0,116,0,20,0,169,0,240,0,93,0,0,0,0,0,30,0,228,0,130,0,184,0,137,0,0,0,0,0,157,0,0,0,17,0,84,0,253,0,144,0,189,0,84,0,170,0,34,0,32,0,0,0,0,0,27,0,69,0,251,0,175,0,163,0,0,0,251,0,28,0,31,0,245,0,47,0,177,0,208,0,121,0,0,0,244,0,244,0,252,0,90,0,115,0,134,0,0,0,178,0,44,0,245,0,135,0,0,0,240,0,177,0,225,0,0,0,21,0,186,0,107,0,0,0,0,0,91,0,158,0,0,0,0,0,14,0,229,0,34,0,236,0,111,0,248,0,0,0,51,0,0,0,53,0,0,0,229,0,0,0,20,0,214,0,37,0,0,0,54,0,177,0,5,0,93,0,58,0,0,0,246,0,57,0,90,0,92,0,2,0,227,0,0,0,212,0,201,0,56,0,247,0,198,0,27,0,0,0,0,0,211,0,0,0,41,0,110,0,174,0,224,0,235,0,0,0,0,0,207,0,127,0,0,0,43,0,204,0,196,0,126,0,0,0,170,0,17,0,91,0,39,0,173,0,0,0,9,0,61,0,208,0,84,0,0,0,164,0,0,0,0,0,0,0,246,0,237,0,8,0,0,0,122,0,33,0,246,0,0,0,25,0,0,0,214,0,82,0,154,0,0,0,108,0,180,0,83,0,251,0,0,0,28,0,80,0,0,0,90,0,254,0,72,0,31,0,159,0,163,0,29,0,156,0,37,0,14,0,233,0,142,0,0,0,149,0,190,0,70,0,52,0,109,0,196,0,97,0,151,0,140,0,0,0,108,0,153,0,229,0,0,0,162,0,239,0,17,0,0,0,223,0,24,0,0,0,251,0,86,0,0,0,121,0,79,0,0,0,146,0,130,0,237,0,130,0,184,0,219,0,0,0,82,0,211,0,109,0,93,0,0,0,136,0,211,0,211,0,0,0,14,0,0,0,246,0,30,0,160,0,147,0,183,0,0,0,0,0,118,0,162,0,59,0,230,0,111,0,97,0,24,0,246,0,237,0,164,0,118,0,241,0,21,0,0,0,224,0,168,0,0,0,39,0,0,0,0,0,244,0,146,0,135,0,252,0,239,0,151,0,211,0,96,0,0,0,151,0,226,0,71,0,1,0,48,0,16,0,71,0,254,0,0,0,183,0,212,0,132,0,0,0,185,0,42,0,79,0,145,0,0,0,82,0,92,0,89,0,195,0,232,0,3,0,58,0,39,0,195,0,150,0,32,0,0,0,218,0,24,0,128,0,28,0,114,0,86,0,0,0,0,0,139,0,57,0,90,0,206,0,163,0,0,0,83,0,193,0,114,0,233,0,11,0,196,0,0,0,123,0,116,0,126,0,218,0,43,0,57,0,185,0,166,0,160,0,217,0,35,0,112,0,210,0,0,0,59,0,217,0,205,0,101,0,247,0,0,0,83,0,0,0,188,0,89,0,188,0,38,0,205,0,0,0,6,0,213,0,232,0,219,0,158,0,0,0,0,0,61,0,243,0,248,0,162,0,120,0,196,0,174,0,188,0,250,0,5,0,101,0,199,0,234,0,124,0,9,0,0,0,162,0,48,0,252,0,166,0,0,0,127,0,184,0,119,0,132,0,196,0,247,0,20,0,182,0,0,0,0,0,132,0,52,0,108,0,114,0,214,0,0,0,0,0,0,0,79,0,50,0,206,0,249,0,0,0,0,0,0,0,18,0,0,0,0,0,147,0,42,0,0,0,178,0,0,0,85,0,214,0,217,0,85,0,118,0,199,0,0,0,143,0,158,0,19,0,213,0,157,0,236,0,158,0,16,0,9,0,182,0,56,0,138,0,236,0,31,0,101,0,71,0,185,0,57,0,227,0,158,0,0,0,98,0,100,0,111,0,187,0,6,0,78,0,116,0,37,0,144,0,144,0,100,0,253,0,179,0,0,0,203,0,99,0,0,0,200,0,72,0,53,0,0,0,210,0,120,0,0,0,154,0,74,0,53,0,47,0,0,0,0,0,0,0,146,0,253,0,202,0,192,0,97,0,246,0,126,0,108,0,167,0,119,0,1,0,81,0,131,0,0,0,199,0,0,0,54,0,82,0,242,0,0,0,222,0,132,0,114,0,46,0,187,0,0,0,255,0,240,0,16,0,143,0,0,0,0,0,126,0,72,0,189,0,119,0,48,0,23,0,77,0,172,0,0,0,194,0,192,0,187,0,0,0,55,0,213,0,204,0,77,0,26,0);
signal scenario_full  : scenario_type := (193,31,60,31,41,31,242,31,120,31,183,31,183,30,183,29,138,31,53,31,1,31,180,31,180,30,180,29,144,31,34,31,120,31,192,31,235,31,45,31,39,31,142,31,142,30,131,31,24,31,251,31,49,31,135,31,154,31,108,31,108,30,235,31,235,30,89,31,50,31,142,31,49,31,66,31,77,31,105,31,100,31,127,31,34,31,191,31,54,31,14,31,162,31,203,31,203,30,178,31,178,31,81,31,69,31,1,31,15,31,123,31,185,31,250,31,48,31,48,30,80,31,57,31,205,31,109,31,109,30,190,31,190,30,51,31,82,31,133,31,200,31,195,31,196,31,168,31,168,30,165,31,45,31,84,31,74,31,38,31,38,30,87,31,174,31,175,31,129,31,86,31,40,31,40,30,26,31,26,30,1,31,22,31,22,30,215,31,33,31,33,30,99,31,12,31,29,31,29,30,29,29,18,31,40,31,254,31,254,30,132,31,185,31,155,31,155,30,17,31,21,31,21,30,146,31,130,31,130,30,164,31,247,31,248,31,116,31,39,31,47,31,47,30,218,31,221,31,221,31,32,31,212,31,212,30,76,31,223,31,227,31,227,30,217,31,181,31,234,31,3,31,133,31,87,31,87,30,98,31,88,31,10,31,108,31,126,31,108,31,185,31,24,31,134,31,85,31,125,31,125,30,69,31,69,30,205,31,247,31,247,30,225,31,1,31,228,31,14,31,204,31,219,31,229,31,2,31,144,31,188,31,188,30,150,31,200,31,195,31,113,31,113,30,77,31,118,31,118,30,169,31,169,30,169,29,189,31,189,30,162,31,33,31,224,31,224,30,10,31,105,31,125,31,82,31,82,30,100,31,100,30,53,31,53,30,36,31,36,30,238,31,25,31,152,31,152,30,243,31,91,31,177,31,177,30,51,31,51,30,229,31,229,30,197,31,123,31,26,31,201,31,127,31,92,31,95,31,218,31,218,30,174,31,34,31,63,31,63,30,228,31,116,31,116,30,105,31,177,31,177,30,184,31,65,31,200,31,88,31,129,31,81,31,252,31,21,31,195,31,195,30,91,31,91,30,31,31,235,31,234,31,242,31,242,30,219,31,130,31,130,30,99,31,57,31,57,30,175,31,175,30,163,31,247,31,210,31,210,30,251,31,251,30,77,31,233,31,221,31,6,31,6,30,6,29,9,31,9,30,106,31,138,31,138,30,19,31,34,31,34,30,116,31,20,31,169,31,240,31,93,31,93,30,93,29,30,31,228,31,130,31,184,31,137,31,137,30,137,29,157,31,157,30,17,31,84,31,253,31,144,31,189,31,84,31,170,31,34,31,32,31,32,30,32,29,27,31,69,31,251,31,175,31,163,31,163,30,251,31,28,31,31,31,245,31,47,31,177,31,208,31,121,31,121,30,244,31,244,31,252,31,90,31,115,31,134,31,134,30,178,31,44,31,245,31,135,31,135,30,240,31,177,31,225,31,225,30,21,31,186,31,107,31,107,30,107,29,91,31,158,31,158,30,158,29,14,31,229,31,34,31,236,31,111,31,248,31,248,30,51,31,51,30,53,31,53,30,229,31,229,30,20,31,214,31,37,31,37,30,54,31,177,31,5,31,93,31,58,31,58,30,246,31,57,31,90,31,92,31,2,31,227,31,227,30,212,31,201,31,56,31,247,31,198,31,27,31,27,30,27,29,211,31,211,30,41,31,110,31,174,31,224,31,235,31,235,30,235,29,207,31,127,31,127,30,43,31,204,31,196,31,126,31,126,30,170,31,17,31,91,31,39,31,173,31,173,30,9,31,61,31,208,31,84,31,84,30,164,31,164,30,164,29,164,28,246,31,237,31,8,31,8,30,122,31,33,31,246,31,246,30,25,31,25,30,214,31,82,31,154,31,154,30,108,31,180,31,83,31,251,31,251,30,28,31,80,31,80,30,90,31,254,31,72,31,31,31,159,31,163,31,29,31,156,31,37,31,14,31,233,31,142,31,142,30,149,31,190,31,70,31,52,31,109,31,196,31,97,31,151,31,140,31,140,30,108,31,153,31,229,31,229,30,162,31,239,31,17,31,17,30,223,31,24,31,24,30,251,31,86,31,86,30,121,31,79,31,79,30,146,31,130,31,237,31,130,31,184,31,219,31,219,30,82,31,211,31,109,31,93,31,93,30,136,31,211,31,211,31,211,30,14,31,14,30,246,31,30,31,160,31,147,31,183,31,183,30,183,29,118,31,162,31,59,31,230,31,111,31,97,31,24,31,246,31,237,31,164,31,118,31,241,31,21,31,21,30,224,31,168,31,168,30,39,31,39,30,39,29,244,31,146,31,135,31,252,31,239,31,151,31,211,31,96,31,96,30,151,31,226,31,71,31,1,31,48,31,16,31,71,31,254,31,254,30,183,31,212,31,132,31,132,30,185,31,42,31,79,31,145,31,145,30,82,31,92,31,89,31,195,31,232,31,3,31,58,31,39,31,195,31,150,31,32,31,32,30,218,31,24,31,128,31,28,31,114,31,86,31,86,30,86,29,139,31,57,31,90,31,206,31,163,31,163,30,83,31,193,31,114,31,233,31,11,31,196,31,196,30,123,31,116,31,126,31,218,31,43,31,57,31,185,31,166,31,160,31,217,31,35,31,112,31,210,31,210,30,59,31,217,31,205,31,101,31,247,31,247,30,83,31,83,30,188,31,89,31,188,31,38,31,205,31,205,30,6,31,213,31,232,31,219,31,158,31,158,30,158,29,61,31,243,31,248,31,162,31,120,31,196,31,174,31,188,31,250,31,5,31,101,31,199,31,234,31,124,31,9,31,9,30,162,31,48,31,252,31,166,31,166,30,127,31,184,31,119,31,132,31,196,31,247,31,20,31,182,31,182,30,182,29,132,31,52,31,108,31,114,31,214,31,214,30,214,29,214,28,79,31,50,31,206,31,249,31,249,30,249,29,249,28,18,31,18,30,18,29,147,31,42,31,42,30,178,31,178,30,85,31,214,31,217,31,85,31,118,31,199,31,199,30,143,31,158,31,19,31,213,31,157,31,236,31,158,31,16,31,9,31,182,31,56,31,138,31,236,31,31,31,101,31,71,31,185,31,57,31,227,31,158,31,158,30,98,31,100,31,111,31,187,31,6,31,78,31,116,31,37,31,144,31,144,31,100,31,253,31,179,31,179,30,203,31,99,31,99,30,200,31,72,31,53,31,53,30,210,31,120,31,120,30,154,31,74,31,53,31,47,31,47,30,47,29,47,28,146,31,253,31,202,31,192,31,97,31,246,31,126,31,108,31,167,31,119,31,1,31,81,31,131,31,131,30,199,31,199,30,54,31,82,31,242,31,242,30,222,31,132,31,114,31,46,31,187,31,187,30,255,31,240,31,16,31,143,31,143,30,143,29,126,31,72,31,189,31,119,31,48,31,23,31,77,31,172,31,172,30,194,31,192,31,187,31,187,30,55,31,213,31,204,31,77,31,26,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
