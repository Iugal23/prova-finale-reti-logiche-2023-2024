-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 834;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (228,0,197,0,0,0,0,0,190,0,40,0,100,0,108,0,140,0,200,0,0,0,206,0,127,0,90,0,177,0,172,0,140,0,141,0,112,0,139,0,62,0,0,0,79,0,8,0,0,0,218,0,251,0,43,0,135,0,0,0,0,0,170,0,115,0,248,0,0,0,94,0,38,0,83,0,150,0,206,0,111,0,48,0,0,0,0,0,0,0,110,0,129,0,0,0,155,0,183,0,51,0,239,0,128,0,164,0,166,0,56,0,116,0,92,0,155,0,162,0,112,0,69,0,0,0,0,0,4,0,47,0,157,0,149,0,0,0,52,0,161,0,186,0,70,0,1,0,165,0,163,0,189,0,186,0,0,0,13,0,59,0,251,0,195,0,211,0,9,0,210,0,78,0,111,0,204,0,109,0,184,0,0,0,194,0,148,0,246,0,12,0,61,0,0,0,105,0,127,0,173,0,170,0,233,0,45,0,153,0,0,0,157,0,51,0,192,0,136,0,241,0,0,0,117,0,139,0,0,0,102,0,214,0,135,0,173,0,76,0,228,0,0,0,42,0,4,0,214,0,24,0,46,0,16,0,26,0,36,0,161,0,55,0,88,0,0,0,0,0,249,0,216,0,119,0,12,0,58,0,2,0,0,0,150,0,159,0,89,0,98,0,248,0,111,0,79,0,187,0,102,0,44,0,0,0,114,0,101,0,170,0,234,0,0,0,134,0,0,0,149,0,0,0,166,0,32,0,118,0,94,0,49,0,35,0,48,0,222,0,0,0,138,0,234,0,128,0,122,0,122,0,216,0,13,0,166,0,0,0,147,0,128,0,0,0,189,0,41,0,78,0,53,0,82,0,0,0,0,0,216,0,172,0,204,0,23,0,75,0,0,0,236,0,38,0,56,0,0,0,11,0,128,0,0,0,216,0,125,0,114,0,49,0,214,0,130,0,198,0,0,0,153,0,56,0,32,0,137,0,196,0,0,0,63,0,155,0,78,0,137,0,0,0,46,0,216,0,185,0,167,0,125,0,0,0,83,0,191,0,37,0,133,0,0,0,152,0,36,0,0,0,137,0,234,0,0,0,226,0,51,0,0,0,205,0,103,0,207,0,207,0,0,0,0,0,147,0,141,0,102,0,185,0,101,0,197,0,130,0,152,0,68,0,2,0,156,0,63,0,166,0,251,0,75,0,117,0,146,0,153,0,63,0,0,0,7,0,171,0,78,0,164,0,0,0,114,0,117,0,0,0,72,0,7,0,158,0,189,0,28,0,188,0,0,0,25,0,119,0,198,0,221,0,0,0,0,0,7,0,32,0,123,0,201,0,3,0,0,0,0,0,195,0,199,0,65,0,98,0,15,0,170,0,0,0,221,0,72,0,163,0,164,0,0,0,134,0,0,0,216,0,90,0,228,0,0,0,196,0,87,0,198,0,189,0,216,0,212,0,19,0,0,0,167,0,231,0,107,0,232,0,232,0,190,0,0,0,0,0,216,0,212,0,0,0,240,0,0,0,251,0,107,0,60,0,0,0,0,0,16,0,116,0,31,0,195,0,176,0,104,0,0,0,169,0,215,0,0,0,157,0,139,0,47,0,0,0,0,0,192,0,11,0,65,0,0,0,84,0,230,0,0,0,1,0,99,0,3,0,188,0,0,0,233,0,140,0,116,0,70,0,75,0,87,0,69,0,34,0,47,0,13,0,34,0,20,0,3,0,245,0,32,0,222,0,177,0,142,0,13,0,38,0,165,0,0,0,175,0,167,0,218,0,107,0,21,0,201,0,147,0,0,0,0,0,22,0,24,0,31,0,54,0,11,0,204,0,38,0,0,0,0,0,186,0,235,0,64,0,0,0,164,0,175,0,143,0,0,0,33,0,147,0,31,0,0,0,3,0,51,0,151,0,206,0,0,0,220,0,154,0,142,0,255,0,106,0,146,0,175,0,0,0,0,0,24,0,20,0,25,0,84,0,224,0,161,0,46,0,0,0,102,0,130,0,151,0,145,0,131,0,19,0,0,0,20,0,18,0,251,0,0,0,15,0,85,0,189,0,181,0,227,0,235,0,50,0,210,0,181,0,74,0,0,0,90,0,216,0,116,0,0,0,9,0,168,0,95,0,0,0,80,0,233,0,0,0,144,0,198,0,0,0,204,0,244,0,16,0,49,0,213,0,72,0,172,0,0,0,209,0,192,0,0,0,0,0,0,0,201,0,22,0,30,0,90,0,213,0,72,0,240,0,87,0,197,0,212,0,153,0,172,0,144,0,180,0,60,0,107,0,101,0,213,0,76,0,192,0,84,0,126,0,220,0,1,0,230,0,201,0,28,0,45,0,234,0,250,0,183,0,214,0,206,0,0,0,225,0,11,0,30,0,118,0,226,0,0,0,159,0,15,0,119,0,28,0,161,0,158,0,119,0,32,0,110,0,8,0,109,0,233,0,0,0,127,0,182,0,104,0,0,0,45,0,255,0,203,0,34,0,26,0,0,0,130,0,199,0,56,0,0,0,6,0,164,0,144,0,118,0,0,0,69,0,139,0,170,0,117,0,35,0,66,0,179,0,0,0,141,0,220,0,33,0,55,0,138,0,0,0,0,0,198,0,0,0,216,0,232,0,108,0,174,0,15,0,0,0,177,0,204,0,250,0,110,0,123,0,155,0,216,0,60,0,209,0,211,0,228,0,0,0,87,0,245,0,110,0,66,0,175,0,110,0,193,0,52,0,117,0,0,0,86,0,142,0,210,0,133,0,0,0,49,0,208,0,77,0,136,0,0,0,26,0,165,0,22,0,138,0,33,0,78,0,141,0,0,0,146,0,208,0,122,0,0,0,131,0,4,0,45,0,33,0,54,0,90,0,137,0,230,0,74,0,219,0,87,0,39,0,217,0,228,0,139,0,155,0,26,0,108,0,113,0,150,0,64,0,217,0,0,0,170,0,69,0,181,0,0,0,99,0,187,0,131,0,129,0,218,0,202,0,87,0,74,0,40,0,78,0,196,0,68,0,42,0,0,0,18,0,201,0,0,0,0,0,0,0,0,0,32,0,250,0,0,0,201,0,88,0,228,0,147,0,77,0,0,0,10,0,0,0,0,0,110,0,118,0,95,0,221,0,87,0,0,0,184,0,173,0,79,0,197,0,255,0,47,0,210,0,1,0,158,0,160,0,16,0,209,0,253,0,129,0,93,0,38,0,46,0,0,0,219,0,80,0,0,0,200,0,245,0,127,0,171,0,195,0,186,0,0,0,19,0,28,0,198,0,188,0,40,0,80,0,118,0,200,0,59,0,23,0,0,0,171,0,252,0,211,0,0,0,165,0,0,0,152,0,172,0,137,0,161,0,68,0,132,0,55,0,65,0,5,0,237,0,23,0,165,0,42,0,186,0,208,0,219,0,44,0,0,0,1,0,143,0,254,0,163,0,0,0,0,0,233,0,114,0,0,0,204,0,64,0,133,0,199,0,15,0,9,0,107,0,202,0,235,0,105,0,125,0,0,0,179,0,0,0,61,0,241,0,0,0,0,0,114,0,0,0,222,0,163,0,0,0,182,0,0,0,171,0,91,0,239,0,231,0,138,0,7,0,75,0,147,0,138,0,119,0,120,0,128,0,218,0,104,0,31,0,124,0,74,0,82,0,242,0,74,0,9,0,81,0,118,0,47,0,13,0,109,0,248,0,0,0,17,0,162,0,49,0,89,0,109,0,67,0,54,0,237,0,163,0,88,0,212,0,0,0,219,0,17,0,238,0);
signal scenario_full  : scenario_type := (228,31,197,31,197,30,197,29,190,31,40,31,100,31,108,31,140,31,200,31,200,30,206,31,127,31,90,31,177,31,172,31,140,31,141,31,112,31,139,31,62,31,62,30,79,31,8,31,8,30,218,31,251,31,43,31,135,31,135,30,135,29,170,31,115,31,248,31,248,30,94,31,38,31,83,31,150,31,206,31,111,31,48,31,48,30,48,29,48,28,110,31,129,31,129,30,155,31,183,31,51,31,239,31,128,31,164,31,166,31,56,31,116,31,92,31,155,31,162,31,112,31,69,31,69,30,69,29,4,31,47,31,157,31,149,31,149,30,52,31,161,31,186,31,70,31,1,31,165,31,163,31,189,31,186,31,186,30,13,31,59,31,251,31,195,31,211,31,9,31,210,31,78,31,111,31,204,31,109,31,184,31,184,30,194,31,148,31,246,31,12,31,61,31,61,30,105,31,127,31,173,31,170,31,233,31,45,31,153,31,153,30,157,31,51,31,192,31,136,31,241,31,241,30,117,31,139,31,139,30,102,31,214,31,135,31,173,31,76,31,228,31,228,30,42,31,4,31,214,31,24,31,46,31,16,31,26,31,36,31,161,31,55,31,88,31,88,30,88,29,249,31,216,31,119,31,12,31,58,31,2,31,2,30,150,31,159,31,89,31,98,31,248,31,111,31,79,31,187,31,102,31,44,31,44,30,114,31,101,31,170,31,234,31,234,30,134,31,134,30,149,31,149,30,166,31,32,31,118,31,94,31,49,31,35,31,48,31,222,31,222,30,138,31,234,31,128,31,122,31,122,31,216,31,13,31,166,31,166,30,147,31,128,31,128,30,189,31,41,31,78,31,53,31,82,31,82,30,82,29,216,31,172,31,204,31,23,31,75,31,75,30,236,31,38,31,56,31,56,30,11,31,128,31,128,30,216,31,125,31,114,31,49,31,214,31,130,31,198,31,198,30,153,31,56,31,32,31,137,31,196,31,196,30,63,31,155,31,78,31,137,31,137,30,46,31,216,31,185,31,167,31,125,31,125,30,83,31,191,31,37,31,133,31,133,30,152,31,36,31,36,30,137,31,234,31,234,30,226,31,51,31,51,30,205,31,103,31,207,31,207,31,207,30,207,29,147,31,141,31,102,31,185,31,101,31,197,31,130,31,152,31,68,31,2,31,156,31,63,31,166,31,251,31,75,31,117,31,146,31,153,31,63,31,63,30,7,31,171,31,78,31,164,31,164,30,114,31,117,31,117,30,72,31,7,31,158,31,189,31,28,31,188,31,188,30,25,31,119,31,198,31,221,31,221,30,221,29,7,31,32,31,123,31,201,31,3,31,3,30,3,29,195,31,199,31,65,31,98,31,15,31,170,31,170,30,221,31,72,31,163,31,164,31,164,30,134,31,134,30,216,31,90,31,228,31,228,30,196,31,87,31,198,31,189,31,216,31,212,31,19,31,19,30,167,31,231,31,107,31,232,31,232,31,190,31,190,30,190,29,216,31,212,31,212,30,240,31,240,30,251,31,107,31,60,31,60,30,60,29,16,31,116,31,31,31,195,31,176,31,104,31,104,30,169,31,215,31,215,30,157,31,139,31,47,31,47,30,47,29,192,31,11,31,65,31,65,30,84,31,230,31,230,30,1,31,99,31,3,31,188,31,188,30,233,31,140,31,116,31,70,31,75,31,87,31,69,31,34,31,47,31,13,31,34,31,20,31,3,31,245,31,32,31,222,31,177,31,142,31,13,31,38,31,165,31,165,30,175,31,167,31,218,31,107,31,21,31,201,31,147,31,147,30,147,29,22,31,24,31,31,31,54,31,11,31,204,31,38,31,38,30,38,29,186,31,235,31,64,31,64,30,164,31,175,31,143,31,143,30,33,31,147,31,31,31,31,30,3,31,51,31,151,31,206,31,206,30,220,31,154,31,142,31,255,31,106,31,146,31,175,31,175,30,175,29,24,31,20,31,25,31,84,31,224,31,161,31,46,31,46,30,102,31,130,31,151,31,145,31,131,31,19,31,19,30,20,31,18,31,251,31,251,30,15,31,85,31,189,31,181,31,227,31,235,31,50,31,210,31,181,31,74,31,74,30,90,31,216,31,116,31,116,30,9,31,168,31,95,31,95,30,80,31,233,31,233,30,144,31,198,31,198,30,204,31,244,31,16,31,49,31,213,31,72,31,172,31,172,30,209,31,192,31,192,30,192,29,192,28,201,31,22,31,30,31,90,31,213,31,72,31,240,31,87,31,197,31,212,31,153,31,172,31,144,31,180,31,60,31,107,31,101,31,213,31,76,31,192,31,84,31,126,31,220,31,1,31,230,31,201,31,28,31,45,31,234,31,250,31,183,31,214,31,206,31,206,30,225,31,11,31,30,31,118,31,226,31,226,30,159,31,15,31,119,31,28,31,161,31,158,31,119,31,32,31,110,31,8,31,109,31,233,31,233,30,127,31,182,31,104,31,104,30,45,31,255,31,203,31,34,31,26,31,26,30,130,31,199,31,56,31,56,30,6,31,164,31,144,31,118,31,118,30,69,31,139,31,170,31,117,31,35,31,66,31,179,31,179,30,141,31,220,31,33,31,55,31,138,31,138,30,138,29,198,31,198,30,216,31,232,31,108,31,174,31,15,31,15,30,177,31,204,31,250,31,110,31,123,31,155,31,216,31,60,31,209,31,211,31,228,31,228,30,87,31,245,31,110,31,66,31,175,31,110,31,193,31,52,31,117,31,117,30,86,31,142,31,210,31,133,31,133,30,49,31,208,31,77,31,136,31,136,30,26,31,165,31,22,31,138,31,33,31,78,31,141,31,141,30,146,31,208,31,122,31,122,30,131,31,4,31,45,31,33,31,54,31,90,31,137,31,230,31,74,31,219,31,87,31,39,31,217,31,228,31,139,31,155,31,26,31,108,31,113,31,150,31,64,31,217,31,217,30,170,31,69,31,181,31,181,30,99,31,187,31,131,31,129,31,218,31,202,31,87,31,74,31,40,31,78,31,196,31,68,31,42,31,42,30,18,31,201,31,201,30,201,29,201,28,201,27,32,31,250,31,250,30,201,31,88,31,228,31,147,31,77,31,77,30,10,31,10,30,10,29,110,31,118,31,95,31,221,31,87,31,87,30,184,31,173,31,79,31,197,31,255,31,47,31,210,31,1,31,158,31,160,31,16,31,209,31,253,31,129,31,93,31,38,31,46,31,46,30,219,31,80,31,80,30,200,31,245,31,127,31,171,31,195,31,186,31,186,30,19,31,28,31,198,31,188,31,40,31,80,31,118,31,200,31,59,31,23,31,23,30,171,31,252,31,211,31,211,30,165,31,165,30,152,31,172,31,137,31,161,31,68,31,132,31,55,31,65,31,5,31,237,31,23,31,165,31,42,31,186,31,208,31,219,31,44,31,44,30,1,31,143,31,254,31,163,31,163,30,163,29,233,31,114,31,114,30,204,31,64,31,133,31,199,31,15,31,9,31,107,31,202,31,235,31,105,31,125,31,125,30,179,31,179,30,61,31,241,31,241,30,241,29,114,31,114,30,222,31,163,31,163,30,182,31,182,30,171,31,91,31,239,31,231,31,138,31,7,31,75,31,147,31,138,31,119,31,120,31,128,31,218,31,104,31,31,31,124,31,74,31,82,31,242,31,74,31,9,31,81,31,118,31,47,31,13,31,109,31,248,31,248,30,17,31,162,31,49,31,89,31,109,31,67,31,54,31,237,31,163,31,88,31,212,31,212,30,219,31,17,31,238,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
