-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 830;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (7,0,41,0,160,0,0,0,12,0,99,0,68,0,226,0,127,0,133,0,103,0,205,0,102,0,234,0,50,0,104,0,131,0,74,0,0,0,97,0,6,0,134,0,3,0,238,0,11,0,211,0,240,0,43,0,25,0,127,0,26,0,0,0,201,0,150,0,0,0,0,0,0,0,232,0,182,0,0,0,46,0,88,0,244,0,235,0,21,0,19,0,53,0,144,0,220,0,140,0,0,0,117,0,205,0,0,0,5,0,0,0,252,0,165,0,141,0,42,0,98,0,0,0,134,0,182,0,0,0,72,0,139,0,168,0,121,0,239,0,124,0,148,0,170,0,91,0,101,0,0,0,213,0,44,0,200,0,186,0,206,0,68,0,0,0,140,0,215,0,251,0,178,0,140,0,44,0,175,0,9,0,45,0,0,0,4,0,150,0,83,0,6,0,7,0,173,0,64,0,94,0,94,0,199,0,10,0,238,0,53,0,197,0,62,0,0,0,214,0,248,0,27,0,85,0,189,0,121,0,158,0,120,0,0,0,66,0,98,0,0,0,0,0,234,0,108,0,196,0,167,0,217,0,212,0,33,0,0,0,128,0,0,0,79,0,62,0,44,0,192,0,12,0,61,0,133,0,119,0,48,0,231,0,102,0,112,0,0,0,85,0,140,0,87,0,139,0,194,0,197,0,225,0,11,0,128,0,193,0,9,0,47,0,40,0,19,0,171,0,145,0,96,0,50,0,68,0,20,0,0,0,146,0,41,0,15,0,27,0,0,0,0,0,35,0,163,0,0,0,133,0,165,0,246,0,0,0,244,0,87,0,62,0,91,0,82,0,172,0,59,0,193,0,243,0,0,0,0,0,196,0,0,0,15,0,255,0,222,0,91,0,202,0,118,0,150,0,177,0,175,0,145,0,108,0,130,0,189,0,197,0,58,0,169,0,87,0,235,0,178,0,0,0,15,0,93,0,114,0,10,0,27,0,51,0,93,0,0,0,254,0,3,0,0,0,56,0,51,0,252,0,211,0,247,0,0,0,175,0,122,0,252,0,0,0,138,0,0,0,148,0,0,0,127,0,166,0,104,0,24,0,0,0,219,0,46,0,6,0,47,0,126,0,0,0,7,0,92,0,68,0,114,0,52,0,50,0,141,0,104,0,70,0,38,0,189,0,117,0,73,0,248,0,0,0,73,0,75,0,150,0,0,0,54,0,110,0,244,0,100,0,93,0,58,0,194,0,0,0,252,0,218,0,153,0,154,0,106,0,171,0,78,0,145,0,0,0,78,0,158,0,0,0,60,0,20,0,245,0,243,0,23,0,0,0,181,0,68,0,215,0,48,0,255,0,0,0,204,0,238,0,146,0,236,0,37,0,221,0,27,0,55,0,65,0,151,0,0,0,168,0,99,0,74,0,205,0,148,0,0,0,195,0,0,0,0,0,0,0,199,0,237,0,0,0,0,0,207,0,70,0,25,0,249,0,143,0,0,0,253,0,242,0,54,0,24,0,11,0,125,0,170,0,197,0,137,0,61,0,0,0,193,0,139,0,144,0,161,0,0,0,34,0,161,0,192,0,174,0,213,0,63,0,0,0,57,0,137,0,197,0,38,0,155,0,238,0,214,0,172,0,172,0,9,0,59,0,191,0,168,0,224,0,231,0,26,0,52,0,0,0,129,0,145,0,108,0,130,0,214,0,0,0,0,0,53,0,18,0,139,0,240,0,0,0,119,0,129,0,16,0,191,0,165,0,0,0,0,0,19,0,39,0,156,0,228,0,90,0,47,0,6,0,151,0,0,0,0,0,40,0,0,0,45,0,153,0,210,0,96,0,21,0,0,0,139,0,25,0,35,0,199,0,28,0,83,0,134,0,182,0,142,0,34,0,81,0,118,0,75,0,228,0,171,0,90,0,0,0,193,0,146,0,126,0,242,0,197,0,0,0,132,0,42,0,1,0,137,0,164,0,230,0,236,0,0,0,1,0,150,0,128,0,250,0,247,0,127,0,0,0,188,0,0,0,233,0,190,0,0,0,73,0,145,0,0,0,208,0,147,0,103,0,83,0,1,0,0,0,11,0,100,0,49,0,239,0,222,0,77,0,21,0,1,0,118,0,10,0,28,0,29,0,24,0,14,0,254,0,0,0,33,0,133,0,118,0,0,0,85,0,0,0,26,0,58,0,120,0,0,0,21,0,75,0,0,0,92,0,0,0,101,0,187,0,0,0,0,0,64,0,87,0,0,0,133,0,0,0,152,0,230,0,0,0,0,0,238,0,187,0,0,0,12,0,210,0,125,0,0,0,222,0,195,0,144,0,168,0,214,0,168,0,213,0,151,0,39,0,243,0,70,0,208,0,0,0,0,0,187,0,149,0,0,0,137,0,214,0,164,0,124,0,49,0,145,0,255,0,48,0,222,0,0,0,148,0,0,0,102,0,132,0,100,0,161,0,127,0,183,0,0,0,139,0,10,0,52,0,115,0,202,0,205,0,170,0,200,0,166,0,255,0,8,0,47,0,240,0,20,0,57,0,100,0,7,0,217,0,165,0,252,0,13,0,6,0,148,0,129,0,13,0,80,0,64,0,87,0,172,0,12,0,0,0,26,0,95,0,226,0,0,0,0,0,170,0,2,0,13,0,0,0,165,0,201,0,1,0,133,0,233,0,156,0,50,0,157,0,60,0,39,0,120,0,226,0,222,0,0,0,212,0,131,0,113,0,0,0,136,0,242,0,75,0,130,0,224,0,118,0,199,0,79,0,74,0,73,0,250,0,28,0,192,0,0,0,56,0,247,0,67,0,45,0,74,0,89,0,0,0,185,0,0,0,0,0,169,0,86,0,186,0,196,0,0,0,200,0,211,0,159,0,113,0,164,0,137,0,23,0,88,0,212,0,255,0,180,0,130,0,137,0,158,0,0,0,79,0,132,0,156,0,169,0,0,0,0,0,236,0,128,0,0,0,0,0,98,0,26,0,5,0,251,0,63,0,0,0,186,0,0,0,104,0,209,0,156,0,85,0,222,0,0,0,137,0,0,0,0,0,120,0,0,0,231,0,0,0,38,0,0,0,0,0,88,0,37,0,83,0,26,0,69,0,213,0,25,0,218,0,0,0,96,0,219,0,146,0,161,0,140,0,0,0,0,0,0,0,137,0,173,0,228,0,77,0,87,0,46,0,42,0,99,0,206,0,68,0,128,0,97,0,214,0,130,0,224,0,134,0,53,0,58,0,0,0,164,0,200,0,147,0,0,0,0,0,90,0,143,0,226,0,90,0,149,0,237,0,0,0,93,0,58,0,0,0,70,0,107,0,224,0,178,0,103,0,37,0,139,0,198,0,232,0,0,0,185,0,86,0,33,0,1,0,226,0,18,0,193,0,126,0,0,0,198,0,89,0,161,0,252,0,48,0,0,0,236,0,250,0,227,0,239,0,102,0,209,0,0,0,20,0,37,0,132,0,45,0,3,0,93,0,102,0,0,0,191,0,0,0,78,0,201,0,243,0,68,0,108,0,38,0,123,0,136,0,79,0,33,0,142,0,163,0,51,0,77,0,237,0,116,0,34,0,100,0,179,0,158,0,152,0,134,0,194,0,213,0,8,0,10,0,232,0,127,0,110,0,229,0,218,0,183,0,133,0,3,0,0,0,111,0,162,0,0,0,127,0,0,0,0,0,0,0,0,0,253,0,55,0,5,0,0,0,176,0,33,0,194,0,0,0,0,0,98,0,82,0);
signal scenario_full  : scenario_type := (7,31,41,31,160,31,160,30,12,31,99,31,68,31,226,31,127,31,133,31,103,31,205,31,102,31,234,31,50,31,104,31,131,31,74,31,74,30,97,31,6,31,134,31,3,31,238,31,11,31,211,31,240,31,43,31,25,31,127,31,26,31,26,30,201,31,150,31,150,30,150,29,150,28,232,31,182,31,182,30,46,31,88,31,244,31,235,31,21,31,19,31,53,31,144,31,220,31,140,31,140,30,117,31,205,31,205,30,5,31,5,30,252,31,165,31,141,31,42,31,98,31,98,30,134,31,182,31,182,30,72,31,139,31,168,31,121,31,239,31,124,31,148,31,170,31,91,31,101,31,101,30,213,31,44,31,200,31,186,31,206,31,68,31,68,30,140,31,215,31,251,31,178,31,140,31,44,31,175,31,9,31,45,31,45,30,4,31,150,31,83,31,6,31,7,31,173,31,64,31,94,31,94,31,199,31,10,31,238,31,53,31,197,31,62,31,62,30,214,31,248,31,27,31,85,31,189,31,121,31,158,31,120,31,120,30,66,31,98,31,98,30,98,29,234,31,108,31,196,31,167,31,217,31,212,31,33,31,33,30,128,31,128,30,79,31,62,31,44,31,192,31,12,31,61,31,133,31,119,31,48,31,231,31,102,31,112,31,112,30,85,31,140,31,87,31,139,31,194,31,197,31,225,31,11,31,128,31,193,31,9,31,47,31,40,31,19,31,171,31,145,31,96,31,50,31,68,31,20,31,20,30,146,31,41,31,15,31,27,31,27,30,27,29,35,31,163,31,163,30,133,31,165,31,246,31,246,30,244,31,87,31,62,31,91,31,82,31,172,31,59,31,193,31,243,31,243,30,243,29,196,31,196,30,15,31,255,31,222,31,91,31,202,31,118,31,150,31,177,31,175,31,145,31,108,31,130,31,189,31,197,31,58,31,169,31,87,31,235,31,178,31,178,30,15,31,93,31,114,31,10,31,27,31,51,31,93,31,93,30,254,31,3,31,3,30,56,31,51,31,252,31,211,31,247,31,247,30,175,31,122,31,252,31,252,30,138,31,138,30,148,31,148,30,127,31,166,31,104,31,24,31,24,30,219,31,46,31,6,31,47,31,126,31,126,30,7,31,92,31,68,31,114,31,52,31,50,31,141,31,104,31,70,31,38,31,189,31,117,31,73,31,248,31,248,30,73,31,75,31,150,31,150,30,54,31,110,31,244,31,100,31,93,31,58,31,194,31,194,30,252,31,218,31,153,31,154,31,106,31,171,31,78,31,145,31,145,30,78,31,158,31,158,30,60,31,20,31,245,31,243,31,23,31,23,30,181,31,68,31,215,31,48,31,255,31,255,30,204,31,238,31,146,31,236,31,37,31,221,31,27,31,55,31,65,31,151,31,151,30,168,31,99,31,74,31,205,31,148,31,148,30,195,31,195,30,195,29,195,28,199,31,237,31,237,30,237,29,207,31,70,31,25,31,249,31,143,31,143,30,253,31,242,31,54,31,24,31,11,31,125,31,170,31,197,31,137,31,61,31,61,30,193,31,139,31,144,31,161,31,161,30,34,31,161,31,192,31,174,31,213,31,63,31,63,30,57,31,137,31,197,31,38,31,155,31,238,31,214,31,172,31,172,31,9,31,59,31,191,31,168,31,224,31,231,31,26,31,52,31,52,30,129,31,145,31,108,31,130,31,214,31,214,30,214,29,53,31,18,31,139,31,240,31,240,30,119,31,129,31,16,31,191,31,165,31,165,30,165,29,19,31,39,31,156,31,228,31,90,31,47,31,6,31,151,31,151,30,151,29,40,31,40,30,45,31,153,31,210,31,96,31,21,31,21,30,139,31,25,31,35,31,199,31,28,31,83,31,134,31,182,31,142,31,34,31,81,31,118,31,75,31,228,31,171,31,90,31,90,30,193,31,146,31,126,31,242,31,197,31,197,30,132,31,42,31,1,31,137,31,164,31,230,31,236,31,236,30,1,31,150,31,128,31,250,31,247,31,127,31,127,30,188,31,188,30,233,31,190,31,190,30,73,31,145,31,145,30,208,31,147,31,103,31,83,31,1,31,1,30,11,31,100,31,49,31,239,31,222,31,77,31,21,31,1,31,118,31,10,31,28,31,29,31,24,31,14,31,254,31,254,30,33,31,133,31,118,31,118,30,85,31,85,30,26,31,58,31,120,31,120,30,21,31,75,31,75,30,92,31,92,30,101,31,187,31,187,30,187,29,64,31,87,31,87,30,133,31,133,30,152,31,230,31,230,30,230,29,238,31,187,31,187,30,12,31,210,31,125,31,125,30,222,31,195,31,144,31,168,31,214,31,168,31,213,31,151,31,39,31,243,31,70,31,208,31,208,30,208,29,187,31,149,31,149,30,137,31,214,31,164,31,124,31,49,31,145,31,255,31,48,31,222,31,222,30,148,31,148,30,102,31,132,31,100,31,161,31,127,31,183,31,183,30,139,31,10,31,52,31,115,31,202,31,205,31,170,31,200,31,166,31,255,31,8,31,47,31,240,31,20,31,57,31,100,31,7,31,217,31,165,31,252,31,13,31,6,31,148,31,129,31,13,31,80,31,64,31,87,31,172,31,12,31,12,30,26,31,95,31,226,31,226,30,226,29,170,31,2,31,13,31,13,30,165,31,201,31,1,31,133,31,233,31,156,31,50,31,157,31,60,31,39,31,120,31,226,31,222,31,222,30,212,31,131,31,113,31,113,30,136,31,242,31,75,31,130,31,224,31,118,31,199,31,79,31,74,31,73,31,250,31,28,31,192,31,192,30,56,31,247,31,67,31,45,31,74,31,89,31,89,30,185,31,185,30,185,29,169,31,86,31,186,31,196,31,196,30,200,31,211,31,159,31,113,31,164,31,137,31,23,31,88,31,212,31,255,31,180,31,130,31,137,31,158,31,158,30,79,31,132,31,156,31,169,31,169,30,169,29,236,31,128,31,128,30,128,29,98,31,26,31,5,31,251,31,63,31,63,30,186,31,186,30,104,31,209,31,156,31,85,31,222,31,222,30,137,31,137,30,137,29,120,31,120,30,231,31,231,30,38,31,38,30,38,29,88,31,37,31,83,31,26,31,69,31,213,31,25,31,218,31,218,30,96,31,219,31,146,31,161,31,140,31,140,30,140,29,140,28,137,31,173,31,228,31,77,31,87,31,46,31,42,31,99,31,206,31,68,31,128,31,97,31,214,31,130,31,224,31,134,31,53,31,58,31,58,30,164,31,200,31,147,31,147,30,147,29,90,31,143,31,226,31,90,31,149,31,237,31,237,30,93,31,58,31,58,30,70,31,107,31,224,31,178,31,103,31,37,31,139,31,198,31,232,31,232,30,185,31,86,31,33,31,1,31,226,31,18,31,193,31,126,31,126,30,198,31,89,31,161,31,252,31,48,31,48,30,236,31,250,31,227,31,239,31,102,31,209,31,209,30,20,31,37,31,132,31,45,31,3,31,93,31,102,31,102,30,191,31,191,30,78,31,201,31,243,31,68,31,108,31,38,31,123,31,136,31,79,31,33,31,142,31,163,31,51,31,77,31,237,31,116,31,34,31,100,31,179,31,158,31,152,31,134,31,194,31,213,31,8,31,10,31,232,31,127,31,110,31,229,31,218,31,183,31,133,31,3,31,3,30,111,31,162,31,162,30,127,31,127,30,127,29,127,28,127,27,253,31,55,31,5,31,5,30,176,31,33,31,194,31,194,30,194,29,98,31,82,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
