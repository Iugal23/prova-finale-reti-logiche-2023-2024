-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_829 is
end project_tb_829;

architecture project_tb_arch_829 of project_tb_829 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 732;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (138,0,96,0,0,0,138,0,0,0,207,0,192,0,221,0,194,0,94,0,115,0,86,0,197,0,150,0,0,0,96,0,220,0,42,0,0,0,184,0,15,0,236,0,177,0,102,0,0,0,135,0,69,0,26,0,0,0,0,0,210,0,147,0,251,0,95,0,165,0,17,0,53,0,179,0,122,0,83,0,14,0,0,0,18,0,180,0,158,0,101,0,57,0,197,0,0,0,33,0,125,0,40,0,255,0,0,0,3,0,82,0,0,0,67,0,240,0,218,0,219,0,248,0,3,0,0,0,0,0,254,0,222,0,215,0,196,0,0,0,0,0,0,0,0,0,232,0,56,0,5,0,92,0,32,0,65,0,140,0,157,0,133,0,153,0,176,0,137,0,60,0,0,0,0,0,32,0,209,0,76,0,121,0,0,0,191,0,145,0,132,0,206,0,57,0,31,0,7,0,238,0,0,0,108,0,59,0,159,0,60,0,129,0,117,0,178,0,32,0,222,0,179,0,221,0,178,0,0,0,185,0,95,0,1,0,170,0,127,0,90,0,25,0,91,0,136,0,140,0,79,0,81,0,0,0,47,0,226,0,191,0,0,0,239,0,160,0,248,0,0,0,107,0,224,0,85,0,248,0,0,0,132,0,0,0,0,0,137,0,160,0,107,0,223,0,0,0,243,0,0,0,46,0,0,0,172,0,171,0,206,0,198,0,0,0,127,0,173,0,9,0,73,0,16,0,0,0,92,0,7,0,11,0,0,0,38,0,56,0,218,0,67,0,94,0,34,0,0,0,184,0,29,0,148,0,127,0,70,0,26,0,229,0,184,0,173,0,113,0,158,0,212,0,130,0,89,0,44,0,179,0,0,0,197,0,0,0,0,0,169,0,128,0,0,0,188,0,0,0,246,0,0,0,127,0,138,0,0,0,211,0,111,0,29,0,48,0,166,0,216,0,16,0,0,0,218,0,40,0,0,0,13,0,196,0,114,0,0,0,99,0,115,0,20,0,93,0,170,0,0,0,101,0,154,0,34,0,0,0,0,0,0,0,0,0,202,0,230,0,0,0,0,0,59,0,0,0,25,0,246,0,162,0,89,0,108,0,101,0,3,0,0,0,22,0,28,0,183,0,199,0,135,0,133,0,77,0,159,0,88,0,219,0,165,0,131,0,27,0,168,0,0,0,235,0,204,0,0,0,179,0,168,0,64,0,150,0,0,0,0,0,102,0,23,0,169,0,15,0,0,0,175,0,242,0,28,0,180,0,115,0,83,0,0,0,160,0,62,0,4,0,200,0,149,0,6,0,202,0,128,0,182,0,104,0,118,0,20,0,254,0,15,0,54,0,73,0,1,0,0,0,156,0,230,0,67,0,114,0,145,0,39,0,251,0,0,0,149,0,0,0,0,0,0,0,89,0,248,0,0,0,173,0,162,0,186,0,253,0,142,0,194,0,235,0,3,0,236,0,178,0,191,0,29,0,117,0,151,0,233,0,185,0,0,0,70,0,129,0,157,0,247,0,60,0,73,0,196,0,187,0,0,0,235,0,0,0,46,0,72,0,42,0,226,0,63,0,0,0,71,0,198,0,8,0,167,0,49,0,150,0,202,0,129,0,0,0,248,0,109,0,255,0,201,0,0,0,251,0,126,0,142,0,66,0,222,0,122,0,176,0,185,0,252,0,208,0,122,0,0,0,16,0,84,0,19,0,0,0,102,0,170,0,168,0,29,0,0,0,0,0,13,0,19,0,246,0,154,0,163,0,0,0,57,0,14,0,121,0,0,0,183,0,147,0,0,0,211,0,128,0,247,0,69,0,117,0,138,0,115,0,0,0,90,0,173,0,229,0,45,0,139,0,0,0,102,0,0,0,96,0,12,0,73,0,101,0,191,0,15,0,107,0,204,0,181,0,138,0,83,0,48,0,0,0,233,0,25,0,244,0,29,0,34,0,0,0,191,0,0,0,246,0,208,0,129,0,0,0,169,0,182,0,195,0,174,0,127,0,103,0,115,0,176,0,35,0,239,0,30,0,101,0,114,0,0,0,104,0,0,0,0,0,144,0,248,0,171,0,0,0,249,0,88,0,40,0,170,0,194,0,102,0,0,0,97,0,44,0,175,0,171,0,183,0,188,0,0,0,226,0,52,0,209,0,188,0,123,0,0,0,0,0,0,0,0,0,0,0,17,0,18,0,250,0,125,0,158,0,152,0,0,0,145,0,206,0,115,0,205,0,0,0,6,0,239,0,78,0,176,0,212,0,0,0,65,0,53,0,43,0,0,0,189,0,0,0,130,0,193,0,0,0,0,0,148,0,54,0,85,0,0,0,198,0,167,0,0,0,98,0,20,0,239,0,91,0,121,0,130,0,228,0,213,0,214,0,0,0,38,0,84,0,0,0,122,0,2,0,79,0,127,0,122,0,26,0,0,0,0,0,226,0,99,0,80,0,165,0,0,0,0,0,0,0,38,0,124,0,212,0,161,0,163,0,3,0,163,0,103,0,142,0,170,0,250,0,245,0,142,0,226,0,172,0,204,0,124,0,117,0,91,0,82,0,252,0,216,0,251,0,241,0,200,0,253,0,84,0,0,0,56,0,249,0,0,0,28,0,244,0,105,0,186,0,166,0,151,0,106,0,157,0,0,0,230,0,127,0,235,0,52,0,138,0,46,0,71,0,227,0,180,0,109,0,147,0,33,0,218,0,0,0,165,0,128,0,0,0,67,0,61,0,0,0,116,0,67,0,66,0,49,0,0,0,0,0,214,0,0,0,0,0,5,0,78,0,80,0,192,0,69,0,173,0,253,0,50,0,151,0,239,0,3,0,42,0,35,0,230,0,167,0,42,0,233,0,97,0,0,0,0,0,15,0,89,0,100,0,78,0,76,0,214,0,204,0,232,0,199,0,148,0,176,0,192,0,52,0,81,0,0,0,0,0,119,0,95,0,186,0,215,0,242,0,0,0,230,0,182,0,103,0,0,0,191,0,6,0,186,0,54,0,39,0,181,0,167,0,235,0,0,0,219,0,76,0,138,0,223,0,0,0,35,0,186,0,0,0,178,0,247,0,0,0,85,0,149,0,250,0,113,0,252,0,0,0,36,0,0,0,21,0,0,0,253,0,86,0,246,0,189,0,77,0,127,0,117,0,0,0,115,0,241,0,219,0,56,0,253,0,0,0,0,0,226,0,18,0,0,0,235,0,0,0,6,0,161,0,14,0,0,0,0,0,199,0,38,0,0,0,237,0,3,0,242,0,197,0,252,0,0,0,154,0,97,0,63,0,0,0,0,0);
signal scenario_full  : scenario_type := (138,31,96,31,96,30,138,31,138,30,207,31,192,31,221,31,194,31,94,31,115,31,86,31,197,31,150,31,150,30,96,31,220,31,42,31,42,30,184,31,15,31,236,31,177,31,102,31,102,30,135,31,69,31,26,31,26,30,26,29,210,31,147,31,251,31,95,31,165,31,17,31,53,31,179,31,122,31,83,31,14,31,14,30,18,31,180,31,158,31,101,31,57,31,197,31,197,30,33,31,125,31,40,31,255,31,255,30,3,31,82,31,82,30,67,31,240,31,218,31,219,31,248,31,3,31,3,30,3,29,254,31,222,31,215,31,196,31,196,30,196,29,196,28,196,27,232,31,56,31,5,31,92,31,32,31,65,31,140,31,157,31,133,31,153,31,176,31,137,31,60,31,60,30,60,29,32,31,209,31,76,31,121,31,121,30,191,31,145,31,132,31,206,31,57,31,31,31,7,31,238,31,238,30,108,31,59,31,159,31,60,31,129,31,117,31,178,31,32,31,222,31,179,31,221,31,178,31,178,30,185,31,95,31,1,31,170,31,127,31,90,31,25,31,91,31,136,31,140,31,79,31,81,31,81,30,47,31,226,31,191,31,191,30,239,31,160,31,248,31,248,30,107,31,224,31,85,31,248,31,248,30,132,31,132,30,132,29,137,31,160,31,107,31,223,31,223,30,243,31,243,30,46,31,46,30,172,31,171,31,206,31,198,31,198,30,127,31,173,31,9,31,73,31,16,31,16,30,92,31,7,31,11,31,11,30,38,31,56,31,218,31,67,31,94,31,34,31,34,30,184,31,29,31,148,31,127,31,70,31,26,31,229,31,184,31,173,31,113,31,158,31,212,31,130,31,89,31,44,31,179,31,179,30,197,31,197,30,197,29,169,31,128,31,128,30,188,31,188,30,246,31,246,30,127,31,138,31,138,30,211,31,111,31,29,31,48,31,166,31,216,31,16,31,16,30,218,31,40,31,40,30,13,31,196,31,114,31,114,30,99,31,115,31,20,31,93,31,170,31,170,30,101,31,154,31,34,31,34,30,34,29,34,28,34,27,202,31,230,31,230,30,230,29,59,31,59,30,25,31,246,31,162,31,89,31,108,31,101,31,3,31,3,30,22,31,28,31,183,31,199,31,135,31,133,31,77,31,159,31,88,31,219,31,165,31,131,31,27,31,168,31,168,30,235,31,204,31,204,30,179,31,168,31,64,31,150,31,150,30,150,29,102,31,23,31,169,31,15,31,15,30,175,31,242,31,28,31,180,31,115,31,83,31,83,30,160,31,62,31,4,31,200,31,149,31,6,31,202,31,128,31,182,31,104,31,118,31,20,31,254,31,15,31,54,31,73,31,1,31,1,30,156,31,230,31,67,31,114,31,145,31,39,31,251,31,251,30,149,31,149,30,149,29,149,28,89,31,248,31,248,30,173,31,162,31,186,31,253,31,142,31,194,31,235,31,3,31,236,31,178,31,191,31,29,31,117,31,151,31,233,31,185,31,185,30,70,31,129,31,157,31,247,31,60,31,73,31,196,31,187,31,187,30,235,31,235,30,46,31,72,31,42,31,226,31,63,31,63,30,71,31,198,31,8,31,167,31,49,31,150,31,202,31,129,31,129,30,248,31,109,31,255,31,201,31,201,30,251,31,126,31,142,31,66,31,222,31,122,31,176,31,185,31,252,31,208,31,122,31,122,30,16,31,84,31,19,31,19,30,102,31,170,31,168,31,29,31,29,30,29,29,13,31,19,31,246,31,154,31,163,31,163,30,57,31,14,31,121,31,121,30,183,31,147,31,147,30,211,31,128,31,247,31,69,31,117,31,138,31,115,31,115,30,90,31,173,31,229,31,45,31,139,31,139,30,102,31,102,30,96,31,12,31,73,31,101,31,191,31,15,31,107,31,204,31,181,31,138,31,83,31,48,31,48,30,233,31,25,31,244,31,29,31,34,31,34,30,191,31,191,30,246,31,208,31,129,31,129,30,169,31,182,31,195,31,174,31,127,31,103,31,115,31,176,31,35,31,239,31,30,31,101,31,114,31,114,30,104,31,104,30,104,29,144,31,248,31,171,31,171,30,249,31,88,31,40,31,170,31,194,31,102,31,102,30,97,31,44,31,175,31,171,31,183,31,188,31,188,30,226,31,52,31,209,31,188,31,123,31,123,30,123,29,123,28,123,27,123,26,17,31,18,31,250,31,125,31,158,31,152,31,152,30,145,31,206,31,115,31,205,31,205,30,6,31,239,31,78,31,176,31,212,31,212,30,65,31,53,31,43,31,43,30,189,31,189,30,130,31,193,31,193,30,193,29,148,31,54,31,85,31,85,30,198,31,167,31,167,30,98,31,20,31,239,31,91,31,121,31,130,31,228,31,213,31,214,31,214,30,38,31,84,31,84,30,122,31,2,31,79,31,127,31,122,31,26,31,26,30,26,29,226,31,99,31,80,31,165,31,165,30,165,29,165,28,38,31,124,31,212,31,161,31,163,31,3,31,163,31,103,31,142,31,170,31,250,31,245,31,142,31,226,31,172,31,204,31,124,31,117,31,91,31,82,31,252,31,216,31,251,31,241,31,200,31,253,31,84,31,84,30,56,31,249,31,249,30,28,31,244,31,105,31,186,31,166,31,151,31,106,31,157,31,157,30,230,31,127,31,235,31,52,31,138,31,46,31,71,31,227,31,180,31,109,31,147,31,33,31,218,31,218,30,165,31,128,31,128,30,67,31,61,31,61,30,116,31,67,31,66,31,49,31,49,30,49,29,214,31,214,30,214,29,5,31,78,31,80,31,192,31,69,31,173,31,253,31,50,31,151,31,239,31,3,31,42,31,35,31,230,31,167,31,42,31,233,31,97,31,97,30,97,29,15,31,89,31,100,31,78,31,76,31,214,31,204,31,232,31,199,31,148,31,176,31,192,31,52,31,81,31,81,30,81,29,119,31,95,31,186,31,215,31,242,31,242,30,230,31,182,31,103,31,103,30,191,31,6,31,186,31,54,31,39,31,181,31,167,31,235,31,235,30,219,31,76,31,138,31,223,31,223,30,35,31,186,31,186,30,178,31,247,31,247,30,85,31,149,31,250,31,113,31,252,31,252,30,36,31,36,30,21,31,21,30,253,31,86,31,246,31,189,31,77,31,127,31,117,31,117,30,115,31,241,31,219,31,56,31,253,31,253,30,253,29,226,31,18,31,18,30,235,31,235,30,6,31,161,31,14,31,14,30,14,29,199,31,38,31,38,30,237,31,3,31,242,31,197,31,252,31,252,30,154,31,97,31,63,31,63,30,63,29);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
