-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 204;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (138,0,36,0,141,0,45,0,60,0,205,0,70,0,0,0,113,0,0,0,156,0,128,0,199,0,105,0,6,0,148,0,60,0,152,0,0,0,211,0,176,0,85,0,1,0,85,0,79,0,79,0,131,0,0,0,62,0,230,0,30,0,154,0,251,0,120,0,55,0,41,0,62,0,0,0,88,0,157,0,0,0,121,0,182,0,140,0,215,0,0,0,3,0,0,0,188,0,166,0,62,0,198,0,64,0,228,0,206,0,35,0,83,0,124,0,49,0,60,0,131,0,192,0,0,0,188,0,73,0,218,0,0,0,222,0,214,0,92,0,94,0,178,0,215,0,0,0,14,0,202,0,61,0,0,0,97,0,138,0,42,0,251,0,52,0,31,0,244,0,158,0,186,0,0,0,181,0,199,0,232,0,243,0,196,0,134,0,245,0,0,0,70,0,227,0,185,0,0,0,140,0,167,0,45,0,250,0,0,0,72,0,232,0,0,0,26,0,15,0,0,0,17,0,229,0,0,0,243,0,31,0,67,0,0,0,56,0,118,0,169,0,30,0,25,0,74,0,209,0,0,0,83,0,0,0,254,0,212,0,0,0,0,0,153,0,20,0,160,0,158,0,204,0,188,0,162,0,0,0,202,0,85,0,83,0,158,0,0,0,195,0,0,0,163,0,212,0,106,0,130,0,128,0,238,0,136,0,5,0,129,0,71,0,221,0,136,0,16,0,0,0,0,0,153,0,52,0,202,0,208,0,76,0,90,0,52,0,108,0,216,0,5,0,200,0,15,0,159,0,237,0,0,0,40,0,209,0,212,0,227,0,175,0,117,0,5,0,0,0,171,0,233,0,94,0,16,0,5,0,201,0,216,0,127,0,150,0,94,0,160,0,117,0,195,0,167,0,68,0,111,0,215,0,127,0,243,0);
signal scenario_full  : scenario_type := (138,31,36,31,141,31,45,31,60,31,205,31,70,31,70,30,113,31,113,30,156,31,128,31,199,31,105,31,6,31,148,31,60,31,152,31,152,30,211,31,176,31,85,31,1,31,85,31,79,31,79,31,131,31,131,30,62,31,230,31,30,31,154,31,251,31,120,31,55,31,41,31,62,31,62,30,88,31,157,31,157,30,121,31,182,31,140,31,215,31,215,30,3,31,3,30,188,31,166,31,62,31,198,31,64,31,228,31,206,31,35,31,83,31,124,31,49,31,60,31,131,31,192,31,192,30,188,31,73,31,218,31,218,30,222,31,214,31,92,31,94,31,178,31,215,31,215,30,14,31,202,31,61,31,61,30,97,31,138,31,42,31,251,31,52,31,31,31,244,31,158,31,186,31,186,30,181,31,199,31,232,31,243,31,196,31,134,31,245,31,245,30,70,31,227,31,185,31,185,30,140,31,167,31,45,31,250,31,250,30,72,31,232,31,232,30,26,31,15,31,15,30,17,31,229,31,229,30,243,31,31,31,67,31,67,30,56,31,118,31,169,31,30,31,25,31,74,31,209,31,209,30,83,31,83,30,254,31,212,31,212,30,212,29,153,31,20,31,160,31,158,31,204,31,188,31,162,31,162,30,202,31,85,31,83,31,158,31,158,30,195,31,195,30,163,31,212,31,106,31,130,31,128,31,238,31,136,31,5,31,129,31,71,31,221,31,136,31,16,31,16,30,16,29,153,31,52,31,202,31,208,31,76,31,90,31,52,31,108,31,216,31,5,31,200,31,15,31,159,31,237,31,237,30,40,31,209,31,212,31,227,31,175,31,117,31,5,31,5,30,171,31,233,31,94,31,16,31,5,31,201,31,216,31,127,31,150,31,94,31,160,31,117,31,195,31,167,31,68,31,111,31,215,31,127,31,243,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
