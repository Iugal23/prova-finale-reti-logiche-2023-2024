-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_998 is
end project_tb_998;

architecture project_tb_arch_998 of project_tb_998 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 820;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (214,0,88,0,132,0,135,0,222,0,128,0,117,0,0,0,11,0,111,0,91,0,214,0,0,0,252,0,0,0,231,0,0,0,178,0,208,0,146,0,87,0,209,0,9,0,0,0,121,0,0,0,169,0,9,0,17,0,0,0,17,0,19,0,221,0,0,0,85,0,0,0,108,0,183,0,215,0,0,0,235,0,147,0,197,0,0,0,0,0,41,0,166,0,159,0,223,0,244,0,124,0,158,0,73,0,0,0,73,0,235,0,58,0,81,0,125,0,217,0,111,0,105,0,0,0,149,0,186,0,0,0,181,0,0,0,2,0,0,0,203,0,9,0,103,0,76,0,44,0,193,0,34,0,187,0,21,0,240,0,0,0,0,0,0,0,158,0,44,0,234,0,176,0,92,0,104,0,0,0,0,0,78,0,17,0,0,0,245,0,42,0,116,0,193,0,0,0,149,0,119,0,210,0,223,0,0,0,140,0,30,0,225,0,249,0,144,0,245,0,155,0,0,0,98,0,220,0,17,0,0,0,107,0,0,0,142,0,2,0,36,0,0,0,0,0,99,0,0,0,9,0,155,0,204,0,209,0,129,0,33,0,152,0,150,0,184,0,77,0,169,0,20,0,204,0,233,0,3,0,102,0,169,0,62,0,83,0,171,0,172,0,246,0,218,0,164,0,55,0,65,0,0,0,0,0,112,0,165,0,140,0,171,0,32,0,197,0,189,0,198,0,222,0,131,0,93,0,0,0,0,0,129,0,175,0,66,0,0,0,139,0,255,0,97,0,98,0,59,0,159,0,90,0,158,0,85,0,148,0,13,0,135,0,0,0,75,0,36,0,174,0,235,0,0,0,129,0,39,0,0,0,0,0,0,0,185,0,188,0,99,0,118,0,159,0,88,0,244,0,225,0,200,0,2,0,0,0,122,0,227,0,66,0,0,0,238,0,83,0,0,0,180,0,122,0,0,0,0,0,48,0,192,0,179,0,191,0,0,0,157,0,185,0,192,0,139,0,0,0,85,0,0,0,222,0,155,0,93,0,0,0,237,0,79,0,243,0,247,0,33,0,0,0,136,0,95,0,80,0,79,0,108,0,247,0,213,0,77,0,184,0,0,0,43,0,57,0,157,0,35,0,220,0,194,0,59,0,0,0,0,0,101,0,169,0,0,0,37,0,201,0,0,0,13,0,129,0,120,0,47,0,0,0,209,0,0,0,0,0,72,0,65,0,84,0,0,0,0,0,214,0,0,0,224,0,0,0,246,0,33,0,137,0,84,0,0,0,217,0,220,0,222,0,254,0,1,0,199,0,138,0,143,0,39,0,104,0,0,0,0,0,16,0,126,0,44,0,0,0,242,0,151,0,41,0,244,0,38,0,0,0,58,0,112,0,82,0,77,0,12,0,240,0,86,0,0,0,51,0,0,0,0,0,254,0,129,0,209,0,129,0,250,0,0,0,0,0,117,0,15,0,188,0,236,0,0,0,45,0,103,0,0,0,0,0,121,0,219,0,209,0,188,0,37,0,13,0,241,0,0,0,154,0,151,0,241,0,83,0,220,0,251,0,142,0,213,0,38,0,0,0,238,0,20,0,36,0,55,0,0,0,250,0,0,0,106,0,0,0,234,0,0,0,0,0,64,0,0,0,133,0,78,0,125,0,174,0,0,0,6,0,14,0,83,0,187,0,75,0,200,0,139,0,0,0,185,0,173,0,155,0,196,0,89,0,223,0,122,0,20,0,0,0,167,0,166,0,87,0,113,0,212,0,137,0,65,0,252,0,182,0,101,0,127,0,201,0,22,0,67,0,0,0,0,0,44,0,77,0,198,0,210,0,92,0,0,0,77,0,15,0,71,0,223,0,40,0,0,0,0,0,12,0,248,0,0,0,143,0,0,0,48,0,184,0,163,0,0,0,195,0,225,0,220,0,188,0,136,0,0,0,190,0,67,0,177,0,4,0,197,0,212,0,4,0,161,0,55,0,0,0,245,0,144,0,24,0,117,0,87,0,182,0,0,0,180,0,68,0,0,0,12,0,213,0,0,0,160,0,228,0,86,0,89,0,15,0,0,0,34,0,152,0,225,0,164,0,55,0,115,0,136,0,190,0,96,0,58,0,81,0,26,0,114,0,213,0,37,0,191,0,161,0,9,0,0,0,177,0,103,0,59,0,0,0,46,0,17,0,246,0,0,0,85,0,159,0,152,0,88,0,56,0,0,0,56,0,81,0,199,0,210,0,209,0,3,0,125,0,177,0,54,0,128,0,0,0,200,0,84,0,52,0,193,0,106,0,130,0,72,0,82,0,132,0,202,0,0,0,156,0,244,0,241,0,17,0,6,0,213,0,36,0,180,0,142,0,0,0,186,0,200,0,126,0,0,0,0,0,81,0,7,0,220,0,8,0,210,0,196,0,198,0,55,0,242,0,58,0,0,0,118,0,109,0,218,0,152,0,159,0,253,0,194,0,238,0,112,0,83,0,182,0,0,0,248,0,118,0,109,0,0,0,0,0,120,0,217,0,27,0,54,0,103,0,0,0,162,0,0,0,246,0,245,0,222,0,223,0,187,0,106,0,56,0,155,0,106,0,0,0,0,0,126,0,0,0,30,0,224,0,0,0,0,0,149,0,67,0,0,0,0,0,248,0,8,0,51,0,0,0,221,0,0,0,0,0,5,0,116,0,52,0,228,0,15,0,40,0,0,0,50,0,0,0,0,0,187,0,0,0,212,0,238,0,251,0,175,0,170,0,144,0,56,0,8,0,181,0,134,0,0,0,0,0,0,0,244,0,31,0,248,0,240,0,111,0,103,0,0,0,92,0,87,0,224,0,173,0,161,0,0,0,53,0,0,0,77,0,101,0,171,0,208,0,186,0,31,0,0,0,0,0,224,0,44,0,255,0,127,0,147,0,136,0,95,0,165,0,0,0,114,0,87,0,236,0,246,0,19,0,58,0,11,0,128,0,219,0,0,0,0,0,0,0,105,0,0,0,82,0,253,0,153,0,187,0,194,0,156,0,206,0,67,0,184,0,22,0,229,0,221,0,28,0,167,0,241,0,230,0,107,0,56,0,0,0,167,0,176,0,161,0,0,0,148,0,39,0,201,0,0,0,97,0,31,0,0,0,156,0,205,0,0,0,0,0,60,0,181,0,0,0,235,0,15,0,214,0,129,0,51,0,12,0,0,0,0,0,18,0,177,0,94,0,27,0,99,0,89,0,51,0,0,0,205,0,242,0,38,0,113,0,239,0,123,0,219,0,142,0,3,0,0,0,0,0,113,0,0,0,0,0,87,0,52,0,100,0,180,0,242,0,93,0,0,0,122,0,159,0,138,0,253,0,225,0,209,0,184,0,142,0,218,0,168,0,0,0,51,0,17,0,219,0,29,0,60,0,151,0,0,0,0,0,0,0,168,0,62,0,150,0,63,0,75,0,53,0,52,0,47,0,59,0,255,0,0,0,181,0,0,0,56,0,96,0,70,0,19,0,0,0,52,0,113,0,31,0,68,0,0,0,20,0,234,0,88,0,69,0,0,0,90,0,34,0,157,0,176,0,115,0,240,0,129,0,99,0,128,0,175,0,0,0,238,0,0,0,212,0,0,0,105,0,22,0,169,0,190,0,31,0,173,0,222,0,107,0,229,0,3,0,52,0,234,0,239,0,179,0,141,0,0,0,100,0,14,0);
signal scenario_full  : scenario_type := (214,31,88,31,132,31,135,31,222,31,128,31,117,31,117,30,11,31,111,31,91,31,214,31,214,30,252,31,252,30,231,31,231,30,178,31,208,31,146,31,87,31,209,31,9,31,9,30,121,31,121,30,169,31,9,31,17,31,17,30,17,31,19,31,221,31,221,30,85,31,85,30,108,31,183,31,215,31,215,30,235,31,147,31,197,31,197,30,197,29,41,31,166,31,159,31,223,31,244,31,124,31,158,31,73,31,73,30,73,31,235,31,58,31,81,31,125,31,217,31,111,31,105,31,105,30,149,31,186,31,186,30,181,31,181,30,2,31,2,30,203,31,9,31,103,31,76,31,44,31,193,31,34,31,187,31,21,31,240,31,240,30,240,29,240,28,158,31,44,31,234,31,176,31,92,31,104,31,104,30,104,29,78,31,17,31,17,30,245,31,42,31,116,31,193,31,193,30,149,31,119,31,210,31,223,31,223,30,140,31,30,31,225,31,249,31,144,31,245,31,155,31,155,30,98,31,220,31,17,31,17,30,107,31,107,30,142,31,2,31,36,31,36,30,36,29,99,31,99,30,9,31,155,31,204,31,209,31,129,31,33,31,152,31,150,31,184,31,77,31,169,31,20,31,204,31,233,31,3,31,102,31,169,31,62,31,83,31,171,31,172,31,246,31,218,31,164,31,55,31,65,31,65,30,65,29,112,31,165,31,140,31,171,31,32,31,197,31,189,31,198,31,222,31,131,31,93,31,93,30,93,29,129,31,175,31,66,31,66,30,139,31,255,31,97,31,98,31,59,31,159,31,90,31,158,31,85,31,148,31,13,31,135,31,135,30,75,31,36,31,174,31,235,31,235,30,129,31,39,31,39,30,39,29,39,28,185,31,188,31,99,31,118,31,159,31,88,31,244,31,225,31,200,31,2,31,2,30,122,31,227,31,66,31,66,30,238,31,83,31,83,30,180,31,122,31,122,30,122,29,48,31,192,31,179,31,191,31,191,30,157,31,185,31,192,31,139,31,139,30,85,31,85,30,222,31,155,31,93,31,93,30,237,31,79,31,243,31,247,31,33,31,33,30,136,31,95,31,80,31,79,31,108,31,247,31,213,31,77,31,184,31,184,30,43,31,57,31,157,31,35,31,220,31,194,31,59,31,59,30,59,29,101,31,169,31,169,30,37,31,201,31,201,30,13,31,129,31,120,31,47,31,47,30,209,31,209,30,209,29,72,31,65,31,84,31,84,30,84,29,214,31,214,30,224,31,224,30,246,31,33,31,137,31,84,31,84,30,217,31,220,31,222,31,254,31,1,31,199,31,138,31,143,31,39,31,104,31,104,30,104,29,16,31,126,31,44,31,44,30,242,31,151,31,41,31,244,31,38,31,38,30,58,31,112,31,82,31,77,31,12,31,240,31,86,31,86,30,51,31,51,30,51,29,254,31,129,31,209,31,129,31,250,31,250,30,250,29,117,31,15,31,188,31,236,31,236,30,45,31,103,31,103,30,103,29,121,31,219,31,209,31,188,31,37,31,13,31,241,31,241,30,154,31,151,31,241,31,83,31,220,31,251,31,142,31,213,31,38,31,38,30,238,31,20,31,36,31,55,31,55,30,250,31,250,30,106,31,106,30,234,31,234,30,234,29,64,31,64,30,133,31,78,31,125,31,174,31,174,30,6,31,14,31,83,31,187,31,75,31,200,31,139,31,139,30,185,31,173,31,155,31,196,31,89,31,223,31,122,31,20,31,20,30,167,31,166,31,87,31,113,31,212,31,137,31,65,31,252,31,182,31,101,31,127,31,201,31,22,31,67,31,67,30,67,29,44,31,77,31,198,31,210,31,92,31,92,30,77,31,15,31,71,31,223,31,40,31,40,30,40,29,12,31,248,31,248,30,143,31,143,30,48,31,184,31,163,31,163,30,195,31,225,31,220,31,188,31,136,31,136,30,190,31,67,31,177,31,4,31,197,31,212,31,4,31,161,31,55,31,55,30,245,31,144,31,24,31,117,31,87,31,182,31,182,30,180,31,68,31,68,30,12,31,213,31,213,30,160,31,228,31,86,31,89,31,15,31,15,30,34,31,152,31,225,31,164,31,55,31,115,31,136,31,190,31,96,31,58,31,81,31,26,31,114,31,213,31,37,31,191,31,161,31,9,31,9,30,177,31,103,31,59,31,59,30,46,31,17,31,246,31,246,30,85,31,159,31,152,31,88,31,56,31,56,30,56,31,81,31,199,31,210,31,209,31,3,31,125,31,177,31,54,31,128,31,128,30,200,31,84,31,52,31,193,31,106,31,130,31,72,31,82,31,132,31,202,31,202,30,156,31,244,31,241,31,17,31,6,31,213,31,36,31,180,31,142,31,142,30,186,31,200,31,126,31,126,30,126,29,81,31,7,31,220,31,8,31,210,31,196,31,198,31,55,31,242,31,58,31,58,30,118,31,109,31,218,31,152,31,159,31,253,31,194,31,238,31,112,31,83,31,182,31,182,30,248,31,118,31,109,31,109,30,109,29,120,31,217,31,27,31,54,31,103,31,103,30,162,31,162,30,246,31,245,31,222,31,223,31,187,31,106,31,56,31,155,31,106,31,106,30,106,29,126,31,126,30,30,31,224,31,224,30,224,29,149,31,67,31,67,30,67,29,248,31,8,31,51,31,51,30,221,31,221,30,221,29,5,31,116,31,52,31,228,31,15,31,40,31,40,30,50,31,50,30,50,29,187,31,187,30,212,31,238,31,251,31,175,31,170,31,144,31,56,31,8,31,181,31,134,31,134,30,134,29,134,28,244,31,31,31,248,31,240,31,111,31,103,31,103,30,92,31,87,31,224,31,173,31,161,31,161,30,53,31,53,30,77,31,101,31,171,31,208,31,186,31,31,31,31,30,31,29,224,31,44,31,255,31,127,31,147,31,136,31,95,31,165,31,165,30,114,31,87,31,236,31,246,31,19,31,58,31,11,31,128,31,219,31,219,30,219,29,219,28,105,31,105,30,82,31,253,31,153,31,187,31,194,31,156,31,206,31,67,31,184,31,22,31,229,31,221,31,28,31,167,31,241,31,230,31,107,31,56,31,56,30,167,31,176,31,161,31,161,30,148,31,39,31,201,31,201,30,97,31,31,31,31,30,156,31,205,31,205,30,205,29,60,31,181,31,181,30,235,31,15,31,214,31,129,31,51,31,12,31,12,30,12,29,18,31,177,31,94,31,27,31,99,31,89,31,51,31,51,30,205,31,242,31,38,31,113,31,239,31,123,31,219,31,142,31,3,31,3,30,3,29,113,31,113,30,113,29,87,31,52,31,100,31,180,31,242,31,93,31,93,30,122,31,159,31,138,31,253,31,225,31,209,31,184,31,142,31,218,31,168,31,168,30,51,31,17,31,219,31,29,31,60,31,151,31,151,30,151,29,151,28,168,31,62,31,150,31,63,31,75,31,53,31,52,31,47,31,59,31,255,31,255,30,181,31,181,30,56,31,96,31,70,31,19,31,19,30,52,31,113,31,31,31,68,31,68,30,20,31,234,31,88,31,69,31,69,30,90,31,34,31,157,31,176,31,115,31,240,31,129,31,99,31,128,31,175,31,175,30,238,31,238,30,212,31,212,30,105,31,22,31,169,31,190,31,31,31,173,31,222,31,107,31,229,31,3,31,52,31,234,31,239,31,179,31,141,31,141,30,100,31,14,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
