-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 251;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (187,0,216,0,41,0,191,0,0,0,62,0,244,0,111,0,26,0,164,0,40,0,19,0,60,0,136,0,0,0,0,0,112,0,25,0,0,0,195,0,235,0,59,0,231,0,129,0,94,0,246,0,47,0,176,0,13,0,123,0,46,0,75,0,172,0,119,0,0,0,15,0,190,0,132,0,0,0,0,0,142,0,7,0,0,0,0,0,102,0,253,0,224,0,74,0,127,0,168,0,115,0,88,0,154,0,167,0,223,0,241,0,244,0,253,0,147,0,104,0,0,0,25,0,184,0,92,0,247,0,0,0,165,0,0,0,0,0,38,0,86,0,0,0,183,0,150,0,69,0,221,0,243,0,92,0,29,0,196,0,152,0,88,0,124,0,147,0,228,0,91,0,113,0,233,0,62,0,250,0,102,0,83,0,51,0,37,0,176,0,236,0,204,0,0,0,161,0,0,0,0,0,0,0,129,0,202,0,77,0,182,0,197,0,202,0,0,0,25,0,0,0,0,0,0,0,65,0,0,0,243,0,0,0,0,0,168,0,0,0,100,0,4,0,44,0,107,0,247,0,130,0,148,0,7,0,160,0,60,0,107,0,255,0,68,0,94,0,169,0,150,0,137,0,160,0,0,0,0,0,101,0,168,0,238,0,49,0,65,0,46,0,199,0,121,0,11,0,95,0,63,0,0,0,0,0,0,0,0,0,134,0,214,0,124,0,113,0,98,0,226,0,42,0,8,0,0,0,0,0,141,0,125,0,150,0,19,0,186,0,191,0,160,0,77,0,235,0,29,0,0,0,0,0,167,0,57,0,120,0,148,0,166,0,134,0,101,0,98,0,232,0,141,0,139,0,251,0,247,0,42,0,155,0,100,0,74,0,0,0,165,0,0,0,161,0,10,0,143,0,212,0,177,0,216,0,1,0,2,0,154,0,188,0,178,0,61,0,0,0,144,0,250,0,229,0,128,0,104,0,0,0,63,0,222,0,173,0,250,0,176,0,230,0,0,0,205,0,1,0,46,0,254,0,91,0,157,0,133,0,0,0,0,0,0,0,0,0,162,0,237,0,26,0,0,0,192,0,251,0,61,0,132,0,117,0,23,0,94,0,0,0,0,0,253,0,185,0,192,0,235,0);
signal scenario_full  : scenario_type := (187,31,216,31,41,31,191,31,191,30,62,31,244,31,111,31,26,31,164,31,40,31,19,31,60,31,136,31,136,30,136,29,112,31,25,31,25,30,195,31,235,31,59,31,231,31,129,31,94,31,246,31,47,31,176,31,13,31,123,31,46,31,75,31,172,31,119,31,119,30,15,31,190,31,132,31,132,30,132,29,142,31,7,31,7,30,7,29,102,31,253,31,224,31,74,31,127,31,168,31,115,31,88,31,154,31,167,31,223,31,241,31,244,31,253,31,147,31,104,31,104,30,25,31,184,31,92,31,247,31,247,30,165,31,165,30,165,29,38,31,86,31,86,30,183,31,150,31,69,31,221,31,243,31,92,31,29,31,196,31,152,31,88,31,124,31,147,31,228,31,91,31,113,31,233,31,62,31,250,31,102,31,83,31,51,31,37,31,176,31,236,31,204,31,204,30,161,31,161,30,161,29,161,28,129,31,202,31,77,31,182,31,197,31,202,31,202,30,25,31,25,30,25,29,25,28,65,31,65,30,243,31,243,30,243,29,168,31,168,30,100,31,4,31,44,31,107,31,247,31,130,31,148,31,7,31,160,31,60,31,107,31,255,31,68,31,94,31,169,31,150,31,137,31,160,31,160,30,160,29,101,31,168,31,238,31,49,31,65,31,46,31,199,31,121,31,11,31,95,31,63,31,63,30,63,29,63,28,63,27,134,31,214,31,124,31,113,31,98,31,226,31,42,31,8,31,8,30,8,29,141,31,125,31,150,31,19,31,186,31,191,31,160,31,77,31,235,31,29,31,29,30,29,29,167,31,57,31,120,31,148,31,166,31,134,31,101,31,98,31,232,31,141,31,139,31,251,31,247,31,42,31,155,31,100,31,74,31,74,30,165,31,165,30,161,31,10,31,143,31,212,31,177,31,216,31,1,31,2,31,154,31,188,31,178,31,61,31,61,30,144,31,250,31,229,31,128,31,104,31,104,30,63,31,222,31,173,31,250,31,176,31,230,31,230,30,205,31,1,31,46,31,254,31,91,31,157,31,133,31,133,30,133,29,133,28,133,27,162,31,237,31,26,31,26,30,192,31,251,31,61,31,132,31,117,31,23,31,94,31,94,30,94,29,253,31,185,31,192,31,235,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
