-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 448;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,71,0,194,0,101,0,0,0,161,0,164,0,47,0,116,0,20,0,36,0,61,0,47,0,243,0,190,0,110,0,0,0,0,0,7,0,0,0,8,0,27,0,170,0,0,0,232,0,238,0,39,0,32,0,86,0,0,0,222,0,23,0,154,0,0,0,0,0,44,0,54,0,140,0,0,0,214,0,25,0,224,0,139,0,0,0,0,0,95,0,0,0,201,0,0,0,96,0,0,0,58,0,96,0,134,0,37,0,198,0,181,0,235,0,135,0,237,0,39,0,40,0,176,0,81,0,139,0,115,0,167,0,77,0,130,0,202,0,40,0,106,0,0,0,253,0,68,0,0,0,0,0,50,0,213,0,160,0,147,0,0,0,141,0,85,0,0,0,173,0,148,0,0,0,159,0,0,0,204,0,0,0,133,0,122,0,165,0,170,0,147,0,11,0,138,0,181,0,0,0,173,0,0,0,138,0,54,0,7,0,170,0,156,0,0,0,118,0,239,0,152,0,104,0,97,0,126,0,150,0,243,0,230,0,0,0,0,0,67,0,0,0,59,0,0,0,83,0,84,0,253,0,108,0,0,0,27,0,45,0,0,0,177,0,192,0,0,0,9,0,0,0,83,0,135,0,176,0,39,0,162,0,0,0,175,0,45,0,0,0,199,0,238,0,186,0,171,0,214,0,63,0,165,0,0,0,0,0,77,0,200,0,110,0,0,0,149,0,184,0,248,0,202,0,73,0,0,0,99,0,72,0,186,0,229,0,167,0,87,0,93,0,28,0,193,0,198,0,95,0,0,0,0,0,120,0,183,0,116,0,0,0,0,0,0,0,145,0,29,0,0,0,80,0,125,0,177,0,193,0,0,0,138,0,0,0,219,0,144,0,19,0,0,0,84,0,253,0,43,0,65,0,52,0,73,0,107,0,179,0,78,0,232,0,38,0,206,0,228,0,103,0,81,0,255,0,169,0,0,0,177,0,184,0,146,0,64,0,204,0,37,0,99,0,88,0,83,0,218,0,163,0,73,0,77,0,110,0,0,0,50,0,165,0,115,0,218,0,205,0,52,0,56,0,166,0,0,0,0,0,173,0,82,0,98,0,33,0,179,0,26,0,214,0,113,0,16,0,0,0,133,0,0,0,0,0,226,0,249,0,0,0,230,0,161,0,241,0,52,0,1,0,137,0,180,0,193,0,0,0,179,0,202,0,237,0,207,0,78,0,93,0,195,0,129,0,60,0,60,0,178,0,194,0,115,0,37,0,95,0,121,0,66,0,0,0,148,0,136,0,146,0,48,0,0,0,239,0,183,0,0,0,157,0,84,0,118,0,19,0,10,0,208,0,0,0,201,0,216,0,80,0,252,0,0,0,59,0,70,0,2,0,40,0,215,0,117,0,173,0,0,0,0,0,214,0,60,0,36,0,252,0,0,0,0,0,242,0,80,0,133,0,114,0,112,0,33,0,147,0,57,0,125,0,5,0,0,0,187,0,240,0,212,0,111,0,122,0,245,0,2,0,165,0,37,0,229,0,19,0,0,0,245,0,173,0,69,0,207,0,63,0,232,0,217,0,200,0,228,0,0,0,214,0,109,0,0,0,16,0,209,0,244,0,18,0,95,0,232,0,162,0,0,0,127,0,89,0,0,0,79,0,158,0,0,0,0,0,47,0,9,0,213,0,0,0,64,0,0,0,203,0,214,0,129,0,0,0,0,0,111,0,89,0,0,0,87,0,179,0,184,0,0,0,224,0,119,0,14,0,252,0,171,0,178,0,184,0,134,0,182,0,53,0,0,0,41,0,23,0,215,0,156,0,196,0,146,0,204,0,0,0,109,0,26,0,0,0,0,0,181,0,45,0,34,0,0,0,143,0,86,0,0,0,185,0,166,0,74,0,0,0,21,0,107,0,209,0,43,0,0,0,0,0,46,0,151,0,72,0,126,0,38,0,133,0,229,0,218,0,0,0,203,0,76,0,0,0,115,0,0,0,138,0,0,0,212,0,159,0,69,0,13,0);
signal scenario_full  : scenario_type := (0,0,71,31,194,31,101,31,101,30,161,31,164,31,47,31,116,31,20,31,36,31,61,31,47,31,243,31,190,31,110,31,110,30,110,29,7,31,7,30,8,31,27,31,170,31,170,30,232,31,238,31,39,31,32,31,86,31,86,30,222,31,23,31,154,31,154,30,154,29,44,31,54,31,140,31,140,30,214,31,25,31,224,31,139,31,139,30,139,29,95,31,95,30,201,31,201,30,96,31,96,30,58,31,96,31,134,31,37,31,198,31,181,31,235,31,135,31,237,31,39,31,40,31,176,31,81,31,139,31,115,31,167,31,77,31,130,31,202,31,40,31,106,31,106,30,253,31,68,31,68,30,68,29,50,31,213,31,160,31,147,31,147,30,141,31,85,31,85,30,173,31,148,31,148,30,159,31,159,30,204,31,204,30,133,31,122,31,165,31,170,31,147,31,11,31,138,31,181,31,181,30,173,31,173,30,138,31,54,31,7,31,170,31,156,31,156,30,118,31,239,31,152,31,104,31,97,31,126,31,150,31,243,31,230,31,230,30,230,29,67,31,67,30,59,31,59,30,83,31,84,31,253,31,108,31,108,30,27,31,45,31,45,30,177,31,192,31,192,30,9,31,9,30,83,31,135,31,176,31,39,31,162,31,162,30,175,31,45,31,45,30,199,31,238,31,186,31,171,31,214,31,63,31,165,31,165,30,165,29,77,31,200,31,110,31,110,30,149,31,184,31,248,31,202,31,73,31,73,30,99,31,72,31,186,31,229,31,167,31,87,31,93,31,28,31,193,31,198,31,95,31,95,30,95,29,120,31,183,31,116,31,116,30,116,29,116,28,145,31,29,31,29,30,80,31,125,31,177,31,193,31,193,30,138,31,138,30,219,31,144,31,19,31,19,30,84,31,253,31,43,31,65,31,52,31,73,31,107,31,179,31,78,31,232,31,38,31,206,31,228,31,103,31,81,31,255,31,169,31,169,30,177,31,184,31,146,31,64,31,204,31,37,31,99,31,88,31,83,31,218,31,163,31,73,31,77,31,110,31,110,30,50,31,165,31,115,31,218,31,205,31,52,31,56,31,166,31,166,30,166,29,173,31,82,31,98,31,33,31,179,31,26,31,214,31,113,31,16,31,16,30,133,31,133,30,133,29,226,31,249,31,249,30,230,31,161,31,241,31,52,31,1,31,137,31,180,31,193,31,193,30,179,31,202,31,237,31,207,31,78,31,93,31,195,31,129,31,60,31,60,31,178,31,194,31,115,31,37,31,95,31,121,31,66,31,66,30,148,31,136,31,146,31,48,31,48,30,239,31,183,31,183,30,157,31,84,31,118,31,19,31,10,31,208,31,208,30,201,31,216,31,80,31,252,31,252,30,59,31,70,31,2,31,40,31,215,31,117,31,173,31,173,30,173,29,214,31,60,31,36,31,252,31,252,30,252,29,242,31,80,31,133,31,114,31,112,31,33,31,147,31,57,31,125,31,5,31,5,30,187,31,240,31,212,31,111,31,122,31,245,31,2,31,165,31,37,31,229,31,19,31,19,30,245,31,173,31,69,31,207,31,63,31,232,31,217,31,200,31,228,31,228,30,214,31,109,31,109,30,16,31,209,31,244,31,18,31,95,31,232,31,162,31,162,30,127,31,89,31,89,30,79,31,158,31,158,30,158,29,47,31,9,31,213,31,213,30,64,31,64,30,203,31,214,31,129,31,129,30,129,29,111,31,89,31,89,30,87,31,179,31,184,31,184,30,224,31,119,31,14,31,252,31,171,31,178,31,184,31,134,31,182,31,53,31,53,30,41,31,23,31,215,31,156,31,196,31,146,31,204,31,204,30,109,31,26,31,26,30,26,29,181,31,45,31,34,31,34,30,143,31,86,31,86,30,185,31,166,31,74,31,74,30,21,31,107,31,209,31,43,31,43,30,43,29,46,31,151,31,72,31,126,31,38,31,133,31,229,31,218,31,218,30,203,31,76,31,76,30,115,31,115,30,138,31,138,30,212,31,159,31,69,31,13,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
