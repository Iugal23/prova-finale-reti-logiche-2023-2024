-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_218 is
end project_tb_218;

architecture project_tb_arch_218 of project_tb_218 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 658;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (174,0,170,0,137,0,0,0,0,0,241,0,163,0,116,0,145,0,0,0,0,0,0,0,67,0,0,0,0,0,0,0,125,0,0,0,246,0,158,0,0,0,138,0,104,0,137,0,235,0,45,0,8,0,143,0,0,0,247,0,177,0,102,0,163,0,58,0,124,0,163,0,251,0,0,0,134,0,201,0,103,0,121,0,0,0,96,0,224,0,127,0,132,0,223,0,137,0,53,0,127,0,187,0,0,0,0,0,0,0,27,0,168,0,143,0,101,0,0,0,65,0,127,0,82,0,0,0,213,0,78,0,47,0,0,0,207,0,152,0,161,0,235,0,37,0,152,0,87,0,185,0,198,0,218,0,205,0,189,0,0,0,0,0,148,0,0,0,91,0,236,0,59,0,171,0,8,0,236,0,2,0,0,0,200,0,136,0,221,0,199,0,77,0,93,0,115,0,187,0,0,0,204,0,207,0,200,0,232,0,0,0,0,0,0,0,250,0,141,0,95,0,136,0,248,0,216,0,42,0,53,0,150,0,4,0,134,0,188,0,0,0,12,0,0,0,0,0,82,0,92,0,0,0,158,0,87,0,184,0,99,0,114,0,0,0,128,0,0,0,248,0,187,0,128,0,30,0,199,0,33,0,40,0,0,0,178,0,232,0,91,0,94,0,220,0,18,0,28,0,235,0,10,0,149,0,0,0,108,0,105,0,243,0,77,0,225,0,189,0,0,0,117,0,42,0,182,0,161,0,26,0,223,0,143,0,70,0,0,0,0,0,178,0,153,0,0,0,250,0,25,0,188,0,0,0,194,0,218,0,76,0,157,0,115,0,0,0,130,0,77,0,231,0,43,0,0,0,45,0,45,0,0,0,0,0,246,0,113,0,125,0,182,0,133,0,0,0,0,0,205,0,29,0,5,0,63,0,0,0,213,0,65,0,233,0,86,0,113,0,0,0,163,0,169,0,205,0,203,0,163,0,0,0,100,0,0,0,0,0,0,0,58,0,248,0,0,0,132,0,91,0,46,0,82,0,0,0,0,0,0,0,40,0,0,0,168,0,129,0,115,0,89,0,53,0,207,0,212,0,94,0,167,0,192,0,181,0,0,0,0,0,181,0,0,0,132,0,147,0,64,0,112,0,31,0,0,0,177,0,0,0,77,0,129,0,170,0,0,0,40,0,172,0,170,0,0,0,0,0,130,0,0,0,71,0,48,0,0,0,20,0,163,0,170,0,38,0,219,0,240,0,237,0,3,0,150,0,131,0,192,0,150,0,169,0,96,0,71,0,129,0,0,0,101,0,182,0,199,0,81,0,252,0,0,0,0,0,236,0,164,0,61,0,225,0,135,0,113,0,243,0,94,0,221,0,130,0,189,0,129,0,0,0,0,0,143,0,148,0,100,0,238,0,253,0,208,0,0,0,24,0,192,0,166,0,47,0,155,0,0,0,198,0,117,0,0,0,177,0,134,0,122,0,204,0,68,0,40,0,149,0,185,0,231,0,227,0,140,0,140,0,114,0,114,0,23,0,68,0,137,0,0,0,125,0,140,0,181,0,142,0,0,0,0,0,180,0,0,0,134,0,0,0,219,0,0,0,24,0,176,0,201,0,113,0,5,0,140,0,169,0,0,0,0,0,0,0,0,0,13,0,0,0,227,0,4,0,228,0,157,0,123,0,245,0,238,0,48,0,78,0,231,0,124,0,117,0,112,0,243,0,66,0,177,0,140,0,8,0,247,0,139,0,194,0,25,0,0,0,49,0,6,0,174,0,0,0,225,0,106,0,0,0,0,0,141,0,181,0,237,0,89,0,0,0,215,0,161,0,0,0,213,0,39,0,0,0,160,0,0,0,0,0,0,0,109,0,10,0,130,0,90,0,0,0,223,0,146,0,230,0,244,0,97,0,96,0,221,0,56,0,208,0,213,0,225,0,0,0,73,0,94,0,43,0,0,0,180,0,7,0,156,0,208,0,219,0,124,0,25,0,149,0,0,0,83,0,199,0,36,0,192,0,74,0,172,0,159,0,87,0,221,0,42,0,56,0,98,0,104,0,104,0,36,0,126,0,87,0,114,0,212,0,133,0,83,0,15,0,153,0,222,0,34,0,80,0,66,0,134,0,51,0,114,0,227,0,255,0,127,0,55,0,195,0,207,0,0,0,105,0,195,0,0,0,231,0,119,0,123,0,126,0,22,0,211,0,96,0,230,0,244,0,130,0,148,0,75,0,7,0,215,0,164,0,240,0,197,0,0,0,152,0,237,0,35,0,37,0,18,0,21,0,186,0,103,0,0,0,230,0,136,0,147,0,57,0,0,0,80,0,5,0,64,0,242,0,134,0,88,0,0,0,1,0,233,0,44,0,81,0,228,0,253,0,180,0,230,0,61,0,127,0,217,0,226,0,54,0,179,0,248,0,216,0,86,0,0,0,1,0,0,0,243,0,39,0,144,0,120,0,36,0,169,0,120,0,162,0,0,0,0,0,0,0,220,0,204,0,0,0,141,0,102,0,123,0,0,0,118,0,0,0,69,0,246,0,52,0,72,0,234,0,224,0,102,0,254,0,65,0,11,0,99,0,0,0,0,0,0,0,204,0,40,0,89,0,180,0,62,0,170,0,0,0,84,0,131,0,65,0,121,0,251,0,204,0,58,0,46,0,84,0,186,0,49,0,64,0,93,0,60,0,0,0,249,0,168,0,0,0,15,0,105,0,7,0,127,0,197,0,42,0,52,0,112,0,238,0,63,0,0,0,195,0,241,0,86,0,116,0,0,0,118,0,202,0,0,0,211,0,55,0,0,0,248,0,56,0,235,0,0,0,0,0,114,0,242,0,136,0,41,0,114,0,30,0,181,0,137,0,0,0,164,0,0,0,57,0,143,0,0,0,108,0,0,0,52,0,0,0,0,0,0,0,240,0,63,0,129,0,207,0,109,0,0,0,162,0,198,0,82,0,61,0);
signal scenario_full  : scenario_type := (174,31,170,31,137,31,137,30,137,29,241,31,163,31,116,31,145,31,145,30,145,29,145,28,67,31,67,30,67,29,67,28,125,31,125,30,246,31,158,31,158,30,138,31,104,31,137,31,235,31,45,31,8,31,143,31,143,30,247,31,177,31,102,31,163,31,58,31,124,31,163,31,251,31,251,30,134,31,201,31,103,31,121,31,121,30,96,31,224,31,127,31,132,31,223,31,137,31,53,31,127,31,187,31,187,30,187,29,187,28,27,31,168,31,143,31,101,31,101,30,65,31,127,31,82,31,82,30,213,31,78,31,47,31,47,30,207,31,152,31,161,31,235,31,37,31,152,31,87,31,185,31,198,31,218,31,205,31,189,31,189,30,189,29,148,31,148,30,91,31,236,31,59,31,171,31,8,31,236,31,2,31,2,30,200,31,136,31,221,31,199,31,77,31,93,31,115,31,187,31,187,30,204,31,207,31,200,31,232,31,232,30,232,29,232,28,250,31,141,31,95,31,136,31,248,31,216,31,42,31,53,31,150,31,4,31,134,31,188,31,188,30,12,31,12,30,12,29,82,31,92,31,92,30,158,31,87,31,184,31,99,31,114,31,114,30,128,31,128,30,248,31,187,31,128,31,30,31,199,31,33,31,40,31,40,30,178,31,232,31,91,31,94,31,220,31,18,31,28,31,235,31,10,31,149,31,149,30,108,31,105,31,243,31,77,31,225,31,189,31,189,30,117,31,42,31,182,31,161,31,26,31,223,31,143,31,70,31,70,30,70,29,178,31,153,31,153,30,250,31,25,31,188,31,188,30,194,31,218,31,76,31,157,31,115,31,115,30,130,31,77,31,231,31,43,31,43,30,45,31,45,31,45,30,45,29,246,31,113,31,125,31,182,31,133,31,133,30,133,29,205,31,29,31,5,31,63,31,63,30,213,31,65,31,233,31,86,31,113,31,113,30,163,31,169,31,205,31,203,31,163,31,163,30,100,31,100,30,100,29,100,28,58,31,248,31,248,30,132,31,91,31,46,31,82,31,82,30,82,29,82,28,40,31,40,30,168,31,129,31,115,31,89,31,53,31,207,31,212,31,94,31,167,31,192,31,181,31,181,30,181,29,181,31,181,30,132,31,147,31,64,31,112,31,31,31,31,30,177,31,177,30,77,31,129,31,170,31,170,30,40,31,172,31,170,31,170,30,170,29,130,31,130,30,71,31,48,31,48,30,20,31,163,31,170,31,38,31,219,31,240,31,237,31,3,31,150,31,131,31,192,31,150,31,169,31,96,31,71,31,129,31,129,30,101,31,182,31,199,31,81,31,252,31,252,30,252,29,236,31,164,31,61,31,225,31,135,31,113,31,243,31,94,31,221,31,130,31,189,31,129,31,129,30,129,29,143,31,148,31,100,31,238,31,253,31,208,31,208,30,24,31,192,31,166,31,47,31,155,31,155,30,198,31,117,31,117,30,177,31,134,31,122,31,204,31,68,31,40,31,149,31,185,31,231,31,227,31,140,31,140,31,114,31,114,31,23,31,68,31,137,31,137,30,125,31,140,31,181,31,142,31,142,30,142,29,180,31,180,30,134,31,134,30,219,31,219,30,24,31,176,31,201,31,113,31,5,31,140,31,169,31,169,30,169,29,169,28,169,27,13,31,13,30,227,31,4,31,228,31,157,31,123,31,245,31,238,31,48,31,78,31,231,31,124,31,117,31,112,31,243,31,66,31,177,31,140,31,8,31,247,31,139,31,194,31,25,31,25,30,49,31,6,31,174,31,174,30,225,31,106,31,106,30,106,29,141,31,181,31,237,31,89,31,89,30,215,31,161,31,161,30,213,31,39,31,39,30,160,31,160,30,160,29,160,28,109,31,10,31,130,31,90,31,90,30,223,31,146,31,230,31,244,31,97,31,96,31,221,31,56,31,208,31,213,31,225,31,225,30,73,31,94,31,43,31,43,30,180,31,7,31,156,31,208,31,219,31,124,31,25,31,149,31,149,30,83,31,199,31,36,31,192,31,74,31,172,31,159,31,87,31,221,31,42,31,56,31,98,31,104,31,104,31,36,31,126,31,87,31,114,31,212,31,133,31,83,31,15,31,153,31,222,31,34,31,80,31,66,31,134,31,51,31,114,31,227,31,255,31,127,31,55,31,195,31,207,31,207,30,105,31,195,31,195,30,231,31,119,31,123,31,126,31,22,31,211,31,96,31,230,31,244,31,130,31,148,31,75,31,7,31,215,31,164,31,240,31,197,31,197,30,152,31,237,31,35,31,37,31,18,31,21,31,186,31,103,31,103,30,230,31,136,31,147,31,57,31,57,30,80,31,5,31,64,31,242,31,134,31,88,31,88,30,1,31,233,31,44,31,81,31,228,31,253,31,180,31,230,31,61,31,127,31,217,31,226,31,54,31,179,31,248,31,216,31,86,31,86,30,1,31,1,30,243,31,39,31,144,31,120,31,36,31,169,31,120,31,162,31,162,30,162,29,162,28,220,31,204,31,204,30,141,31,102,31,123,31,123,30,118,31,118,30,69,31,246,31,52,31,72,31,234,31,224,31,102,31,254,31,65,31,11,31,99,31,99,30,99,29,99,28,204,31,40,31,89,31,180,31,62,31,170,31,170,30,84,31,131,31,65,31,121,31,251,31,204,31,58,31,46,31,84,31,186,31,49,31,64,31,93,31,60,31,60,30,249,31,168,31,168,30,15,31,105,31,7,31,127,31,197,31,42,31,52,31,112,31,238,31,63,31,63,30,195,31,241,31,86,31,116,31,116,30,118,31,202,31,202,30,211,31,55,31,55,30,248,31,56,31,235,31,235,30,235,29,114,31,242,31,136,31,41,31,114,31,30,31,181,31,137,31,137,30,164,31,164,30,57,31,143,31,143,30,108,31,108,30,52,31,52,30,52,29,52,28,240,31,63,31,129,31,207,31,109,31,109,30,162,31,198,31,82,31,61,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
