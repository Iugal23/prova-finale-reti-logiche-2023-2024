-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_984 is
end project_tb_984;

architecture project_tb_arch_984 of project_tb_984 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 746;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (9,0,0,0,52,0,0,0,141,0,0,0,29,0,88,0,127,0,142,0,0,0,36,0,29,0,229,0,8,0,72,0,184,0,196,0,33,0,159,0,0,0,251,0,31,0,0,0,4,0,182,0,35,0,117,0,116,0,255,0,0,0,0,0,0,0,37,0,0,0,17,0,118,0,59,0,225,0,0,0,195,0,251,0,214,0,95,0,165,0,152,0,115,0,56,0,24,0,150,0,235,0,66,0,195,0,164,0,0,0,93,0,218,0,157,0,72,0,223,0,44,0,166,0,5,0,9,0,0,0,40,0,76,0,224,0,173,0,0,0,95,0,43,0,161,0,237,0,231,0,0,0,0,0,149,0,192,0,0,0,26,0,164,0,247,0,23,0,195,0,0,0,40,0,135,0,174,0,205,0,43,0,42,0,0,0,95,0,72,0,103,0,169,0,187,0,232,0,143,0,204,0,179,0,117,0,50,0,163,0,151,0,242,0,157,0,214,0,198,0,179,0,135,0,237,0,58,0,33,0,0,0,184,0,19,0,103,0,197,0,147,0,120,0,47,0,69,0,150,0,5,0,197,0,231,0,205,0,192,0,146,0,46,0,15,0,32,0,180,0,235,0,230,0,168,0,0,0,165,0,0,0,108,0,161,0,230,0,223,0,210,0,245,0,196,0,85,0,158,0,0,0,176,0,158,0,79,0,226,0,158,0,129,0,109,0,0,0,0,0,109,0,0,0,0,0,6,0,27,0,173,0,68,0,132,0,132,0,154,0,151,0,0,0,220,0,0,0,132,0,76,0,0,0,23,0,74,0,34,0,216,0,78,0,3,0,0,0,12,0,10,0,90,0,162,0,88,0,75,0,0,0,204,0,231,0,0,0,237,0,230,0,129,0,246,0,126,0,133,0,219,0,141,0,164,0,0,0,81,0,85,0,135,0,105,0,3,0,0,0,0,0,235,0,55,0,0,0,126,0,2,0,181,0,161,0,129,0,231,0,42,0,182,0,249,0,31,0,0,0,172,0,141,0,172,0,59,0,0,0,178,0,109,0,157,0,58,0,242,0,21,0,122,0,0,0,152,0,194,0,0,0,218,0,239,0,156,0,0,0,0,0,108,0,0,0,219,0,88,0,221,0,35,0,15,0,3,0,22,0,0,0,254,0,194,0,235,0,118,0,0,0,117,0,243,0,138,0,81,0,78,0,66,0,81,0,224,0,0,0,198,0,57,0,45,0,200,0,57,0,9,0,136,0,197,0,148,0,1,0,85,0,159,0,0,0,127,0,0,0,36,0,195,0,102,0,0,0,0,0,243,0,73,0,188,0,0,0,136,0,52,0,103,0,161,0,22,0,67,0,74,0,32,0,76,0,217,0,55,0,225,0,0,0,0,0,121,0,91,0,255,0,14,0,60,0,197,0,60,0,220,0,43,0,32,0,126,0,51,0,20,0,189,0,0,0,204,0,229,0,149,0,190,0,0,0,0,0,0,0,0,0,69,0,75,0,151,0,127,0,5,0,37,0,0,0,154,0,61,0,60,0,169,0,144,0,198,0,202,0,247,0,255,0,248,0,13,0,0,0,19,0,55,0,227,0,184,0,71,0,0,0,74,0,59,0,70,0,96,0,54,0,118,0,0,0,174,0,7,0,32,0,58,0,16,0,127,0,224,0,148,0,137,0,146,0,28,0,0,0,122,0,77,0,177,0,242,0,227,0,133,0,196,0,13,0,0,0,167,0,0,0,0,0,251,0,179,0,244,0,0,0,25,0,246,0,87,0,0,0,46,0,94,0,161,0,0,0,78,0,163,0,116,0,193,0,38,0,245,0,0,0,81,0,159,0,0,0,8,0,16,0,0,0,127,0,0,0,0,0,174,0,233,0,77,0,0,0,120,0,251,0,216,0,195,0,114,0,143,0,229,0,113,0,224,0,0,0,116,0,56,0,0,0,0,0,0,0,157,0,245,0,91,0,241,0,244,0,224,0,0,0,81,0,239,0,19,0,186,0,222,0,4,0,0,0,135,0,0,0,144,0,238,0,30,0,228,0,159,0,253,0,6,0,111,0,0,0,0,0,228,0,244,0,187,0,135,0,0,0,80,0,200,0,234,0,0,0,218,0,0,0,250,0,137,0,204,0,220,0,0,0,0,0,68,0,26,0,144,0,76,0,170,0,59,0,5,0,197,0,239,0,0,0,251,0,205,0,199,0,0,0,117,0,38,0,117,0,73,0,64,0,33,0,197,0,57,0,115,0,0,0,11,0,240,0,233,0,52,0,214,0,191,0,176,0,219,0,0,0,125,0,24,0,0,0,32,0,225,0,158,0,199,0,0,0,26,0,0,0,0,0,255,0,60,0,171,0,44,0,179,0,137,0,161,0,188,0,110,0,26,0,0,0,243,0,110,0,101,0,220,0,82,0,28,0,126,0,105,0,234,0,97,0,198,0,31,0,87,0,10,0,193,0,0,0,0,0,0,0,135,0,47,0,171,0,0,0,112,0,247,0,71,0,146,0,59,0,190,0,186,0,10,0,151,0,0,0,81,0,114,0,51,0,160,0,0,0,120,0,193,0,101,0,2,0,162,0,0,0,239,0,189,0,197,0,16,0,0,0,79,0,57,0,3,0,33,0,11,0,221,0,218,0,185,0,126,0,0,0,117,0,154,0,36,0,150,0,0,0,239,0,56,0,201,0,245,0,3,0,0,0,161,0,0,0,120,0,229,0,0,0,163,0,34,0,101,0,0,0,0,0,226,0,150,0,176,0,166,0,137,0,62,0,124,0,10,0,0,0,0,0,0,0,230,0,116,0,156,0,31,0,136,0,128,0,120,0,182,0,68,0,175,0,0,0,107,0,0,0,1,0,164,0,81,0,0,0,221,0,211,0,7,0,199,0,180,0,225,0,227,0,161,0,20,0,83,0,104,0,180,0,34,0,176,0,250,0,73,0,0,0,134,0,133,0,50,0,14,0,150,0,197,0,0,0,128,0,25,0,248,0,128,0,57,0,106,0,189,0,0,0,134,0,28,0,29,0,0,0,226,0,49,0,96,0,143,0,72,0,0,0,229,0,27,0,201,0,195,0,0,0,126,0,22,0,90,0,0,0,0,0,0,0,84,0,95,0,61,0,143,0,66,0,208,0,48,0,196,0,0,0,239,0,24,0,56,0,154,0,133,0,0,0,0,0,119,0,220,0,40,0,0,0,1,0,184,0,51,0,63,0,29,0,130,0,138,0,237,0,0,0,47,0,174,0,250,0,86,0,15,0,185,0,79,0,120,0,185,0,144,0,215,0,50,0,162,0,228,0,241,0,127,0,143,0,255,0,64,0,123,0,160,0,184,0,14,0,117,0,0,0);
signal scenario_full  : scenario_type := (9,31,9,30,52,31,52,30,141,31,141,30,29,31,88,31,127,31,142,31,142,30,36,31,29,31,229,31,8,31,72,31,184,31,196,31,33,31,159,31,159,30,251,31,31,31,31,30,4,31,182,31,35,31,117,31,116,31,255,31,255,30,255,29,255,28,37,31,37,30,17,31,118,31,59,31,225,31,225,30,195,31,251,31,214,31,95,31,165,31,152,31,115,31,56,31,24,31,150,31,235,31,66,31,195,31,164,31,164,30,93,31,218,31,157,31,72,31,223,31,44,31,166,31,5,31,9,31,9,30,40,31,76,31,224,31,173,31,173,30,95,31,43,31,161,31,237,31,231,31,231,30,231,29,149,31,192,31,192,30,26,31,164,31,247,31,23,31,195,31,195,30,40,31,135,31,174,31,205,31,43,31,42,31,42,30,95,31,72,31,103,31,169,31,187,31,232,31,143,31,204,31,179,31,117,31,50,31,163,31,151,31,242,31,157,31,214,31,198,31,179,31,135,31,237,31,58,31,33,31,33,30,184,31,19,31,103,31,197,31,147,31,120,31,47,31,69,31,150,31,5,31,197,31,231,31,205,31,192,31,146,31,46,31,15,31,32,31,180,31,235,31,230,31,168,31,168,30,165,31,165,30,108,31,161,31,230,31,223,31,210,31,245,31,196,31,85,31,158,31,158,30,176,31,158,31,79,31,226,31,158,31,129,31,109,31,109,30,109,29,109,31,109,30,109,29,6,31,27,31,173,31,68,31,132,31,132,31,154,31,151,31,151,30,220,31,220,30,132,31,76,31,76,30,23,31,74,31,34,31,216,31,78,31,3,31,3,30,12,31,10,31,90,31,162,31,88,31,75,31,75,30,204,31,231,31,231,30,237,31,230,31,129,31,246,31,126,31,133,31,219,31,141,31,164,31,164,30,81,31,85,31,135,31,105,31,3,31,3,30,3,29,235,31,55,31,55,30,126,31,2,31,181,31,161,31,129,31,231,31,42,31,182,31,249,31,31,31,31,30,172,31,141,31,172,31,59,31,59,30,178,31,109,31,157,31,58,31,242,31,21,31,122,31,122,30,152,31,194,31,194,30,218,31,239,31,156,31,156,30,156,29,108,31,108,30,219,31,88,31,221,31,35,31,15,31,3,31,22,31,22,30,254,31,194,31,235,31,118,31,118,30,117,31,243,31,138,31,81,31,78,31,66,31,81,31,224,31,224,30,198,31,57,31,45,31,200,31,57,31,9,31,136,31,197,31,148,31,1,31,85,31,159,31,159,30,127,31,127,30,36,31,195,31,102,31,102,30,102,29,243,31,73,31,188,31,188,30,136,31,52,31,103,31,161,31,22,31,67,31,74,31,32,31,76,31,217,31,55,31,225,31,225,30,225,29,121,31,91,31,255,31,14,31,60,31,197,31,60,31,220,31,43,31,32,31,126,31,51,31,20,31,189,31,189,30,204,31,229,31,149,31,190,31,190,30,190,29,190,28,190,27,69,31,75,31,151,31,127,31,5,31,37,31,37,30,154,31,61,31,60,31,169,31,144,31,198,31,202,31,247,31,255,31,248,31,13,31,13,30,19,31,55,31,227,31,184,31,71,31,71,30,74,31,59,31,70,31,96,31,54,31,118,31,118,30,174,31,7,31,32,31,58,31,16,31,127,31,224,31,148,31,137,31,146,31,28,31,28,30,122,31,77,31,177,31,242,31,227,31,133,31,196,31,13,31,13,30,167,31,167,30,167,29,251,31,179,31,244,31,244,30,25,31,246,31,87,31,87,30,46,31,94,31,161,31,161,30,78,31,163,31,116,31,193,31,38,31,245,31,245,30,81,31,159,31,159,30,8,31,16,31,16,30,127,31,127,30,127,29,174,31,233,31,77,31,77,30,120,31,251,31,216,31,195,31,114,31,143,31,229,31,113,31,224,31,224,30,116,31,56,31,56,30,56,29,56,28,157,31,245,31,91,31,241,31,244,31,224,31,224,30,81,31,239,31,19,31,186,31,222,31,4,31,4,30,135,31,135,30,144,31,238,31,30,31,228,31,159,31,253,31,6,31,111,31,111,30,111,29,228,31,244,31,187,31,135,31,135,30,80,31,200,31,234,31,234,30,218,31,218,30,250,31,137,31,204,31,220,31,220,30,220,29,68,31,26,31,144,31,76,31,170,31,59,31,5,31,197,31,239,31,239,30,251,31,205,31,199,31,199,30,117,31,38,31,117,31,73,31,64,31,33,31,197,31,57,31,115,31,115,30,11,31,240,31,233,31,52,31,214,31,191,31,176,31,219,31,219,30,125,31,24,31,24,30,32,31,225,31,158,31,199,31,199,30,26,31,26,30,26,29,255,31,60,31,171,31,44,31,179,31,137,31,161,31,188,31,110,31,26,31,26,30,243,31,110,31,101,31,220,31,82,31,28,31,126,31,105,31,234,31,97,31,198,31,31,31,87,31,10,31,193,31,193,30,193,29,193,28,135,31,47,31,171,31,171,30,112,31,247,31,71,31,146,31,59,31,190,31,186,31,10,31,151,31,151,30,81,31,114,31,51,31,160,31,160,30,120,31,193,31,101,31,2,31,162,31,162,30,239,31,189,31,197,31,16,31,16,30,79,31,57,31,3,31,33,31,11,31,221,31,218,31,185,31,126,31,126,30,117,31,154,31,36,31,150,31,150,30,239,31,56,31,201,31,245,31,3,31,3,30,161,31,161,30,120,31,229,31,229,30,163,31,34,31,101,31,101,30,101,29,226,31,150,31,176,31,166,31,137,31,62,31,124,31,10,31,10,30,10,29,10,28,230,31,116,31,156,31,31,31,136,31,128,31,120,31,182,31,68,31,175,31,175,30,107,31,107,30,1,31,164,31,81,31,81,30,221,31,211,31,7,31,199,31,180,31,225,31,227,31,161,31,20,31,83,31,104,31,180,31,34,31,176,31,250,31,73,31,73,30,134,31,133,31,50,31,14,31,150,31,197,31,197,30,128,31,25,31,248,31,128,31,57,31,106,31,189,31,189,30,134,31,28,31,29,31,29,30,226,31,49,31,96,31,143,31,72,31,72,30,229,31,27,31,201,31,195,31,195,30,126,31,22,31,90,31,90,30,90,29,90,28,84,31,95,31,61,31,143,31,66,31,208,31,48,31,196,31,196,30,239,31,24,31,56,31,154,31,133,31,133,30,133,29,119,31,220,31,40,31,40,30,1,31,184,31,51,31,63,31,29,31,130,31,138,31,237,31,237,30,47,31,174,31,250,31,86,31,15,31,185,31,79,31,120,31,185,31,144,31,215,31,50,31,162,31,228,31,241,31,127,31,143,31,255,31,64,31,123,31,160,31,184,31,14,31,117,31,117,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
