-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_32 is
end project_tb_32;

architecture project_tb_arch_32 of project_tb_32 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 951;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (167,0,71,0,48,0,138,0,83,0,0,0,75,0,0,0,0,0,133,0,0,0,245,0,246,0,19,0,85,0,5,0,235,0,187,0,154,0,43,0,39,0,137,0,152,0,85,0,34,0,75,0,193,0,206,0,158,0,77,0,249,0,248,0,82,0,231,0,6,0,149,0,240,0,88,0,114,0,0,0,0,0,36,0,107,0,55,0,0,0,155,0,215,0,35,0,71,0,225,0,140,0,130,0,127,0,54,0,207,0,194,0,194,0,71,0,155,0,63,0,254,0,23,0,212,0,178,0,19,0,182,0,71,0,38,0,117,0,153,0,36,0,158,0,157,0,0,0,140,0,0,0,251,0,238,0,126,0,218,0,17,0,158,0,179,0,221,0,151,0,186,0,220,0,0,0,251,0,0,0,91,0,10,0,38,0,64,0,0,0,27,0,227,0,99,0,0,0,157,0,107,0,159,0,221,0,92,0,201,0,0,0,214,0,221,0,0,0,101,0,0,0,72,0,0,0,0,0,227,0,0,0,206,0,213,0,182,0,71,0,124,0,0,0,219,0,234,0,38,0,0,0,128,0,20,0,5,0,0,0,14,0,25,0,0,0,28,0,74,0,0,0,104,0,236,0,80,0,74,0,202,0,133,0,46,0,176,0,0,0,1,0,38,0,108,0,234,0,237,0,47,0,0,0,167,0,65,0,0,0,202,0,241,0,66,0,134,0,0,0,230,0,0,0,91,0,56,0,0,0,0,0,183,0,136,0,71,0,0,0,0,0,175,0,88,0,19,0,197,0,0,0,197,0,31,0,191,0,200,0,139,0,97,0,232,0,167,0,246,0,47,0,197,0,58,0,254,0,182,0,0,0,0,0,140,0,146,0,0,0,58,0,205,0,134,0,88,0,0,0,29,0,84,0,16,0,246,0,252,0,242,0,51,0,86,0,14,0,247,0,179,0,131,0,140,0,204,0,147,0,116,0,213,0,0,0,139,0,138,0,170,0,147,0,98,0,5,0,249,0,0,0,250,0,168,0,238,0,141,0,126,0,8,0,219,0,0,0,172,0,167,0,82,0,248,0,16,0,241,0,161,0,248,0,0,0,128,0,87,0,15,0,187,0,0,0,0,0,0,0,195,0,52,0,160,0,239,0,180,0,0,0,61,0,185,0,207,0,101,0,185,0,57,0,77,0,0,0,69,0,161,0,206,0,154,0,0,0,127,0,35,0,224,0,0,0,70,0,128,0,233,0,161,0,218,0,158,0,127,0,0,0,230,0,0,0,0,0,236,0,11,0,143,0,0,0,0,0,214,0,66,0,240,0,28,0,124,0,0,0,38,0,165,0,8,0,86,0,153,0,201,0,247,0,245,0,33,0,0,0,57,0,246,0,19,0,122,0,0,0,0,0,43,0,108,0,218,0,21,0,244,0,159,0,0,0,0,0,0,0,0,0,19,0,170,0,49,0,78,0,67,0,82,0,57,0,0,0,181,0,13,0,196,0,35,0,0,0,124,0,12,0,45,0,202,0,130,0,0,0,59,0,44,0,0,0,0,0,9,0,72,0,0,0,168,0,217,0,35,0,57,0,50,0,151,0,197,0,188,0,79,0,72,0,237,0,0,0,0,0,68,0,125,0,217,0,34,0,160,0,80,0,0,0,254,0,0,0,43,0,0,0,15,0,63,0,0,0,149,0,158,0,0,0,170,0,35,0,147,0,131,0,113,0,91,0,37,0,0,0,116,0,56,0,249,0,0,0,0,0,58,0,166,0,173,0,12,0,221,0,217,0,118,0,28,0,0,0,254,0,41,0,183,0,207,0,47,0,243,0,0,0,74,0,0,0,80,0,197,0,173,0,29,0,0,0,222,0,197,0,105,0,231,0,238,0,0,0,83,0,76,0,49,0,24,0,107,0,171,0,200,0,61,0,79,0,25,0,236,0,0,0,23,0,147,0,112,0,238,0,17,0,84,0,206,0,144,0,149,0,107,0,73,0,112,0,188,0,113,0,48,0,185,0,0,0,107,0,77,0,225,0,0,0,13,0,0,0,210,0,159,0,0,0,0,0,0,0,17,0,123,0,236,0,118,0,8,0,157,0,169,0,224,0,26,0,31,0,74,0,33,0,238,0,44,0,236,0,31,0,0,0,98,0,117,0,115,0,20,0,58,0,180,0,0,0,129,0,15,0,0,0,78,0,36,0,252,0,192,0,0,0,216,0,0,0,160,0,0,0,204,0,0,0,220,0,182,0,164,0,76,0,0,0,178,0,201,0,0,0,161,0,230,0,250,0,0,0,133,0,11,0,209,0,10,0,218,0,49,0,109,0,45,0,24,0,149,0,98,0,133,0,167,0,0,0,0,0,57,0,0,0,182,0,0,0,113,0,47,0,54,0,183,0,12,0,71,0,232,0,108,0,168,0,173,0,0,0,109,0,78,0,4,0,0,0,150,0,173,0,12,0,230,0,158,0,65,0,183,0,153,0,209,0,230,0,32,0,43,0,0,0,104,0,161,0,130,0,12,0,2,0,0,0,254,0,6,0,0,0,67,0,159,0,19,0,180,0,248,0,0,0,207,0,115,0,111,0,253,0,229,0,0,0,241,0,86,0,13,0,137,0,181,0,38,0,0,0,0,0,92,0,0,0,198,0,239,0,72,0,108,0,201,0,123,0,4,0,166,0,209,0,207,0,0,0,17,0,0,0,237,0,179,0,112,0,192,0,0,0,114,0,232,0,146,0,251,0,1,0,241,0,205,0,31,0,243,0,81,0,114,0,235,0,64,0,0,0,212,0,180,0,148,0,48,0,182,0,40,0,0,0,0,0,159,0,142,0,105,0,8,0,247,0,195,0,45,0,0,0,0,0,96,0,76,0,93,0,158,0,41,0,187,0,0,0,41,0,238,0,186,0,168,0,118,0,153,0,143,0,194,0,27,0,0,0,0,0,151,0,89,0,175,0,65,0,229,0,147,0,199,0,40,0,107,0,75,0,0,0,169,0,0,0,214,0,153,0,0,0,246,0,190,0,145,0,122,0,0,0,201,0,178,0,110,0,104,0,172,0,210,0,174,0,194,0,107,0,4,0,46,0,243,0,241,0,138,0,0,0,0,0,50,0,16,0,0,0,43,0,226,0,46,0,141,0,175,0,182,0,84,0,140,0,0,0,61,0,123,0,216,0,0,0,19,0,219,0,152,0,168,0,65,0,167,0,150,0,189,0,162,0,109,0,171,0,108,0,149,0,0,0,50,0,107,0,161,0,0,0,112,0,132,0,38,0,26,0,202,0,75,0,122,0,255,0,229,0,0,0,117,0,125,0,49,0,38,0,162,0,106,0,0,0,0,0,168,0,0,0,62,0,74,0,55,0,62,0,142,0,234,0,18,0,211,0,194,0,31,0,81,0,0,0,227,0,235,0,150,0,196,0,99,0,179,0,181,0,234,0,0,0,201,0,249,0,131,0,0,0,99,0,70,0,0,0,255,0,154,0,108,0,131,0,197,0,0,0,0,0,0,0,180,0,176,0,162,0,159,0,0,0,83,0,49,0,203,0,2,0,37,0,230,0,226,0,198,0,15,0,18,0,0,0,59,0,116,0,61,0,196,0,130,0,89,0,218,0,101,0,144,0,65,0,0,0,30,0,139,0,227,0,172,0,0,0,54,0,237,0,100,0,71,0,102,0,0,0,90,0,163,0,30,0,45,0,0,0,234,0,2,0,114,0,239,0,107,0,74,0,197,0,151,0,153,0,84,0,187,0,37,0,225,0,62,0,117,0,101,0,22,0,0,0,0,0,171,0,150,0,215,0,0,0,164,0,172,0,0,0,216,0,218,0,139,0,251,0,0,0,28,0,0,0,0,0,48,0,155,0,182,0,138,0,213,0,104,0,9,0,18,0,243,0,70,0,0,0,147,0,253,0,131,0,56,0,139,0,165,0,0,0,0,0,0,0,94,0,0,0,0,0,123,0,0,0,171,0,176,0,123,0,69,0,157,0,67,0,0,0,66,0,191,0,230,0,101,0,179,0,28,0,212,0,105,0,109,0,157,0,85,0,136,0,100,0,88,0,117,0,97,0,0,0,38,0,0,0,126,0,0,0,0,0,65,0,228,0,19,0,145,0,98,0,234,0,150,0,225,0,0,0,223,0,0,0,56,0,185,0,180,0,198,0,150,0,167,0,124,0,179,0,144,0,86,0,239,0,90,0,28,0,0,0,151,0,136,0,29,0,75,0,187,0,167,0,136,0,199,0,0,0,83,0,73,0,11,0,196,0,0,0);
signal scenario_full  : scenario_type := (167,31,71,31,48,31,138,31,83,31,83,30,75,31,75,30,75,29,133,31,133,30,245,31,246,31,19,31,85,31,5,31,235,31,187,31,154,31,43,31,39,31,137,31,152,31,85,31,34,31,75,31,193,31,206,31,158,31,77,31,249,31,248,31,82,31,231,31,6,31,149,31,240,31,88,31,114,31,114,30,114,29,36,31,107,31,55,31,55,30,155,31,215,31,35,31,71,31,225,31,140,31,130,31,127,31,54,31,207,31,194,31,194,31,71,31,155,31,63,31,254,31,23,31,212,31,178,31,19,31,182,31,71,31,38,31,117,31,153,31,36,31,158,31,157,31,157,30,140,31,140,30,251,31,238,31,126,31,218,31,17,31,158,31,179,31,221,31,151,31,186,31,220,31,220,30,251,31,251,30,91,31,10,31,38,31,64,31,64,30,27,31,227,31,99,31,99,30,157,31,107,31,159,31,221,31,92,31,201,31,201,30,214,31,221,31,221,30,101,31,101,30,72,31,72,30,72,29,227,31,227,30,206,31,213,31,182,31,71,31,124,31,124,30,219,31,234,31,38,31,38,30,128,31,20,31,5,31,5,30,14,31,25,31,25,30,28,31,74,31,74,30,104,31,236,31,80,31,74,31,202,31,133,31,46,31,176,31,176,30,1,31,38,31,108,31,234,31,237,31,47,31,47,30,167,31,65,31,65,30,202,31,241,31,66,31,134,31,134,30,230,31,230,30,91,31,56,31,56,30,56,29,183,31,136,31,71,31,71,30,71,29,175,31,88,31,19,31,197,31,197,30,197,31,31,31,191,31,200,31,139,31,97,31,232,31,167,31,246,31,47,31,197,31,58,31,254,31,182,31,182,30,182,29,140,31,146,31,146,30,58,31,205,31,134,31,88,31,88,30,29,31,84,31,16,31,246,31,252,31,242,31,51,31,86,31,14,31,247,31,179,31,131,31,140,31,204,31,147,31,116,31,213,31,213,30,139,31,138,31,170,31,147,31,98,31,5,31,249,31,249,30,250,31,168,31,238,31,141,31,126,31,8,31,219,31,219,30,172,31,167,31,82,31,248,31,16,31,241,31,161,31,248,31,248,30,128,31,87,31,15,31,187,31,187,30,187,29,187,28,195,31,52,31,160,31,239,31,180,31,180,30,61,31,185,31,207,31,101,31,185,31,57,31,77,31,77,30,69,31,161,31,206,31,154,31,154,30,127,31,35,31,224,31,224,30,70,31,128,31,233,31,161,31,218,31,158,31,127,31,127,30,230,31,230,30,230,29,236,31,11,31,143,31,143,30,143,29,214,31,66,31,240,31,28,31,124,31,124,30,38,31,165,31,8,31,86,31,153,31,201,31,247,31,245,31,33,31,33,30,57,31,246,31,19,31,122,31,122,30,122,29,43,31,108,31,218,31,21,31,244,31,159,31,159,30,159,29,159,28,159,27,19,31,170,31,49,31,78,31,67,31,82,31,57,31,57,30,181,31,13,31,196,31,35,31,35,30,124,31,12,31,45,31,202,31,130,31,130,30,59,31,44,31,44,30,44,29,9,31,72,31,72,30,168,31,217,31,35,31,57,31,50,31,151,31,197,31,188,31,79,31,72,31,237,31,237,30,237,29,68,31,125,31,217,31,34,31,160,31,80,31,80,30,254,31,254,30,43,31,43,30,15,31,63,31,63,30,149,31,158,31,158,30,170,31,35,31,147,31,131,31,113,31,91,31,37,31,37,30,116,31,56,31,249,31,249,30,249,29,58,31,166,31,173,31,12,31,221,31,217,31,118,31,28,31,28,30,254,31,41,31,183,31,207,31,47,31,243,31,243,30,74,31,74,30,80,31,197,31,173,31,29,31,29,30,222,31,197,31,105,31,231,31,238,31,238,30,83,31,76,31,49,31,24,31,107,31,171,31,200,31,61,31,79,31,25,31,236,31,236,30,23,31,147,31,112,31,238,31,17,31,84,31,206,31,144,31,149,31,107,31,73,31,112,31,188,31,113,31,48,31,185,31,185,30,107,31,77,31,225,31,225,30,13,31,13,30,210,31,159,31,159,30,159,29,159,28,17,31,123,31,236,31,118,31,8,31,157,31,169,31,224,31,26,31,31,31,74,31,33,31,238,31,44,31,236,31,31,31,31,30,98,31,117,31,115,31,20,31,58,31,180,31,180,30,129,31,15,31,15,30,78,31,36,31,252,31,192,31,192,30,216,31,216,30,160,31,160,30,204,31,204,30,220,31,182,31,164,31,76,31,76,30,178,31,201,31,201,30,161,31,230,31,250,31,250,30,133,31,11,31,209,31,10,31,218,31,49,31,109,31,45,31,24,31,149,31,98,31,133,31,167,31,167,30,167,29,57,31,57,30,182,31,182,30,113,31,47,31,54,31,183,31,12,31,71,31,232,31,108,31,168,31,173,31,173,30,109,31,78,31,4,31,4,30,150,31,173,31,12,31,230,31,158,31,65,31,183,31,153,31,209,31,230,31,32,31,43,31,43,30,104,31,161,31,130,31,12,31,2,31,2,30,254,31,6,31,6,30,67,31,159,31,19,31,180,31,248,31,248,30,207,31,115,31,111,31,253,31,229,31,229,30,241,31,86,31,13,31,137,31,181,31,38,31,38,30,38,29,92,31,92,30,198,31,239,31,72,31,108,31,201,31,123,31,4,31,166,31,209,31,207,31,207,30,17,31,17,30,237,31,179,31,112,31,192,31,192,30,114,31,232,31,146,31,251,31,1,31,241,31,205,31,31,31,243,31,81,31,114,31,235,31,64,31,64,30,212,31,180,31,148,31,48,31,182,31,40,31,40,30,40,29,159,31,142,31,105,31,8,31,247,31,195,31,45,31,45,30,45,29,96,31,76,31,93,31,158,31,41,31,187,31,187,30,41,31,238,31,186,31,168,31,118,31,153,31,143,31,194,31,27,31,27,30,27,29,151,31,89,31,175,31,65,31,229,31,147,31,199,31,40,31,107,31,75,31,75,30,169,31,169,30,214,31,153,31,153,30,246,31,190,31,145,31,122,31,122,30,201,31,178,31,110,31,104,31,172,31,210,31,174,31,194,31,107,31,4,31,46,31,243,31,241,31,138,31,138,30,138,29,50,31,16,31,16,30,43,31,226,31,46,31,141,31,175,31,182,31,84,31,140,31,140,30,61,31,123,31,216,31,216,30,19,31,219,31,152,31,168,31,65,31,167,31,150,31,189,31,162,31,109,31,171,31,108,31,149,31,149,30,50,31,107,31,161,31,161,30,112,31,132,31,38,31,26,31,202,31,75,31,122,31,255,31,229,31,229,30,117,31,125,31,49,31,38,31,162,31,106,31,106,30,106,29,168,31,168,30,62,31,74,31,55,31,62,31,142,31,234,31,18,31,211,31,194,31,31,31,81,31,81,30,227,31,235,31,150,31,196,31,99,31,179,31,181,31,234,31,234,30,201,31,249,31,131,31,131,30,99,31,70,31,70,30,255,31,154,31,108,31,131,31,197,31,197,30,197,29,197,28,180,31,176,31,162,31,159,31,159,30,83,31,49,31,203,31,2,31,37,31,230,31,226,31,198,31,15,31,18,31,18,30,59,31,116,31,61,31,196,31,130,31,89,31,218,31,101,31,144,31,65,31,65,30,30,31,139,31,227,31,172,31,172,30,54,31,237,31,100,31,71,31,102,31,102,30,90,31,163,31,30,31,45,31,45,30,234,31,2,31,114,31,239,31,107,31,74,31,197,31,151,31,153,31,84,31,187,31,37,31,225,31,62,31,117,31,101,31,22,31,22,30,22,29,171,31,150,31,215,31,215,30,164,31,172,31,172,30,216,31,218,31,139,31,251,31,251,30,28,31,28,30,28,29,48,31,155,31,182,31,138,31,213,31,104,31,9,31,18,31,243,31,70,31,70,30,147,31,253,31,131,31,56,31,139,31,165,31,165,30,165,29,165,28,94,31,94,30,94,29,123,31,123,30,171,31,176,31,123,31,69,31,157,31,67,31,67,30,66,31,191,31,230,31,101,31,179,31,28,31,212,31,105,31,109,31,157,31,85,31,136,31,100,31,88,31,117,31,97,31,97,30,38,31,38,30,126,31,126,30,126,29,65,31,228,31,19,31,145,31,98,31,234,31,150,31,225,31,225,30,223,31,223,30,56,31,185,31,180,31,198,31,150,31,167,31,124,31,179,31,144,31,86,31,239,31,90,31,28,31,28,30,151,31,136,31,29,31,75,31,187,31,167,31,136,31,199,31,199,30,83,31,73,31,11,31,196,31,196,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
