-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_375 is
end project_tb_375;

architecture project_tb_arch_375 of project_tb_375 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 697;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (105,0,20,0,123,0,152,0,19,0,0,0,178,0,88,0,48,0,106,0,156,0,0,0,175,0,16,0,9,0,179,0,216,0,0,0,86,0,154,0,41,0,0,0,49,0,134,0,51,0,216,0,145,0,58,0,0,0,0,0,113,0,4,0,0,0,241,0,233,0,0,0,8,0,9,0,138,0,129,0,113,0,247,0,184,0,113,0,144,0,0,0,185,0,26,0,38,0,63,0,175,0,12,0,251,0,127,0,42,0,150,0,71,0,134,0,0,0,195,0,210,0,0,0,231,0,0,0,0,0,176,0,246,0,21,0,14,0,168,0,0,0,234,0,0,0,31,0,241,0,76,0,83,0,91,0,217,0,123,0,0,0,132,0,0,0,0,0,0,0,114,0,29,0,212,0,203,0,85,0,203,0,29,0,0,0,251,0,220,0,0,0,159,0,220,0,0,0,89,0,0,0,176,0,76,0,0,0,41,0,0,0,138,0,101,0,200,0,127,0,252,0,0,0,32,0,170,0,120,0,0,0,66,0,0,0,77,0,68,0,0,0,134,0,0,0,173,0,166,0,41,0,134,0,0,0,73,0,50,0,111,0,19,0,229,0,7,0,125,0,9,0,173,0,127,0,161,0,146,0,0,0,0,0,15,0,0,0,94,0,0,0,92,0,0,0,198,0,162,0,0,0,11,0,231,0,251,0,105,0,154,0,0,0,0,0,0,0,82,0,6,0,201,0,71,0,223,0,224,0,0,0,14,0,52,0,132,0,107,0,101,0,23,0,0,0,170,0,172,0,0,0,25,0,144,0,186,0,220,0,133,0,17,0,46,0,32,0,195,0,100,0,233,0,0,0,131,0,6,0,190,0,85,0,105,0,74,0,112,0,211,0,196,0,230,0,68,0,127,0,142,0,204,0,235,0,12,0,0,0,0,0,188,0,175,0,19,0,141,0,149,0,88,0,31,0,229,0,84,0,230,0,20,0,0,0,175,0,42,0,165,0,4,0,153,0,203,0,235,0,161,0,179,0,0,0,222,0,44,0,109,0,56,0,46,0,166,0,135,0,0,0,0,0,234,0,0,0,0,0,4,0,19,0,132,0,0,0,0,0,139,0,65,0,169,0,118,0,84,0,28,0,100,0,154,0,17,0,14,0,175,0,0,0,0,0,0,0,0,0,146,0,255,0,167,0,98,0,218,0,37,0,110,0,0,0,88,0,196,0,57,0,0,0,0,0,0,0,228,0,148,0,14,0,27,0,149,0,129,0,0,0,79,0,136,0,5,0,155,0,10,0,0,0,192,0,0,0,0,0,157,0,97,0,0,0,74,0,131,0,26,0,14,0,4,0,71,0,221,0,8,0,170,0,244,0,117,0,114,0,103,0,0,0,0,0,0,0,199,0,22,0,89,0,230,0,246,0,167,0,14,0,252,0,73,0,108,0,0,0,0,0,0,0,155,0,92,0,201,0,20,0,113,0,0,0,0,0,171,0,0,0,37,0,249,0,13,0,109,0,98,0,187,0,0,0,19,0,184,0,136,0,101,0,174,0,174,0,3,0,136,0,0,0,71,0,99,0,108,0,67,0,109,0,60,0,162,0,192,0,221,0,113,0,192,0,7,0,219,0,67,0,229,0,100,0,236,0,0,0,0,0,177,0,184,0,214,0,13,0,79,0,0,0,0,0,0,0,31,0,13,0,141,0,25,0,111,0,13,0,10,0,193,0,78,0,57,0,198,0,66,0,23,0,136,0,73,0,0,0,195,0,72,0,165,0,251,0,187,0,111,0,16,0,235,0,0,0,245,0,109,0,12,0,253,0,43,0,219,0,31,0,98,0,17,0,175,0,191,0,176,0,230,0,53,0,202,0,125,0,183,0,74,0,24,0,86,0,173,0,149,0,201,0,36,0,70,0,0,0,14,0,0,0,177,0,41,0,0,0,0,0,10,0,0,0,144,0,108,0,204,0,16,0,0,0,229,0,206,0,245,0,176,0,12,0,46,0,52,0,58,0,175,0,69,0,105,0,241,0,62,0,102,0,189,0,73,0,111,0,134,0,122,0,0,0,115,0,205,0,242,0,137,0,246,0,0,0,87,0,30,0,109,0,3,0,0,0,155,0,80,0,0,0,25,0,0,0,121,0,95,0,235,0,0,0,209,0,0,0,24,0,148,0,208,0,153,0,194,0,136,0,249,0,157,0,253,0,104,0,71,0,206,0,119,0,94,0,244,0,1,0,236,0,88,0,126,0,21,0,0,0,109,0,155,0,0,0,0,0,103,0,161,0,0,0,26,0,76,0,115,0,225,0,48,0,107,0,228,0,0,0,0,0,0,0,77,0,194,0,165,0,9,0,0,0,13,0,55,0,241,0,224,0,251,0,169,0,0,0,0,0,0,0,42,0,0,0,65,0,63,0,9,0,128,0,10,0,68,0,0,0,0,0,0,0,27,0,0,0,241,0,2,0,143,0,0,0,117,0,127,0,43,0,220,0,244,0,95,0,142,0,84,0,81,0,139,0,0,0,169,0,159,0,91,0,0,0,0,0,165,0,147,0,216,0,73,0,0,0,58,0,52,0,0,0,0,0,0,0,40,0,164,0,69,0,163,0,0,0,0,0,73,0,166,0,155,0,206,0,14,0,11,0,177,0,89,0,0,0,252,0,179,0,220,0,6,0,155,0,142,0,0,0,0,0,0,0,0,0,194,0,180,0,0,0,7,0,46,0,149,0,49,0,144,0,3,0,249,0,182,0,2,0,60,0,212,0,115,0,68,0,199,0,216,0,252,0,184,0,226,0,66,0,135,0,96,0,0,0,156,0,46,0,39,0,0,0,243,0,0,0,249,0,26,0,126,0,45,0,156,0,249,0,117,0,221,0,0,0,93,0,47,0,48,0,0,0,29,0,160,0,0,0,96,0,221,0,237,0,149,0,198,0,247,0,66,0,234,0,101,0,192,0,74,0,0,0,173,0,19,0,103,0,144,0,17,0,168,0,147,0,58,0,0,0,213,0,204,0,245,0,24,0,247,0,223,0,156,0,144,0,0,0,229,0,225,0,176,0,229,0,170,0,30,0,230,0,218,0,30,0,183,0,15,0,236,0,197,0,69,0,196,0,112,0,0,0,0,0,60,0,127,0);
signal scenario_full  : scenario_type := (105,31,20,31,123,31,152,31,19,31,19,30,178,31,88,31,48,31,106,31,156,31,156,30,175,31,16,31,9,31,179,31,216,31,216,30,86,31,154,31,41,31,41,30,49,31,134,31,51,31,216,31,145,31,58,31,58,30,58,29,113,31,4,31,4,30,241,31,233,31,233,30,8,31,9,31,138,31,129,31,113,31,247,31,184,31,113,31,144,31,144,30,185,31,26,31,38,31,63,31,175,31,12,31,251,31,127,31,42,31,150,31,71,31,134,31,134,30,195,31,210,31,210,30,231,31,231,30,231,29,176,31,246,31,21,31,14,31,168,31,168,30,234,31,234,30,31,31,241,31,76,31,83,31,91,31,217,31,123,31,123,30,132,31,132,30,132,29,132,28,114,31,29,31,212,31,203,31,85,31,203,31,29,31,29,30,251,31,220,31,220,30,159,31,220,31,220,30,89,31,89,30,176,31,76,31,76,30,41,31,41,30,138,31,101,31,200,31,127,31,252,31,252,30,32,31,170,31,120,31,120,30,66,31,66,30,77,31,68,31,68,30,134,31,134,30,173,31,166,31,41,31,134,31,134,30,73,31,50,31,111,31,19,31,229,31,7,31,125,31,9,31,173,31,127,31,161,31,146,31,146,30,146,29,15,31,15,30,94,31,94,30,92,31,92,30,198,31,162,31,162,30,11,31,231,31,251,31,105,31,154,31,154,30,154,29,154,28,82,31,6,31,201,31,71,31,223,31,224,31,224,30,14,31,52,31,132,31,107,31,101,31,23,31,23,30,170,31,172,31,172,30,25,31,144,31,186,31,220,31,133,31,17,31,46,31,32,31,195,31,100,31,233,31,233,30,131,31,6,31,190,31,85,31,105,31,74,31,112,31,211,31,196,31,230,31,68,31,127,31,142,31,204,31,235,31,12,31,12,30,12,29,188,31,175,31,19,31,141,31,149,31,88,31,31,31,229,31,84,31,230,31,20,31,20,30,175,31,42,31,165,31,4,31,153,31,203,31,235,31,161,31,179,31,179,30,222,31,44,31,109,31,56,31,46,31,166,31,135,31,135,30,135,29,234,31,234,30,234,29,4,31,19,31,132,31,132,30,132,29,139,31,65,31,169,31,118,31,84,31,28,31,100,31,154,31,17,31,14,31,175,31,175,30,175,29,175,28,175,27,146,31,255,31,167,31,98,31,218,31,37,31,110,31,110,30,88,31,196,31,57,31,57,30,57,29,57,28,228,31,148,31,14,31,27,31,149,31,129,31,129,30,79,31,136,31,5,31,155,31,10,31,10,30,192,31,192,30,192,29,157,31,97,31,97,30,74,31,131,31,26,31,14,31,4,31,71,31,221,31,8,31,170,31,244,31,117,31,114,31,103,31,103,30,103,29,103,28,199,31,22,31,89,31,230,31,246,31,167,31,14,31,252,31,73,31,108,31,108,30,108,29,108,28,155,31,92,31,201,31,20,31,113,31,113,30,113,29,171,31,171,30,37,31,249,31,13,31,109,31,98,31,187,31,187,30,19,31,184,31,136,31,101,31,174,31,174,31,3,31,136,31,136,30,71,31,99,31,108,31,67,31,109,31,60,31,162,31,192,31,221,31,113,31,192,31,7,31,219,31,67,31,229,31,100,31,236,31,236,30,236,29,177,31,184,31,214,31,13,31,79,31,79,30,79,29,79,28,31,31,13,31,141,31,25,31,111,31,13,31,10,31,193,31,78,31,57,31,198,31,66,31,23,31,136,31,73,31,73,30,195,31,72,31,165,31,251,31,187,31,111,31,16,31,235,31,235,30,245,31,109,31,12,31,253,31,43,31,219,31,31,31,98,31,17,31,175,31,191,31,176,31,230,31,53,31,202,31,125,31,183,31,74,31,24,31,86,31,173,31,149,31,201,31,36,31,70,31,70,30,14,31,14,30,177,31,41,31,41,30,41,29,10,31,10,30,144,31,108,31,204,31,16,31,16,30,229,31,206,31,245,31,176,31,12,31,46,31,52,31,58,31,175,31,69,31,105,31,241,31,62,31,102,31,189,31,73,31,111,31,134,31,122,31,122,30,115,31,205,31,242,31,137,31,246,31,246,30,87,31,30,31,109,31,3,31,3,30,155,31,80,31,80,30,25,31,25,30,121,31,95,31,235,31,235,30,209,31,209,30,24,31,148,31,208,31,153,31,194,31,136,31,249,31,157,31,253,31,104,31,71,31,206,31,119,31,94,31,244,31,1,31,236,31,88,31,126,31,21,31,21,30,109,31,155,31,155,30,155,29,103,31,161,31,161,30,26,31,76,31,115,31,225,31,48,31,107,31,228,31,228,30,228,29,228,28,77,31,194,31,165,31,9,31,9,30,13,31,55,31,241,31,224,31,251,31,169,31,169,30,169,29,169,28,42,31,42,30,65,31,63,31,9,31,128,31,10,31,68,31,68,30,68,29,68,28,27,31,27,30,241,31,2,31,143,31,143,30,117,31,127,31,43,31,220,31,244,31,95,31,142,31,84,31,81,31,139,31,139,30,169,31,159,31,91,31,91,30,91,29,165,31,147,31,216,31,73,31,73,30,58,31,52,31,52,30,52,29,52,28,40,31,164,31,69,31,163,31,163,30,163,29,73,31,166,31,155,31,206,31,14,31,11,31,177,31,89,31,89,30,252,31,179,31,220,31,6,31,155,31,142,31,142,30,142,29,142,28,142,27,194,31,180,31,180,30,7,31,46,31,149,31,49,31,144,31,3,31,249,31,182,31,2,31,60,31,212,31,115,31,68,31,199,31,216,31,252,31,184,31,226,31,66,31,135,31,96,31,96,30,156,31,46,31,39,31,39,30,243,31,243,30,249,31,26,31,126,31,45,31,156,31,249,31,117,31,221,31,221,30,93,31,47,31,48,31,48,30,29,31,160,31,160,30,96,31,221,31,237,31,149,31,198,31,247,31,66,31,234,31,101,31,192,31,74,31,74,30,173,31,19,31,103,31,144,31,17,31,168,31,147,31,58,31,58,30,213,31,204,31,245,31,24,31,247,31,223,31,156,31,144,31,144,30,229,31,225,31,176,31,229,31,170,31,30,31,230,31,218,31,30,31,183,31,15,31,236,31,197,31,69,31,196,31,112,31,112,30,112,29,60,31,127,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
