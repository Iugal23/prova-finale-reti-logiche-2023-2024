-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_287 is
end project_tb_287;

architecture project_tb_arch_287 of project_tb_287 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 632;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,134,0,26,0,158,0,138,0,112,0,18,0,249,0,214,0,123,0,26,0,41,0,0,0,235,0,170,0,53,0,68,0,60,0,0,0,16,0,46,0,93,0,202,0,200,0,0,0,179,0,59,0,197,0,49,0,133,0,174,0,29,0,160,0,49,0,25,0,0,0,242,0,177,0,0,0,0,0,132,0,103,0,205,0,138,0,173,0,190,0,81,0,0,0,40,0,0,0,238,0,0,0,110,0,237,0,0,0,0,0,153,0,0,0,201,0,32,0,0,0,255,0,219,0,247,0,28,0,0,0,199,0,195,0,6,0,65,0,40,0,240,0,6,0,51,0,72,0,120,0,85,0,232,0,28,0,208,0,250,0,5,0,159,0,0,0,102,0,174,0,94,0,0,0,31,0,74,0,247,0,19,0,70,0,246,0,150,0,129,0,131,0,188,0,123,0,158,0,0,0,13,0,173,0,106,0,118,0,135,0,233,0,44,0,60,0,111,0,199,0,2,0,34,0,212,0,156,0,27,0,60,0,185,0,251,0,0,0,0,0,190,0,124,0,94,0,43,0,0,0,0,0,0,0,103,0,0,0,247,0,182,0,167,0,109,0,244,0,203,0,0,0,0,0,136,0,0,0,184,0,119,0,127,0,128,0,142,0,186,0,183,0,19,0,0,0,0,0,0,0,160,0,0,0,192,0,0,0,28,0,1,0,5,0,147,0,112,0,24,0,0,0,126,0,41,0,224,0,186,0,76,0,216,0,0,0,51,0,165,0,220,0,19,0,170,0,171,0,0,0,222,0,0,0,67,0,72,0,107,0,222,0,224,0,1,0,173,0,245,0,0,0,0,0,180,0,0,0,99,0,64,0,53,0,0,0,104,0,251,0,183,0,100,0,136,0,207,0,140,0,2,0,4,0,101,0,49,0,201,0,0,0,0,0,206,0,184,0,186,0,95,0,177,0,0,0,216,0,86,0,74,0,0,0,61,0,156,0,72,0,140,0,61,0,170,0,31,0,59,0,134,0,202,0,228,0,151,0,137,0,214,0,0,0,210,0,104,0,28,0,255,0,114,0,0,0,0,0,190,0,0,0,164,0,12,0,106,0,206,0,98,0,250,0,174,0,90,0,92,0,27,0,0,0,167,0,99,0,29,0,40,0,0,0,103,0,109,0,252,0,50,0,71,0,23,0,0,0,208,0,74,0,0,0,0,0,0,0,226,0,90,0,102,0,20,0,30,0,0,0,251,0,42,0,252,0,18,0,192,0,219,0,198,0,0,0,250,0,208,0,253,0,106,0,38,0,186,0,104,0,249,0,8,0,132,0,24,0,0,0,204,0,197,0,15,0,111,0,236,0,132,0,0,0,249,0,103,0,82,0,2,0,40,0,0,0,84,0,205,0,179,0,183,0,0,0,229,0,219,0,23,0,248,0,0,0,100,0,230,0,153,0,0,0,151,0,145,0,192,0,70,0,33,0,141,0,78,0,0,0,66,0,0,0,187,0,120,0,65,0,234,0,213,0,139,0,200,0,38,0,0,0,165,0,137,0,22,0,0,0,245,0,16,0,38,0,240,0,255,0,162,0,0,0,76,0,0,0,71,0,248,0,0,0,148,0,196,0,0,0,76,0,252,0,16,0,0,0,91,0,51,0,200,0,77,0,177,0,4,0,117,0,85,0,240,0,0,0,99,0,248,0,0,0,123,0,184,0,176,0,56,0,28,0,199,0,20,0,20,0,90,0,35,0,30,0,0,0,202,0,0,0,147,0,97,0,27,0,254,0,86,0,0,0,0,0,0,0,92,0,81,0,27,0,216,0,68,0,189,0,217,0,171,0,182,0,0,0,170,0,0,0,0,0,150,0,111,0,0,0,183,0,177,0,234,0,0,0,100,0,106,0,88,0,74,0,183,0,68,0,245,0,24,0,154,0,223,0,60,0,0,0,114,0,183,0,76,0,208,0,117,0,0,0,74,0,0,0,223,0,0,0,53,0,155,0,125,0,223,0,71,0,39,0,0,0,4,0,105,0,89,0,98,0,0,0,0,0,0,0,123,0,206,0,48,0,221,0,0,0,15,0,123,0,139,0,167,0,123,0,22,0,130,0,60,0,0,0,16,0,189,0,14,0,250,0,58,0,249,0,194,0,50,0,0,0,0,0,72,0,136,0,18,0,24,0,142,0,100,0,0,0,0,0,130,0,111,0,8,0,28,0,52,0,202,0,248,0,0,0,0,0,0,0,230,0,0,0,83,0,171,0,0,0,10,0,182,0,167,0,119,0,136,0,15,0,169,0,134,0,176,0,50,0,144,0,103,0,160,0,6,0,170,0,82,0,214,0,0,0,224,0,0,0,229,0,190,0,253,0,225,0,19,0,38,0,18,0,83,0,221,0,3,0,80,0,70,0,88,0,239,0,86,0,160,0,154,0,231,0,0,0,172,0,143,0,147,0,233,0,59,0,64,0,206,0,112,0,30,0,207,0,0,0,239,0,178,0,239,0,170,0,28,0,198,0,47,0,10,0,254,0,0,0,0,0,0,0,230,0,14,0,51,0,0,0,0,0,21,0,0,0,36,0,11,0,145,0,137,0,122,0,0,0,0,0,78,0,135,0,0,0,0,0,70,0,48,0,38,0,124,0,151,0,196,0,225,0,16,0,24,0,91,0,126,0,116,0,8,0,178,0,167,0,0,0,0,0,201,0,66,0,187,0,18,0,213,0,0,0,0,0,67,0,123,0,240,0,0,0,49,0,194,0,89,0,237,0,0,0,0,0,89,0,138,0,150,0,87,0,9,0,78,0,17,0,184,0,213,0,63,0,5,0,97,0,191,0,232,0,2,0);
signal scenario_full  : scenario_type := (0,0,134,31,26,31,158,31,138,31,112,31,18,31,249,31,214,31,123,31,26,31,41,31,41,30,235,31,170,31,53,31,68,31,60,31,60,30,16,31,46,31,93,31,202,31,200,31,200,30,179,31,59,31,197,31,49,31,133,31,174,31,29,31,160,31,49,31,25,31,25,30,242,31,177,31,177,30,177,29,132,31,103,31,205,31,138,31,173,31,190,31,81,31,81,30,40,31,40,30,238,31,238,30,110,31,237,31,237,30,237,29,153,31,153,30,201,31,32,31,32,30,255,31,219,31,247,31,28,31,28,30,199,31,195,31,6,31,65,31,40,31,240,31,6,31,51,31,72,31,120,31,85,31,232,31,28,31,208,31,250,31,5,31,159,31,159,30,102,31,174,31,94,31,94,30,31,31,74,31,247,31,19,31,70,31,246,31,150,31,129,31,131,31,188,31,123,31,158,31,158,30,13,31,173,31,106,31,118,31,135,31,233,31,44,31,60,31,111,31,199,31,2,31,34,31,212,31,156,31,27,31,60,31,185,31,251,31,251,30,251,29,190,31,124,31,94,31,43,31,43,30,43,29,43,28,103,31,103,30,247,31,182,31,167,31,109,31,244,31,203,31,203,30,203,29,136,31,136,30,184,31,119,31,127,31,128,31,142,31,186,31,183,31,19,31,19,30,19,29,19,28,160,31,160,30,192,31,192,30,28,31,1,31,5,31,147,31,112,31,24,31,24,30,126,31,41,31,224,31,186,31,76,31,216,31,216,30,51,31,165,31,220,31,19,31,170,31,171,31,171,30,222,31,222,30,67,31,72,31,107,31,222,31,224,31,1,31,173,31,245,31,245,30,245,29,180,31,180,30,99,31,64,31,53,31,53,30,104,31,251,31,183,31,100,31,136,31,207,31,140,31,2,31,4,31,101,31,49,31,201,31,201,30,201,29,206,31,184,31,186,31,95,31,177,31,177,30,216,31,86,31,74,31,74,30,61,31,156,31,72,31,140,31,61,31,170,31,31,31,59,31,134,31,202,31,228,31,151,31,137,31,214,31,214,30,210,31,104,31,28,31,255,31,114,31,114,30,114,29,190,31,190,30,164,31,12,31,106,31,206,31,98,31,250,31,174,31,90,31,92,31,27,31,27,30,167,31,99,31,29,31,40,31,40,30,103,31,109,31,252,31,50,31,71,31,23,31,23,30,208,31,74,31,74,30,74,29,74,28,226,31,90,31,102,31,20,31,30,31,30,30,251,31,42,31,252,31,18,31,192,31,219,31,198,31,198,30,250,31,208,31,253,31,106,31,38,31,186,31,104,31,249,31,8,31,132,31,24,31,24,30,204,31,197,31,15,31,111,31,236,31,132,31,132,30,249,31,103,31,82,31,2,31,40,31,40,30,84,31,205,31,179,31,183,31,183,30,229,31,219,31,23,31,248,31,248,30,100,31,230,31,153,31,153,30,151,31,145,31,192,31,70,31,33,31,141,31,78,31,78,30,66,31,66,30,187,31,120,31,65,31,234,31,213,31,139,31,200,31,38,31,38,30,165,31,137,31,22,31,22,30,245,31,16,31,38,31,240,31,255,31,162,31,162,30,76,31,76,30,71,31,248,31,248,30,148,31,196,31,196,30,76,31,252,31,16,31,16,30,91,31,51,31,200,31,77,31,177,31,4,31,117,31,85,31,240,31,240,30,99,31,248,31,248,30,123,31,184,31,176,31,56,31,28,31,199,31,20,31,20,31,90,31,35,31,30,31,30,30,202,31,202,30,147,31,97,31,27,31,254,31,86,31,86,30,86,29,86,28,92,31,81,31,27,31,216,31,68,31,189,31,217,31,171,31,182,31,182,30,170,31,170,30,170,29,150,31,111,31,111,30,183,31,177,31,234,31,234,30,100,31,106,31,88,31,74,31,183,31,68,31,245,31,24,31,154,31,223,31,60,31,60,30,114,31,183,31,76,31,208,31,117,31,117,30,74,31,74,30,223,31,223,30,53,31,155,31,125,31,223,31,71,31,39,31,39,30,4,31,105,31,89,31,98,31,98,30,98,29,98,28,123,31,206,31,48,31,221,31,221,30,15,31,123,31,139,31,167,31,123,31,22,31,130,31,60,31,60,30,16,31,189,31,14,31,250,31,58,31,249,31,194,31,50,31,50,30,50,29,72,31,136,31,18,31,24,31,142,31,100,31,100,30,100,29,130,31,111,31,8,31,28,31,52,31,202,31,248,31,248,30,248,29,248,28,230,31,230,30,83,31,171,31,171,30,10,31,182,31,167,31,119,31,136,31,15,31,169,31,134,31,176,31,50,31,144,31,103,31,160,31,6,31,170,31,82,31,214,31,214,30,224,31,224,30,229,31,190,31,253,31,225,31,19,31,38,31,18,31,83,31,221,31,3,31,80,31,70,31,88,31,239,31,86,31,160,31,154,31,231,31,231,30,172,31,143,31,147,31,233,31,59,31,64,31,206,31,112,31,30,31,207,31,207,30,239,31,178,31,239,31,170,31,28,31,198,31,47,31,10,31,254,31,254,30,254,29,254,28,230,31,14,31,51,31,51,30,51,29,21,31,21,30,36,31,11,31,145,31,137,31,122,31,122,30,122,29,78,31,135,31,135,30,135,29,70,31,48,31,38,31,124,31,151,31,196,31,225,31,16,31,24,31,91,31,126,31,116,31,8,31,178,31,167,31,167,30,167,29,201,31,66,31,187,31,18,31,213,31,213,30,213,29,67,31,123,31,240,31,240,30,49,31,194,31,89,31,237,31,237,30,237,29,89,31,138,31,150,31,87,31,9,31,78,31,17,31,184,31,213,31,63,31,5,31,97,31,191,31,232,31,2,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
