-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 568;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (220,0,193,0,131,0,1,0,200,0,170,0,108,0,219,0,209,0,9,0,0,0,0,0,0,0,40,0,75,0,0,0,166,0,74,0,95,0,171,0,247,0,157,0,231,0,142,0,252,0,0,0,41,0,137,0,104,0,146,0,187,0,153,0,140,0,230,0,120,0,250,0,0,0,102,0,0,0,148,0,123,0,71,0,0,0,190,0,198,0,0,0,0,0,105,0,11,0,141,0,137,0,169,0,216,0,90,0,210,0,174,0,206,0,27,0,210,0,85,0,225,0,126,0,31,0,195,0,185,0,213,0,136,0,57,0,168,0,10,0,51,0,0,0,152,0,0,0,168,0,0,0,39,0,0,0,14,0,127,0,42,0,185,0,0,0,153,0,226,0,62,0,157,0,111,0,0,0,5,0,238,0,194,0,21,0,220,0,81,0,199,0,47,0,168,0,141,0,23,0,0,0,125,0,205,0,127,0,138,0,31,0,0,0,112,0,0,0,159,0,0,0,0,0,245,0,0,0,70,0,94,0,148,0,0,0,217,0,0,0,132,0,0,0,0,0,251,0,230,0,0,0,63,0,206,0,213,0,118,0,246,0,10,0,174,0,211,0,71,0,252,0,105,0,0,0,178,0,0,0,0,0,52,0,207,0,195,0,156,0,101,0,167,0,200,0,20,0,0,0,77,0,103,0,0,0,47,0,0,0,200,0,1,0,6,0,243,0,102,0,45,0,60,0,185,0,245,0,0,0,42,0,79,0,173,0,0,0,184,0,0,0,24,0,157,0,113,0,189,0,252,0,115,0,139,0,245,0,3,0,64,0,35,0,0,0,12,0,25,0,87,0,127,0,2,0,64,0,162,0,121,0,0,0,0,0,196,0,0,0,219,0,228,0,165,0,119,0,248,0,160,0,74,0,0,0,0,0,0,0,9,0,3,0,205,0,17,0,0,0,251,0,112,0,14,0,106,0,154,0,181,0,95,0,128,0,122,0,173,0,179,0,35,0,21,0,238,0,31,0,202,0,0,0,0,0,96,0,238,0,142,0,9,0,128,0,155,0,162,0,197,0,4,0,92,0,195,0,156,0,183,0,0,0,217,0,42,0,0,0,36,0,72,0,203,0,0,0,79,0,198,0,201,0,0,0,117,0,0,0,0,0,48,0,0,0,1,0,113,0,1,0,169,0,0,0,208,0,6,0,0,0,99,0,52,0,0,0,249,0,250,0,63,0,156,0,33,0,197,0,48,0,226,0,228,0,34,0,125,0,76,0,84,0,0,0,109,0,0,0,194,0,0,0,4,0,0,0,57,0,183,0,234,0,224,0,183,0,104,0,10,0,104,0,100,0,0,0,0,0,0,0,0,0,0,0,114,0,202,0,184,0,18,0,212,0,55,0,61,0,54,0,0,0,0,0,191,0,0,0,234,0,77,0,197,0,0,0,31,0,0,0,75,0,173,0,27,0,0,0,158,0,98,0,0,0,7,0,55,0,199,0,168,0,0,0,141,0,0,0,242,0,221,0,149,0,94,0,74,0,173,0,0,0,0,0,148,0,204,0,27,0,42,0,183,0,176,0,72,0,107,0,151,0,0,0,0,0,97,0,68,0,94,0,219,0,18,0,195,0,39,0,193,0,214,0,142,0,19,0,0,0,185,0,16,0,243,0,183,0,243,0,22,0,63,0,0,0,0,0,7,0,36,0,221,0,117,0,0,0,74,0,191,0,0,0,79,0,232,0,183,0,86,0,84,0,90,0,244,0,42,0,0,0,58,0,19,0,252,0,122,0,244,0,0,0,70,0,187,0,0,0,127,0,209,0,19,0,0,0,73,0,109,0,0,0,0,0,9,0,194,0,10,0,33,0,210,0,103,0,120,0,240,0,187,0,182,0,168,0,78,0,23,0,56,0,48,0,251,0,237,0,21,0,26,0,30,0,197,0,161,0,75,0,0,0,30,0,57,0,126,0,0,0,17,0,140,0,0,0,92,0,49,0,165,0,187,0,210,0,139,0,0,0,164,0,105,0,123,0,109,0,0,0,6,0,134,0,250,0,93,0,0,0,0,0,230,0,132,0,156,0,188,0,76,0,229,0,69,0,155,0,135,0,0,0,80,0,175,0,85,0,7,0,244,0,199,0,210,0,180,0,50,0,14,0,26,0,41,0,0,0,171,0,180,0,0,0,205,0,55,0,0,0,0,0,198,0,0,0,4,0,247,0,0,0,8,0,26,0,158,0,222,0,199,0,137,0,185,0,241,0,0,0,187,0,0,0,97,0,13,0,211,0,30,0,0,0,91,0,58,0,121,0,0,0,42,0,19,0,0,0,137,0,164,0,124,0,0,0,143,0,223,0,2,0,190,0,252,0,24,0,0,0,17,0,11,0,77,0,29,0,131,0,213,0,249,0,0,0,59,0,12,0,0,0,85,0,55,0,0,0,29,0,76,0,243,0,230,0,135,0,87,0,0,0,79,0,32,0,0,0,170,0,202,0,184,0,192,0,177,0,19,0,0,0,0,0,83,0,68,0,250,0,0,0,185,0,232,0,0,0,182,0,142,0);
signal scenario_full  : scenario_type := (220,31,193,31,131,31,1,31,200,31,170,31,108,31,219,31,209,31,9,31,9,30,9,29,9,28,40,31,75,31,75,30,166,31,74,31,95,31,171,31,247,31,157,31,231,31,142,31,252,31,252,30,41,31,137,31,104,31,146,31,187,31,153,31,140,31,230,31,120,31,250,31,250,30,102,31,102,30,148,31,123,31,71,31,71,30,190,31,198,31,198,30,198,29,105,31,11,31,141,31,137,31,169,31,216,31,90,31,210,31,174,31,206,31,27,31,210,31,85,31,225,31,126,31,31,31,195,31,185,31,213,31,136,31,57,31,168,31,10,31,51,31,51,30,152,31,152,30,168,31,168,30,39,31,39,30,14,31,127,31,42,31,185,31,185,30,153,31,226,31,62,31,157,31,111,31,111,30,5,31,238,31,194,31,21,31,220,31,81,31,199,31,47,31,168,31,141,31,23,31,23,30,125,31,205,31,127,31,138,31,31,31,31,30,112,31,112,30,159,31,159,30,159,29,245,31,245,30,70,31,94,31,148,31,148,30,217,31,217,30,132,31,132,30,132,29,251,31,230,31,230,30,63,31,206,31,213,31,118,31,246,31,10,31,174,31,211,31,71,31,252,31,105,31,105,30,178,31,178,30,178,29,52,31,207,31,195,31,156,31,101,31,167,31,200,31,20,31,20,30,77,31,103,31,103,30,47,31,47,30,200,31,1,31,6,31,243,31,102,31,45,31,60,31,185,31,245,31,245,30,42,31,79,31,173,31,173,30,184,31,184,30,24,31,157,31,113,31,189,31,252,31,115,31,139,31,245,31,3,31,64,31,35,31,35,30,12,31,25,31,87,31,127,31,2,31,64,31,162,31,121,31,121,30,121,29,196,31,196,30,219,31,228,31,165,31,119,31,248,31,160,31,74,31,74,30,74,29,74,28,9,31,3,31,205,31,17,31,17,30,251,31,112,31,14,31,106,31,154,31,181,31,95,31,128,31,122,31,173,31,179,31,35,31,21,31,238,31,31,31,202,31,202,30,202,29,96,31,238,31,142,31,9,31,128,31,155,31,162,31,197,31,4,31,92,31,195,31,156,31,183,31,183,30,217,31,42,31,42,30,36,31,72,31,203,31,203,30,79,31,198,31,201,31,201,30,117,31,117,30,117,29,48,31,48,30,1,31,113,31,1,31,169,31,169,30,208,31,6,31,6,30,99,31,52,31,52,30,249,31,250,31,63,31,156,31,33,31,197,31,48,31,226,31,228,31,34,31,125,31,76,31,84,31,84,30,109,31,109,30,194,31,194,30,4,31,4,30,57,31,183,31,234,31,224,31,183,31,104,31,10,31,104,31,100,31,100,30,100,29,100,28,100,27,100,26,114,31,202,31,184,31,18,31,212,31,55,31,61,31,54,31,54,30,54,29,191,31,191,30,234,31,77,31,197,31,197,30,31,31,31,30,75,31,173,31,27,31,27,30,158,31,98,31,98,30,7,31,55,31,199,31,168,31,168,30,141,31,141,30,242,31,221,31,149,31,94,31,74,31,173,31,173,30,173,29,148,31,204,31,27,31,42,31,183,31,176,31,72,31,107,31,151,31,151,30,151,29,97,31,68,31,94,31,219,31,18,31,195,31,39,31,193,31,214,31,142,31,19,31,19,30,185,31,16,31,243,31,183,31,243,31,22,31,63,31,63,30,63,29,7,31,36,31,221,31,117,31,117,30,74,31,191,31,191,30,79,31,232,31,183,31,86,31,84,31,90,31,244,31,42,31,42,30,58,31,19,31,252,31,122,31,244,31,244,30,70,31,187,31,187,30,127,31,209,31,19,31,19,30,73,31,109,31,109,30,109,29,9,31,194,31,10,31,33,31,210,31,103,31,120,31,240,31,187,31,182,31,168,31,78,31,23,31,56,31,48,31,251,31,237,31,21,31,26,31,30,31,197,31,161,31,75,31,75,30,30,31,57,31,126,31,126,30,17,31,140,31,140,30,92,31,49,31,165,31,187,31,210,31,139,31,139,30,164,31,105,31,123,31,109,31,109,30,6,31,134,31,250,31,93,31,93,30,93,29,230,31,132,31,156,31,188,31,76,31,229,31,69,31,155,31,135,31,135,30,80,31,175,31,85,31,7,31,244,31,199,31,210,31,180,31,50,31,14,31,26,31,41,31,41,30,171,31,180,31,180,30,205,31,55,31,55,30,55,29,198,31,198,30,4,31,247,31,247,30,8,31,26,31,158,31,222,31,199,31,137,31,185,31,241,31,241,30,187,31,187,30,97,31,13,31,211,31,30,31,30,30,91,31,58,31,121,31,121,30,42,31,19,31,19,30,137,31,164,31,124,31,124,30,143,31,223,31,2,31,190,31,252,31,24,31,24,30,17,31,11,31,77,31,29,31,131,31,213,31,249,31,249,30,59,31,12,31,12,30,85,31,55,31,55,30,29,31,76,31,243,31,230,31,135,31,87,31,87,30,79,31,32,31,32,30,170,31,202,31,184,31,192,31,177,31,19,31,19,30,19,29,83,31,68,31,250,31,250,30,185,31,232,31,232,30,182,31,142,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
