-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 664;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (147,0,87,0,55,0,51,0,0,0,0,0,77,0,191,0,0,0,157,0,227,0,196,0,150,0,97,0,0,0,112,0,82,0,198,0,0,0,197,0,246,0,150,0,235,0,30,0,0,0,204,0,51,0,0,0,189,0,200,0,227,0,246,0,0,0,146,0,132,0,133,0,117,0,0,0,244,0,16,0,61,0,38,0,0,0,96,0,186,0,0,0,0,0,133,0,86,0,0,0,133,0,78,0,0,0,2,0,76,0,130,0,0,0,57,0,123,0,31,0,25,0,254,0,0,0,67,0,12,0,110,0,186,0,204,0,41,0,203,0,171,0,178,0,217,0,30,0,165,0,0,0,135,0,119,0,178,0,51,0,108,0,0,0,10,0,133,0,60,0,179,0,0,0,185,0,0,0,129,0,121,0,204,0,82,0,0,0,251,0,81,0,85,0,8,0,17,0,134,0,0,0,61,0,115,0,192,0,192,0,72,0,241,0,193,0,223,0,123,0,28,0,0,0,247,0,76,0,147,0,0,0,0,0,217,0,113,0,156,0,86,0,42,0,188,0,53,0,196,0,58,0,255,0,0,0,176,0,89,0,165,0,0,0,0,0,93,0,238,0,165,0,73,0,25,0,60,0,0,0,0,0,60,0,0,0,174,0,184,0,98,0,32,0,0,0,246,0,251,0,159,0,0,0,147,0,83,0,107,0,163,0,79,0,50,0,0,0,195,0,65,0,34,0,48,0,235,0,59,0,111,0,30,0,251,0,0,0,186,0,87,0,75,0,168,0,5,0,8,0,111,0,90,0,108,0,40,0,69,0,0,0,232,0,0,0,227,0,126,0,224,0,185,0,0,0,77,0,158,0,0,0,18,0,105,0,103,0,148,0,208,0,0,0,108,0,179,0,44,0,190,0,126,0,85,0,255,0,44,0,0,0,225,0,158,0,40,0,25,0,0,0,103,0,0,0,72,0,0,0,248,0,69,0,95,0,101,0,54,0,88,0,124,0,38,0,168,0,128,0,100,0,0,0,174,0,100,0,0,0,138,0,121,0,122,0,139,0,163,0,10,0,0,0,0,0,142,0,235,0,0,0,198,0,184,0,68,0,85,0,0,0,192,0,159,0,27,0,0,0,135,0,147,0,231,0,0,0,100,0,62,0,236,0,255,0,240,0,150,0,25,0,0,0,0,0,139,0,0,0,27,0,0,0,0,0,249,0,189,0,199,0,18,0,194,0,195,0,201,0,113,0,116,0,0,0,0,0,209,0,155,0,186,0,148,0,226,0,110,0,161,0,146,0,94,0,19,0,207,0,0,0,23,0,90,0,4,0,107,0,6,0,228,0,0,0,213,0,221,0,165,0,134,0,0,0,113,0,169,0,215,0,60,0,39,0,44,0,0,0,0,0,39,0,243,0,163,0,78,0,176,0,0,0,151,0,231,0,7,0,162,0,152,0,17,0,0,0,231,0,249,0,252,0,105,0,127,0,137,0,35,0,109,0,106,0,0,0,208,0,0,0,86,0,0,0,238,0,151,0,103,0,0,0,206,0,114,0,127,0,3,0,0,0,147,0,69,0,96,0,157,0,150,0,175,0,232,0,99,0,66,0,83,0,115,0,0,0,184,0,44,0,139,0,64,0,0,0,93,0,111,0,173,0,108,0,142,0,45,0,3,0,65,0,13,0,3,0,105,0,150,0,17,0,125,0,188,0,102,0,222,0,0,0,78,0,86,0,135,0,4,0,225,0,249,0,198,0,163,0,63,0,82,0,1,0,89,0,9,0,0,0,239,0,0,0,62,0,27,0,197,0,206,0,0,0,33,0,57,0,140,0,109,0,227,0,210,0,0,0,0,0,1,0,0,0,11,0,225,0,174,0,4,0,69,0,121,0,151,0,98,0,16,0,7,0,50,0,232,0,1,0,175,0,47,0,0,0,212,0,194,0,220,0,0,0,233,0,116,0,0,0,82,0,209,0,0,0,37,0,221,0,236,0,58,0,112,0,0,0,45,0,0,0,129,0,252,0,160,0,77,0,172,0,178,0,118,0,1,0,178,0,82,0,104,0,175,0,205,0,102,0,245,0,44,0,229,0,12,0,66,0,0,0,180,0,154,0,185,0,140,0,81,0,162,0,164,0,87,0,138,0,10,0,65,0,231,0,152,0,0,0,236,0,0,0,143,0,0,0,215,0,3,0,131,0,211,0,234,0,57,0,186,0,187,0,0,0,41,0,66,0,72,0,133,0,0,0,237,0,60,0,13,0,33,0,233,0,30,0,131,0,0,0,21,0,40,0,218,0,167,0,0,0,242,0,0,0,0,0,78,0,213,0,71,0,114,0,0,0,0,0,59,0,209,0,225,0,114,0,171,0,41,0,9,0,91,0,171,0,59,0,38,0,192,0,136,0,186,0,40,0,221,0,246,0,239,0,211,0,112,0,138,0,0,0,39,0,228,0,0,0,245,0,142,0,20,0,42,0,196,0,177,0,226,0,251,0,39,0,0,0,223,0,16,0,0,0,0,0,0,0,121,0,0,0,250,0,246,0,127,0,156,0,156,0,0,0,0,0,145,0,198,0,0,0,135,0,76,0,78,0,0,0,197,0,88,0,140,0,25,0,37,0,181,0,132,0,9,0,108,0,27,0,84,0,141,0,0,0,248,0,30,0,0,0,36,0,41,0,0,0,129,0,84,0,52,0,217,0,225,0,123,0,209,0,0,0,0,0,101,0,194,0,158,0,124,0,0,0,240,0,118,0,129,0,134,0,12,0,50,0,0,0,216,0,94,0,121,0,253,0,161,0,95,0,250,0,0,0,0,0,166,0,176,0,0,0,179,0,0,0,0,0,149,0,182,0,0,0,151,0,0,0,24,0,238,0,0,0,0,0,0,0,230,0,0,0,204,0,53,0,227,0,0,0,166,0,209,0,246,0,238,0,116,0,13,0,24,0,3,0,0,0,83,0,0,0,143,0,139,0,182,0,5,0,71,0);
signal scenario_full  : scenario_type := (147,31,87,31,55,31,51,31,51,30,51,29,77,31,191,31,191,30,157,31,227,31,196,31,150,31,97,31,97,30,112,31,82,31,198,31,198,30,197,31,246,31,150,31,235,31,30,31,30,30,204,31,51,31,51,30,189,31,200,31,227,31,246,31,246,30,146,31,132,31,133,31,117,31,117,30,244,31,16,31,61,31,38,31,38,30,96,31,186,31,186,30,186,29,133,31,86,31,86,30,133,31,78,31,78,30,2,31,76,31,130,31,130,30,57,31,123,31,31,31,25,31,254,31,254,30,67,31,12,31,110,31,186,31,204,31,41,31,203,31,171,31,178,31,217,31,30,31,165,31,165,30,135,31,119,31,178,31,51,31,108,31,108,30,10,31,133,31,60,31,179,31,179,30,185,31,185,30,129,31,121,31,204,31,82,31,82,30,251,31,81,31,85,31,8,31,17,31,134,31,134,30,61,31,115,31,192,31,192,31,72,31,241,31,193,31,223,31,123,31,28,31,28,30,247,31,76,31,147,31,147,30,147,29,217,31,113,31,156,31,86,31,42,31,188,31,53,31,196,31,58,31,255,31,255,30,176,31,89,31,165,31,165,30,165,29,93,31,238,31,165,31,73,31,25,31,60,31,60,30,60,29,60,31,60,30,174,31,184,31,98,31,32,31,32,30,246,31,251,31,159,31,159,30,147,31,83,31,107,31,163,31,79,31,50,31,50,30,195,31,65,31,34,31,48,31,235,31,59,31,111,31,30,31,251,31,251,30,186,31,87,31,75,31,168,31,5,31,8,31,111,31,90,31,108,31,40,31,69,31,69,30,232,31,232,30,227,31,126,31,224,31,185,31,185,30,77,31,158,31,158,30,18,31,105,31,103,31,148,31,208,31,208,30,108,31,179,31,44,31,190,31,126,31,85,31,255,31,44,31,44,30,225,31,158,31,40,31,25,31,25,30,103,31,103,30,72,31,72,30,248,31,69,31,95,31,101,31,54,31,88,31,124,31,38,31,168,31,128,31,100,31,100,30,174,31,100,31,100,30,138,31,121,31,122,31,139,31,163,31,10,31,10,30,10,29,142,31,235,31,235,30,198,31,184,31,68,31,85,31,85,30,192,31,159,31,27,31,27,30,135,31,147,31,231,31,231,30,100,31,62,31,236,31,255,31,240,31,150,31,25,31,25,30,25,29,139,31,139,30,27,31,27,30,27,29,249,31,189,31,199,31,18,31,194,31,195,31,201,31,113,31,116,31,116,30,116,29,209,31,155,31,186,31,148,31,226,31,110,31,161,31,146,31,94,31,19,31,207,31,207,30,23,31,90,31,4,31,107,31,6,31,228,31,228,30,213,31,221,31,165,31,134,31,134,30,113,31,169,31,215,31,60,31,39,31,44,31,44,30,44,29,39,31,243,31,163,31,78,31,176,31,176,30,151,31,231,31,7,31,162,31,152,31,17,31,17,30,231,31,249,31,252,31,105,31,127,31,137,31,35,31,109,31,106,31,106,30,208,31,208,30,86,31,86,30,238,31,151,31,103,31,103,30,206,31,114,31,127,31,3,31,3,30,147,31,69,31,96,31,157,31,150,31,175,31,232,31,99,31,66,31,83,31,115,31,115,30,184,31,44,31,139,31,64,31,64,30,93,31,111,31,173,31,108,31,142,31,45,31,3,31,65,31,13,31,3,31,105,31,150,31,17,31,125,31,188,31,102,31,222,31,222,30,78,31,86,31,135,31,4,31,225,31,249,31,198,31,163,31,63,31,82,31,1,31,89,31,9,31,9,30,239,31,239,30,62,31,27,31,197,31,206,31,206,30,33,31,57,31,140,31,109,31,227,31,210,31,210,30,210,29,1,31,1,30,11,31,225,31,174,31,4,31,69,31,121,31,151,31,98,31,16,31,7,31,50,31,232,31,1,31,175,31,47,31,47,30,212,31,194,31,220,31,220,30,233,31,116,31,116,30,82,31,209,31,209,30,37,31,221,31,236,31,58,31,112,31,112,30,45,31,45,30,129,31,252,31,160,31,77,31,172,31,178,31,118,31,1,31,178,31,82,31,104,31,175,31,205,31,102,31,245,31,44,31,229,31,12,31,66,31,66,30,180,31,154,31,185,31,140,31,81,31,162,31,164,31,87,31,138,31,10,31,65,31,231,31,152,31,152,30,236,31,236,30,143,31,143,30,215,31,3,31,131,31,211,31,234,31,57,31,186,31,187,31,187,30,41,31,66,31,72,31,133,31,133,30,237,31,60,31,13,31,33,31,233,31,30,31,131,31,131,30,21,31,40,31,218,31,167,31,167,30,242,31,242,30,242,29,78,31,213,31,71,31,114,31,114,30,114,29,59,31,209,31,225,31,114,31,171,31,41,31,9,31,91,31,171,31,59,31,38,31,192,31,136,31,186,31,40,31,221,31,246,31,239,31,211,31,112,31,138,31,138,30,39,31,228,31,228,30,245,31,142,31,20,31,42,31,196,31,177,31,226,31,251,31,39,31,39,30,223,31,16,31,16,30,16,29,16,28,121,31,121,30,250,31,246,31,127,31,156,31,156,31,156,30,156,29,145,31,198,31,198,30,135,31,76,31,78,31,78,30,197,31,88,31,140,31,25,31,37,31,181,31,132,31,9,31,108,31,27,31,84,31,141,31,141,30,248,31,30,31,30,30,36,31,41,31,41,30,129,31,84,31,52,31,217,31,225,31,123,31,209,31,209,30,209,29,101,31,194,31,158,31,124,31,124,30,240,31,118,31,129,31,134,31,12,31,50,31,50,30,216,31,94,31,121,31,253,31,161,31,95,31,250,31,250,30,250,29,166,31,176,31,176,30,179,31,179,30,179,29,149,31,182,31,182,30,151,31,151,30,24,31,238,31,238,30,238,29,238,28,230,31,230,30,204,31,53,31,227,31,227,30,166,31,209,31,246,31,238,31,116,31,13,31,24,31,3,31,3,30,83,31,83,30,143,31,139,31,182,31,5,31,71,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
