-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_21 is
end project_tb_21;

architecture project_tb_arch_21 of project_tb_21 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 447;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (6,0,146,0,197,0,0,0,2,0,173,0,25,0,113,0,0,0,115,0,54,0,35,0,57,0,0,0,71,0,0,0,73,0,209,0,102,0,68,0,111,0,0,0,88,0,126,0,114,0,0,0,0,0,122,0,118,0,0,0,0,0,229,0,240,0,178,0,0,0,187,0,0,0,139,0,106,0,146,0,27,0,37,0,49,0,141,0,15,0,21,0,93,0,54,0,0,0,126,0,6,0,216,0,112,0,160,0,15,0,186,0,139,0,173,0,125,0,0,0,88,0,0,0,169,0,47,0,115,0,34,0,13,0,251,0,0,0,95,0,98,0,147,0,126,0,90,0,40,0,76,0,126,0,3,0,242,0,78,0,0,0,113,0,0,0,59,0,124,0,67,0,208,0,22,0,70,0,5,0,238,0,13,0,81,0,54,0,0,0,0,0,78,0,0,0,85,0,84,0,31,0,241,0,87,0,27,0,40,0,142,0,165,0,0,0,3,0,206,0,131,0,0,0,147,0,165,0,174,0,0,0,154,0,217,0,75,0,0,0,118,0,86,0,0,0,0,0,60,0,26,0,57,0,110,0,44,0,244,0,249,0,235,0,0,0,247,0,125,0,167,0,134,0,42,0,192,0,26,0,86,0,130,0,218,0,197,0,223,0,169,0,9,0,252,0,0,0,89,0,95,0,184,0,229,0,75,0,154,0,249,0,30,0,116,0,187,0,165,0,0,0,203,0,58,0,146,0,225,0,242,0,172,0,0,0,0,0,120,0,114,0,0,0,76,0,228,0,169,0,253,0,215,0,58,0,200,0,202,0,0,0,0,0,127,0,127,0,152,0,26,0,197,0,0,0,0,0,93,0,0,0,42,0,0,0,74,0,78,0,85,0,163,0,172,0,18,0,9,0,207,0,170,0,161,0,0,0,17,0,185,0,85,0,0,0,124,0,54,0,143,0,57,0,138,0,234,0,235,0,0,0,19,0,183,0,200,0,0,0,104,0,0,0,192,0,0,0,137,0,0,0,189,0,24,0,175,0,0,0,74,0,151,0,223,0,0,0,0,0,0,0,68,0,177,0,184,0,25,0,18,0,0,0,140,0,171,0,164,0,224,0,0,0,44,0,21,0,112,0,3,0,207,0,210,0,118,0,203,0,106,0,21,0,187,0,15,0,0,0,151,0,154,0,0,0,146,0,0,0,87,0,0,0,6,0,246,0,0,0,0,0,139,0,214,0,141,0,0,0,254,0,129,0,234,0,242,0,148,0,178,0,236,0,218,0,77,0,136,0,0,0,205,0,0,0,26,0,185,0,135,0,236,0,144,0,72,0,74,0,251,0,0,0,0,0,180,0,0,0,245,0,0,0,203,0,71,0,225,0,0,0,72,0,63,0,75,0,0,0,161,0,229,0,105,0,0,0,0,0,18,0,62,0,0,0,35,0,17,0,236,0,144,0,77,0,16,0,177,0,118,0,93,0,163,0,0,0,22,0,238,0,42,0,80,0,255,0,116,0,2,0,29,0,16,0,178,0,226,0,247,0,239,0,51,0,245,0,116,0,0,0,0,0,242,0,206,0,11,0,171,0,156,0,61,0,0,0,119,0,247,0,163,0,0,0,161,0,0,0,220,0,147,0,238,0,40,0,0,0,182,0,95,0,151,0,22,0,55,0,43,0,0,0,0,0,0,0,147,0,89,0,109,0,0,0,35,0,0,0,113,0,132,0,188,0,106,0,229,0,182,0,73,0,67,0,213,0,197,0,229,0,41,0,236,0,12,0,0,0,0,0,47,0,0,0,233,0,232,0,156,0,0,0,73,0,217,0,166,0,0,0,146,0,80,0,169,0,61,0,164,0,56,0,168,0,251,0,32,0,160,0,208,0,27,0,207,0,72,0,129,0,0,0,0,0,0,0,75,0,123,0,209,0,0,0,0,0,0,0,69,0,245,0,229,0,69,0,178,0,255,0,179,0,229,0,28,0,147,0,0,0,57,0,251,0,0,0,0,0,0,0,0,0);
signal scenario_full  : scenario_type := (6,31,146,31,197,31,197,30,2,31,173,31,25,31,113,31,113,30,115,31,54,31,35,31,57,31,57,30,71,31,71,30,73,31,209,31,102,31,68,31,111,31,111,30,88,31,126,31,114,31,114,30,114,29,122,31,118,31,118,30,118,29,229,31,240,31,178,31,178,30,187,31,187,30,139,31,106,31,146,31,27,31,37,31,49,31,141,31,15,31,21,31,93,31,54,31,54,30,126,31,6,31,216,31,112,31,160,31,15,31,186,31,139,31,173,31,125,31,125,30,88,31,88,30,169,31,47,31,115,31,34,31,13,31,251,31,251,30,95,31,98,31,147,31,126,31,90,31,40,31,76,31,126,31,3,31,242,31,78,31,78,30,113,31,113,30,59,31,124,31,67,31,208,31,22,31,70,31,5,31,238,31,13,31,81,31,54,31,54,30,54,29,78,31,78,30,85,31,84,31,31,31,241,31,87,31,27,31,40,31,142,31,165,31,165,30,3,31,206,31,131,31,131,30,147,31,165,31,174,31,174,30,154,31,217,31,75,31,75,30,118,31,86,31,86,30,86,29,60,31,26,31,57,31,110,31,44,31,244,31,249,31,235,31,235,30,247,31,125,31,167,31,134,31,42,31,192,31,26,31,86,31,130,31,218,31,197,31,223,31,169,31,9,31,252,31,252,30,89,31,95,31,184,31,229,31,75,31,154,31,249,31,30,31,116,31,187,31,165,31,165,30,203,31,58,31,146,31,225,31,242,31,172,31,172,30,172,29,120,31,114,31,114,30,76,31,228,31,169,31,253,31,215,31,58,31,200,31,202,31,202,30,202,29,127,31,127,31,152,31,26,31,197,31,197,30,197,29,93,31,93,30,42,31,42,30,74,31,78,31,85,31,163,31,172,31,18,31,9,31,207,31,170,31,161,31,161,30,17,31,185,31,85,31,85,30,124,31,54,31,143,31,57,31,138,31,234,31,235,31,235,30,19,31,183,31,200,31,200,30,104,31,104,30,192,31,192,30,137,31,137,30,189,31,24,31,175,31,175,30,74,31,151,31,223,31,223,30,223,29,223,28,68,31,177,31,184,31,25,31,18,31,18,30,140,31,171,31,164,31,224,31,224,30,44,31,21,31,112,31,3,31,207,31,210,31,118,31,203,31,106,31,21,31,187,31,15,31,15,30,151,31,154,31,154,30,146,31,146,30,87,31,87,30,6,31,246,31,246,30,246,29,139,31,214,31,141,31,141,30,254,31,129,31,234,31,242,31,148,31,178,31,236,31,218,31,77,31,136,31,136,30,205,31,205,30,26,31,185,31,135,31,236,31,144,31,72,31,74,31,251,31,251,30,251,29,180,31,180,30,245,31,245,30,203,31,71,31,225,31,225,30,72,31,63,31,75,31,75,30,161,31,229,31,105,31,105,30,105,29,18,31,62,31,62,30,35,31,17,31,236,31,144,31,77,31,16,31,177,31,118,31,93,31,163,31,163,30,22,31,238,31,42,31,80,31,255,31,116,31,2,31,29,31,16,31,178,31,226,31,247,31,239,31,51,31,245,31,116,31,116,30,116,29,242,31,206,31,11,31,171,31,156,31,61,31,61,30,119,31,247,31,163,31,163,30,161,31,161,30,220,31,147,31,238,31,40,31,40,30,182,31,95,31,151,31,22,31,55,31,43,31,43,30,43,29,43,28,147,31,89,31,109,31,109,30,35,31,35,30,113,31,132,31,188,31,106,31,229,31,182,31,73,31,67,31,213,31,197,31,229,31,41,31,236,31,12,31,12,30,12,29,47,31,47,30,233,31,232,31,156,31,156,30,73,31,217,31,166,31,166,30,146,31,80,31,169,31,61,31,164,31,56,31,168,31,251,31,32,31,160,31,208,31,27,31,207,31,72,31,129,31,129,30,129,29,129,28,75,31,123,31,209,31,209,30,209,29,209,28,69,31,245,31,229,31,69,31,178,31,255,31,179,31,229,31,28,31,147,31,147,30,57,31,251,31,251,30,251,29,251,28,251,27);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
