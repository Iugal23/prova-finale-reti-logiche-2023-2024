-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1021;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (212,0,0,0,172,0,51,0,0,0,99,0,21,0,0,0,219,0,254,0,184,0,217,0,158,0,24,0,3,0,98,0,244,0,247,0,0,0,110,0,54,0,0,0,0,0,74,0,171,0,184,0,140,0,73,0,137,0,143,0,62,0,243,0,80,0,126,0,95,0,87,0,86,0,0,0,32,0,10,0,0,0,74,0,0,0,192,0,37,0,187,0,169,0,0,0,143,0,126,0,18,0,145,0,156,0,210,0,196,0,0,0,198,0,96,0,170,0,15,0,2,0,155,0,145,0,130,0,0,0,0,0,0,0,171,0,180,0,148,0,39,0,129,0,88,0,4,0,43,0,0,0,81,0,22,0,70,0,165,0,100,0,16,0,68,0,191,0,218,0,124,0,3,0,0,0,0,0,61,0,238,0,49,0,103,0,108,0,0,0,0,0,103,0,140,0,246,0,130,0,126,0,43,0,64,0,0,0,0,0,95,0,153,0,243,0,0,0,0,0,32,0,63,0,89,0,76,0,150,0,169,0,157,0,3,0,0,0,107,0,233,0,229,0,145,0,199,0,248,0,113,0,184,0,51,0,189,0,0,0,109,0,202,0,27,0,0,0,106,0,201,0,19,0,71,0,167,0,99,0,162,0,0,0,0,0,0,0,140,0,11,0,164,0,70,0,150,0,35,0,100,0,0,0,61,0,0,0,0,0,216,0,2,0,90,0,145,0,238,0,136,0,159,0,22,0,0,0,242,0,162,0,34,0,137,0,102,0,228,0,67,0,0,0,215,0,68,0,253,0,0,0,213,0,4,0,123,0,16,0,104,0,10,0,106,0,164,0,0,0,243,0,116,0,0,0,159,0,45,0,0,0,71,0,205,0,34,0,121,0,29,0,0,0,168,0,51,0,0,0,245,0,163,0,72,0,195,0,0,0,0,0,13,0,172,0,121,0,0,0,11,0,108,0,137,0,68,0,153,0,0,0,189,0,250,0,222,0,0,0,0,0,181,0,135,0,57,0,0,0,145,0,0,0,71,0,0,0,153,0,28,0,125,0,0,0,247,0,46,0,210,0,0,0,236,0,138,0,177,0,127,0,177,0,236,0,0,0,7,0,85,0,1,0,0,0,125,0,38,0,24,0,185,0,172,0,0,0,158,0,209,0,128,0,36,0,0,0,217,0,185,0,150,0,58,0,17,0,211,0,164,0,165,0,0,0,75,0,134,0,5,0,169,0,0,0,138,0,203,0,101,0,246,0,244,0,0,0,157,0,153,0,180,0,0,0,0,0,255,0,241,0,227,0,39,0,0,0,67,0,61,0,158,0,0,0,114,0,31,0,0,0,223,0,194,0,247,0,231,0,107,0,131,0,151,0,21,0,152,0,0,0,16,0,0,0,90,0,102,0,133,0,0,0,0,0,231,0,0,0,216,0,59,0,0,0,108,0,0,0,167,0,216,0,34,0,75,0,255,0,241,0,0,0,45,0,198,0,204,0,206,0,0,0,44,0,140,0,139,0,94,0,166,0,0,0,130,0,48,0,88,0,116,0,72,0,246,0,223,0,158,0,213,0,223,0,250,0,0,0,74,0,225,0,225,0,0,0,169,0,0,0,0,0,154,0,0,0,109,0,149,0,0,0,116,0,119,0,241,0,0,0,249,0,151,0,11,0,134,0,59,0,161,0,226,0,178,0,118,0,60,0,0,0,134,0,48,0,52,0,0,0,0,0,128,0,58,0,22,0,106,0,0,0,55,0,165,0,65,0,216,0,251,0,121,0,138,0,88,0,159,0,104,0,67,0,61,0,201,0,9,0,0,0,54,0,35,0,100,0,26,0,148,0,127,0,0,0,119,0,27,0,131,0,121,0,8,0,0,0,80,0,203,0,27,0,152,0,90,0,106,0,165,0,142,0,128,0,221,0,65,0,67,0,190,0,0,0,0,0,165,0,0,0,164,0,27,0,159,0,149,0,141,0,153,0,0,0,0,0,233,0,79,0,29,0,3,0,234,0,114,0,159,0,0,0,14,0,234,0,0,0,165,0,12,0,213,0,0,0,244,0,66,0,241,0,8,0,183,0,0,0,40,0,10,0,0,0,197,0,195,0,249,0,202,0,77,0,217,0,40,0,68,0,36,0,173,0,78,0,193,0,20,0,157,0,0,0,33,0,201,0,121,0,129,0,201,0,0,0,174,0,55,0,0,0,0,0,0,0,147,0,240,0,0,0,237,0,0,0,0,0,3,0,0,0,68,0,243,0,18,0,208,0,253,0,160,0,55,0,0,0,103,0,246,0,167,0,0,0,179,0,137,0,0,0,239,0,157,0,64,0,215,0,23,0,7,0,228,0,223,0,28,0,117,0,0,0,96,0,228,0,199,0,154,0,20,0,197,0,38,0,206,0,15,0,13,0,112,0,213,0,12,0,240,0,46,0,107,0,215,0,208,0,142,0,85,0,26,0,60,0,0,0,151,0,0,0,59,0,71,0,222,0,75,0,208,0,202,0,152,0,33,0,248,0,93,0,128,0,181,0,232,0,177,0,84,0,212,0,0,0,199,0,104,0,130,0,122,0,120,0,19,0,86,0,230,0,0,0,232,0,0,0,10,0,166,0,137,0,0,0,20,0,244,0,199,0,225,0,86,0,186,0,0,0,166,0,146,0,170,0,61,0,245,0,0,0,61,0,179,0,38,0,253,0,127,0,30,0,223,0,161,0,171,0,12,0,187,0,16,0,144,0,178,0,32,0,171,0,136,0,130,0,24,0,65,0,0,0,3,0,221,0,190,0,195,0,107,0,25,0,0,0,193,0,111,0,80,0,99,0,0,0,140,0,25,0,252,0,95,0,59,0,139,0,161,0,92,0,9,0,212,0,96,0,62,0,0,0,125,0,0,0,38,0,89,0,79,0,101,0,220,0,0,0,53,0,88,0,71,0,186,0,101,0,142,0,213,0,0,0,130,0,36,0,59,0,41,0,0,0,184,0,173,0,0,0,8,0,153,0,0,0,165,0,8,0,178,0,0,0,0,0,145,0,39,0,0,0,33,0,127,0,152,0,177,0,92,0,132,0,60,0,74,0,47,0,189,0,0,0,39,0,92,0,128,0,0,0,93,0,0,0,53,0,69,0,213,0,0,0,143,0,187,0,0,0,0,0,0,0,128,0,120,0,199,0,166,0,0,0,117,0,95,0,0,0,161,0,58,0,58,0,0,0,191,0,46,0,155,0,0,0,142,0,166,0,113,0,204,0,106,0,45,0,197,0,203,0,127,0,94,0,149,0,0,0,255,0,0,0,143,0,107,0,6,0,160,0,102,0,198,0,80,0,119,0,0,0,97,0,8,0,57,0,106,0,174,0,0,0,147,0,0,0,68,0,159,0,0,0,185,0,193,0,153,0,133,0,47,0,144,0,11,0,72,0,0,0,88,0,22,0,95,0,15,0,0,0,0,0,86,0,24,0,16,0,19,0,7,0,60,0,0,0,38,0,0,0,73,0,241,0,53,0,170,0,98,0,0,0,112,0,0,0,60,0,49,0,40,0,158,0,29,0,22,0,113,0,0,0,52,0,167,0,221,0,154,0,218,0,0,0,120,0,0,0,45,0,0,0,78,0,230,0,211,0,135,0,172,0,129,0,157,0,185,0,211,0,118,0,0,0,60,0,253,0,202,0,93,0,83,0,190,0,19,0,50,0,100,0,0,0,0,0,202,0,0,0,250,0,0,0,250,0,129,0,108,0,193,0,109,0,160,0,12,0,31,0,0,0,47,0,234,0,0,0,103,0,182,0,0,0,0,0,87,0,181,0,187,0,58,0,239,0,0,0,129,0,173,0,172,0,5,0,70,0,217,0,0,0,104,0,71,0,77,0,56,0,0,0,195,0,255,0,0,0,0,0,226,0,198,0,0,0,241,0,0,0,111,0,26,0,31,0,64,0,181,0,77,0,55,0,0,0,0,0,19,0,57,0,102,0,166,0,126,0,255,0,165,0,0,0,234,0,130,0,57,0,50,0,42,0,120,0,0,0,157,0,0,0,147,0,209,0,192,0,36,0,0,0,0,0,35,0,46,0,248,0,113,0,72,0,85,0,0,0,238,0,92,0,122,0,106,0,6,0,53,0,187,0,53,0,17,0,0,0,152,0,20,0,0,0,87,0,173,0,0,0,81,0,0,0,4,0,227,0,251,0,0,0,101,0,195,0,253,0,193,0,25,0,75,0,61,0,30,0,142,0,215,0,157,0,85,0,56,0,25,0,93,0,159,0,173,0,0,0,0,0,145,0,173,0,143,0,109,0,35,0,124,0,109,0,165,0,31,0,100,0,10,0,28,0,216,0,216,0,103,0,61,0,54,0,0,0,0,0,0,0,153,0,0,0,12,0,54,0,68,0,226,0,0,0,0,0,82,0,225,0,26,0,65,0,135,0,237,0,140,0,163,0,4,0,170,0,98,0,145,0,104,0,69,0,208,0,161,0,0,0,99,0,183,0,221,0,0,0,196,0,74,0,98,0,96,0,0,0,0,0,170,0,116,0,152,0,125,0,0,0,221,0,36,0,161,0,166,0,0,0,162,0,151,0,96,0,228,0,221,0,17,0);
signal scenario_full  : scenario_type := (212,31,212,30,172,31,51,31,51,30,99,31,21,31,21,30,219,31,254,31,184,31,217,31,158,31,24,31,3,31,98,31,244,31,247,31,247,30,110,31,54,31,54,30,54,29,74,31,171,31,184,31,140,31,73,31,137,31,143,31,62,31,243,31,80,31,126,31,95,31,87,31,86,31,86,30,32,31,10,31,10,30,74,31,74,30,192,31,37,31,187,31,169,31,169,30,143,31,126,31,18,31,145,31,156,31,210,31,196,31,196,30,198,31,96,31,170,31,15,31,2,31,155,31,145,31,130,31,130,30,130,29,130,28,171,31,180,31,148,31,39,31,129,31,88,31,4,31,43,31,43,30,81,31,22,31,70,31,165,31,100,31,16,31,68,31,191,31,218,31,124,31,3,31,3,30,3,29,61,31,238,31,49,31,103,31,108,31,108,30,108,29,103,31,140,31,246,31,130,31,126,31,43,31,64,31,64,30,64,29,95,31,153,31,243,31,243,30,243,29,32,31,63,31,89,31,76,31,150,31,169,31,157,31,3,31,3,30,107,31,233,31,229,31,145,31,199,31,248,31,113,31,184,31,51,31,189,31,189,30,109,31,202,31,27,31,27,30,106,31,201,31,19,31,71,31,167,31,99,31,162,31,162,30,162,29,162,28,140,31,11,31,164,31,70,31,150,31,35,31,100,31,100,30,61,31,61,30,61,29,216,31,2,31,90,31,145,31,238,31,136,31,159,31,22,31,22,30,242,31,162,31,34,31,137,31,102,31,228,31,67,31,67,30,215,31,68,31,253,31,253,30,213,31,4,31,123,31,16,31,104,31,10,31,106,31,164,31,164,30,243,31,116,31,116,30,159,31,45,31,45,30,71,31,205,31,34,31,121,31,29,31,29,30,168,31,51,31,51,30,245,31,163,31,72,31,195,31,195,30,195,29,13,31,172,31,121,31,121,30,11,31,108,31,137,31,68,31,153,31,153,30,189,31,250,31,222,31,222,30,222,29,181,31,135,31,57,31,57,30,145,31,145,30,71,31,71,30,153,31,28,31,125,31,125,30,247,31,46,31,210,31,210,30,236,31,138,31,177,31,127,31,177,31,236,31,236,30,7,31,85,31,1,31,1,30,125,31,38,31,24,31,185,31,172,31,172,30,158,31,209,31,128,31,36,31,36,30,217,31,185,31,150,31,58,31,17,31,211,31,164,31,165,31,165,30,75,31,134,31,5,31,169,31,169,30,138,31,203,31,101,31,246,31,244,31,244,30,157,31,153,31,180,31,180,30,180,29,255,31,241,31,227,31,39,31,39,30,67,31,61,31,158,31,158,30,114,31,31,31,31,30,223,31,194,31,247,31,231,31,107,31,131,31,151,31,21,31,152,31,152,30,16,31,16,30,90,31,102,31,133,31,133,30,133,29,231,31,231,30,216,31,59,31,59,30,108,31,108,30,167,31,216,31,34,31,75,31,255,31,241,31,241,30,45,31,198,31,204,31,206,31,206,30,44,31,140,31,139,31,94,31,166,31,166,30,130,31,48,31,88,31,116,31,72,31,246,31,223,31,158,31,213,31,223,31,250,31,250,30,74,31,225,31,225,31,225,30,169,31,169,30,169,29,154,31,154,30,109,31,149,31,149,30,116,31,119,31,241,31,241,30,249,31,151,31,11,31,134,31,59,31,161,31,226,31,178,31,118,31,60,31,60,30,134,31,48,31,52,31,52,30,52,29,128,31,58,31,22,31,106,31,106,30,55,31,165,31,65,31,216,31,251,31,121,31,138,31,88,31,159,31,104,31,67,31,61,31,201,31,9,31,9,30,54,31,35,31,100,31,26,31,148,31,127,31,127,30,119,31,27,31,131,31,121,31,8,31,8,30,80,31,203,31,27,31,152,31,90,31,106,31,165,31,142,31,128,31,221,31,65,31,67,31,190,31,190,30,190,29,165,31,165,30,164,31,27,31,159,31,149,31,141,31,153,31,153,30,153,29,233,31,79,31,29,31,3,31,234,31,114,31,159,31,159,30,14,31,234,31,234,30,165,31,12,31,213,31,213,30,244,31,66,31,241,31,8,31,183,31,183,30,40,31,10,31,10,30,197,31,195,31,249,31,202,31,77,31,217,31,40,31,68,31,36,31,173,31,78,31,193,31,20,31,157,31,157,30,33,31,201,31,121,31,129,31,201,31,201,30,174,31,55,31,55,30,55,29,55,28,147,31,240,31,240,30,237,31,237,30,237,29,3,31,3,30,68,31,243,31,18,31,208,31,253,31,160,31,55,31,55,30,103,31,246,31,167,31,167,30,179,31,137,31,137,30,239,31,157,31,64,31,215,31,23,31,7,31,228,31,223,31,28,31,117,31,117,30,96,31,228,31,199,31,154,31,20,31,197,31,38,31,206,31,15,31,13,31,112,31,213,31,12,31,240,31,46,31,107,31,215,31,208,31,142,31,85,31,26,31,60,31,60,30,151,31,151,30,59,31,71,31,222,31,75,31,208,31,202,31,152,31,33,31,248,31,93,31,128,31,181,31,232,31,177,31,84,31,212,31,212,30,199,31,104,31,130,31,122,31,120,31,19,31,86,31,230,31,230,30,232,31,232,30,10,31,166,31,137,31,137,30,20,31,244,31,199,31,225,31,86,31,186,31,186,30,166,31,146,31,170,31,61,31,245,31,245,30,61,31,179,31,38,31,253,31,127,31,30,31,223,31,161,31,171,31,12,31,187,31,16,31,144,31,178,31,32,31,171,31,136,31,130,31,24,31,65,31,65,30,3,31,221,31,190,31,195,31,107,31,25,31,25,30,193,31,111,31,80,31,99,31,99,30,140,31,25,31,252,31,95,31,59,31,139,31,161,31,92,31,9,31,212,31,96,31,62,31,62,30,125,31,125,30,38,31,89,31,79,31,101,31,220,31,220,30,53,31,88,31,71,31,186,31,101,31,142,31,213,31,213,30,130,31,36,31,59,31,41,31,41,30,184,31,173,31,173,30,8,31,153,31,153,30,165,31,8,31,178,31,178,30,178,29,145,31,39,31,39,30,33,31,127,31,152,31,177,31,92,31,132,31,60,31,74,31,47,31,189,31,189,30,39,31,92,31,128,31,128,30,93,31,93,30,53,31,69,31,213,31,213,30,143,31,187,31,187,30,187,29,187,28,128,31,120,31,199,31,166,31,166,30,117,31,95,31,95,30,161,31,58,31,58,31,58,30,191,31,46,31,155,31,155,30,142,31,166,31,113,31,204,31,106,31,45,31,197,31,203,31,127,31,94,31,149,31,149,30,255,31,255,30,143,31,107,31,6,31,160,31,102,31,198,31,80,31,119,31,119,30,97,31,8,31,57,31,106,31,174,31,174,30,147,31,147,30,68,31,159,31,159,30,185,31,193,31,153,31,133,31,47,31,144,31,11,31,72,31,72,30,88,31,22,31,95,31,15,31,15,30,15,29,86,31,24,31,16,31,19,31,7,31,60,31,60,30,38,31,38,30,73,31,241,31,53,31,170,31,98,31,98,30,112,31,112,30,60,31,49,31,40,31,158,31,29,31,22,31,113,31,113,30,52,31,167,31,221,31,154,31,218,31,218,30,120,31,120,30,45,31,45,30,78,31,230,31,211,31,135,31,172,31,129,31,157,31,185,31,211,31,118,31,118,30,60,31,253,31,202,31,93,31,83,31,190,31,19,31,50,31,100,31,100,30,100,29,202,31,202,30,250,31,250,30,250,31,129,31,108,31,193,31,109,31,160,31,12,31,31,31,31,30,47,31,234,31,234,30,103,31,182,31,182,30,182,29,87,31,181,31,187,31,58,31,239,31,239,30,129,31,173,31,172,31,5,31,70,31,217,31,217,30,104,31,71,31,77,31,56,31,56,30,195,31,255,31,255,30,255,29,226,31,198,31,198,30,241,31,241,30,111,31,26,31,31,31,64,31,181,31,77,31,55,31,55,30,55,29,19,31,57,31,102,31,166,31,126,31,255,31,165,31,165,30,234,31,130,31,57,31,50,31,42,31,120,31,120,30,157,31,157,30,147,31,209,31,192,31,36,31,36,30,36,29,35,31,46,31,248,31,113,31,72,31,85,31,85,30,238,31,92,31,122,31,106,31,6,31,53,31,187,31,53,31,17,31,17,30,152,31,20,31,20,30,87,31,173,31,173,30,81,31,81,30,4,31,227,31,251,31,251,30,101,31,195,31,253,31,193,31,25,31,75,31,61,31,30,31,142,31,215,31,157,31,85,31,56,31,25,31,93,31,159,31,173,31,173,30,173,29,145,31,173,31,143,31,109,31,35,31,124,31,109,31,165,31,31,31,100,31,10,31,28,31,216,31,216,31,103,31,61,31,54,31,54,30,54,29,54,28,153,31,153,30,12,31,54,31,68,31,226,31,226,30,226,29,82,31,225,31,26,31,65,31,135,31,237,31,140,31,163,31,4,31,170,31,98,31,145,31,104,31,69,31,208,31,161,31,161,30,99,31,183,31,221,31,221,30,196,31,74,31,98,31,96,31,96,30,96,29,170,31,116,31,152,31,125,31,125,30,221,31,36,31,161,31,166,31,166,30,162,31,151,31,96,31,228,31,221,31,17,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
