-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_726 is
end project_tb_726;

architecture project_tb_arch_726 of project_tb_726 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 856;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (113,0,0,0,0,0,179,0,230,0,3,0,113,0,0,0,43,0,231,0,139,0,64,0,0,0,87,0,242,0,30,0,20,0,0,0,31,0,168,0,114,0,167,0,227,0,91,0,69,0,255,0,110,0,31,0,0,0,0,0,61,0,55,0,235,0,0,0,0,0,70,0,91,0,90,0,0,0,230,0,189,0,232,0,122,0,164,0,28,0,124,0,178,0,0,0,20,0,139,0,228,0,251,0,21,0,177,0,74,0,152,0,252,0,199,0,0,0,73,0,0,0,229,0,0,0,0,0,86,0,32,0,112,0,41,0,0,0,89,0,213,0,0,0,55,0,204,0,215,0,219,0,0,0,83,0,175,0,55,0,0,0,0,0,0,0,203,0,144,0,150,0,0,0,99,0,248,0,45,0,109,0,44,0,0,0,33,0,116,0,143,0,33,0,112,0,147,0,100,0,53,0,239,0,202,0,59,0,28,0,102,0,220,0,0,0,72,0,187,0,170,0,0,0,227,0,250,0,51,0,19,0,0,0,143,0,203,0,216,0,0,0,166,0,83,0,253,0,131,0,200,0,0,0,232,0,67,0,243,0,110,0,189,0,0,0,128,0,0,0,0,0,50,0,0,0,220,0,221,0,180,0,151,0,87,0,0,0,8,0,55,0,89,0,0,0,196,0,12,0,134,0,196,0,170,0,90,0,0,0,29,0,169,0,27,0,0,0,159,0,3,0,163,0,243,0,57,0,232,0,30,0,55,0,8,0,0,0,31,0,213,0,102,0,90,0,214,0,0,0,209,0,182,0,199,0,0,0,96,0,133,0,194,0,67,0,0,0,237,0,215,0,0,0,251,0,200,0,252,0,18,0,107,0,133,0,181,0,0,0,132,0,1,0,51,0,153,0,9,0,235,0,113,0,32,0,69,0,90,0,101,0,34,0,0,0,112,0,137,0,154,0,248,0,97,0,223,0,244,0,23,0,0,0,162,0,0,0,191,0,190,0,84,0,156,0,18,0,162,0,209,0,0,0,64,0,50,0,23,0,189,0,0,0,241,0,24,0,0,0,0,0,140,0,143,0,64,0,111,0,0,0,244,0,198,0,114,0,11,0,76,0,82,0,106,0,219,0,0,0,25,0,180,0,0,0,0,0,157,0,0,0,109,0,140,0,139,0,124,0,36,0,142,0,134,0,152,0,73,0,15,0,175,0,60,0,0,0,21,0,149,0,109,0,83,0,7,0,0,0,225,0,141,0,187,0,0,0,238,0,208,0,112,0,161,0,0,0,93,0,0,0,46,0,18,0,0,0,198,0,143,0,205,0,164,0,80,0,92,0,25,0,0,0,0,0,150,0,0,0,0,0,224,0,0,0,0,0,31,0,0,0,21,0,203,0,0,0,176,0,158,0,41,0,73,0,55,0,0,0,36,0,227,0,153,0,200,0,156,0,42,0,43,0,150,0,160,0,0,0,131,0,129,0,24,0,130,0,86,0,114,0,0,0,119,0,66,0,123,0,59,0,168,0,181,0,45,0,36,0,0,0,140,0,232,0,194,0,105,0,205,0,89,0,240,0,104,0,84,0,183,0,36,0,104,0,231,0,59,0,130,0,0,0,0,0,223,0,0,0,39,0,255,0,43,0,0,0,145,0,147,0,0,0,35,0,180,0,249,0,27,0,0,0,0,0,183,0,251,0,117,0,87,0,3,0,0,0,37,0,0,0,124,0,219,0,193,0,56,0,0,0,0,0,114,0,93,0,122,0,132,0,169,0,0,0,28,0,0,0,205,0,56,0,28,0,0,0,0,0,251,0,217,0,43,0,156,0,36,0,33,0,35,0,22,0,163,0,187,0,219,0,81,0,84,0,0,0,210,0,135,0,91,0,144,0,0,0,202,0,15,0,176,0,164,0,0,0,48,0,158,0,89,0,67,0,0,0,0,0,113,0,195,0,172,0,0,0,0,0,220,0,0,0,162,0,103,0,58,0,69,0,129,0,136,0,20,0,178,0,210,0,216,0,143,0,134,0,142,0,170,0,92,0,14,0,0,0,121,0,0,0,94,0,0,0,30,0,217,0,189,0,168,0,249,0,54,0,0,0,215,0,36,0,171,0,39,0,207,0,28,0,158,0,53,0,160,0,45,0,51,0,214,0,60,0,0,0,23,0,76,0,177,0,0,0,0,0,197,0,242,0,124,0,136,0,0,0,91,0,6,0,42,0,0,0,23,0,108,0,0,0,142,0,0,0,152,0,189,0,153,0,0,0,80,0,105,0,73,0,13,0,54,0,24,0,128,0,0,0,161,0,0,0,0,0,3,0,0,0,177,0,46,0,58,0,0,0,103,0,0,0,230,0,182,0,0,0,141,0,118,0,36,0,191,0,233,0,191,0,254,0,176,0,123,0,0,0,243,0,189,0,41,0,218,0,0,0,131,0,0,0,251,0,88,0,114,0,0,0,0,0,69,0,0,0,0,0,123,0,0,0,154,0,192,0,29,0,0,0,17,0,154,0,0,0,103,0,0,0,152,0,226,0,223,0,205,0,85,0,136,0,205,0,209,0,35,0,26,0,0,0,0,0,106,0,197,0,0,0,0,0,39,0,213,0,116,0,74,0,95,0,174,0,0,0,146,0,186,0,0,0,0,0,89,0,0,0,191,0,0,0,171,0,181,0,131,0,151,0,41,0,249,0,0,0,0,0,132,0,178,0,71,0,0,0,127,0,159,0,31,0,40,0,29,0,163,0,187,0,173,0,106,0,241,0,218,0,4,0,225,0,134,0,64,0,154,0,178,0,137,0,136,0,0,0,151,0,39,0,82,0,32,0,0,0,10,0,161,0,32,0,170,0,104,0,0,0,0,0,161,0,113,0,67,0,253,0,23,0,121,0,20,0,0,0,68,0,70,0,47,0,82,0,0,0,250,0,109,0,58,0,225,0,78,0,160,0,55,0,0,0,170,0,119,0,0,0,39,0,125,0,0,0,11,0,206,0,0,0,63,0,154,0,172,0,241,0,129,0,0,0,189,0,184,0,99,0,1,0,0,0,90,0,0,0,0,0,20,0,0,0,91,0,4,0,92,0,0,0,196,0,35,0,167,0,0,0,40,0,150,0,42,0,216,0,13,0,232,0,210,0,228,0,128,0,41,0,38,0,53,0,12,0,216,0,0,0,17,0,125,0,59,0,147,0,109,0,190,0,149,0,175,0,65,0,186,0,83,0,131,0,91,0,139,0,201,0,169,0,255,0,169,0,23,0,227,0,0,0,151,0,223,0,110,0,0,0,0,0,7,0,0,0,244,0,219,0,159,0,0,0,116,0,187,0,0,0,169,0,163,0,184,0,220,0,242,0,184,0,221,0,225,0,216,0,213,0,245,0,150,0,38,0,191,0,0,0,196,0,0,0,64,0,101,0,170,0,217,0,156,0,135,0,47,0,121,0,169,0,27,0,157,0,214,0,121,0,0,0,0,0,41,0,181,0,38,0,184,0,135,0,126,0,139,0,0,0,108,0,147,0,140,0,0,0,35,0,0,0,159,0,71,0,0,0,58,0,249,0,159,0,3,0,12,0,98,0,115,0,17,0,0,0,0,0,218,0,236,0,222,0,61,0,188,0,0,0,82,0,255,0,0,0,86,0,0,0,154,0,212,0,247,0,86,0,6,0,232,0,79,0,115,0,154,0,0,0,243,0,121,0,15,0,209,0,39,0,119,0,0,0,112,0,0,0,170,0,185,0,0,0,140,0,162,0,1,0,238,0,72,0,0,0,107,0,0,0,22,0,75,0,39,0,185,0,53,0,140,0,0,0,12,0,0,0,152,0,105,0,0,0,178,0,0,0,148,0,174,0,0,0);
signal scenario_full  : scenario_type := (113,31,113,30,113,29,179,31,230,31,3,31,113,31,113,30,43,31,231,31,139,31,64,31,64,30,87,31,242,31,30,31,20,31,20,30,31,31,168,31,114,31,167,31,227,31,91,31,69,31,255,31,110,31,31,31,31,30,31,29,61,31,55,31,235,31,235,30,235,29,70,31,91,31,90,31,90,30,230,31,189,31,232,31,122,31,164,31,28,31,124,31,178,31,178,30,20,31,139,31,228,31,251,31,21,31,177,31,74,31,152,31,252,31,199,31,199,30,73,31,73,30,229,31,229,30,229,29,86,31,32,31,112,31,41,31,41,30,89,31,213,31,213,30,55,31,204,31,215,31,219,31,219,30,83,31,175,31,55,31,55,30,55,29,55,28,203,31,144,31,150,31,150,30,99,31,248,31,45,31,109,31,44,31,44,30,33,31,116,31,143,31,33,31,112,31,147,31,100,31,53,31,239,31,202,31,59,31,28,31,102,31,220,31,220,30,72,31,187,31,170,31,170,30,227,31,250,31,51,31,19,31,19,30,143,31,203,31,216,31,216,30,166,31,83,31,253,31,131,31,200,31,200,30,232,31,67,31,243,31,110,31,189,31,189,30,128,31,128,30,128,29,50,31,50,30,220,31,221,31,180,31,151,31,87,31,87,30,8,31,55,31,89,31,89,30,196,31,12,31,134,31,196,31,170,31,90,31,90,30,29,31,169,31,27,31,27,30,159,31,3,31,163,31,243,31,57,31,232,31,30,31,55,31,8,31,8,30,31,31,213,31,102,31,90,31,214,31,214,30,209,31,182,31,199,31,199,30,96,31,133,31,194,31,67,31,67,30,237,31,215,31,215,30,251,31,200,31,252,31,18,31,107,31,133,31,181,31,181,30,132,31,1,31,51,31,153,31,9,31,235,31,113,31,32,31,69,31,90,31,101,31,34,31,34,30,112,31,137,31,154,31,248,31,97,31,223,31,244,31,23,31,23,30,162,31,162,30,191,31,190,31,84,31,156,31,18,31,162,31,209,31,209,30,64,31,50,31,23,31,189,31,189,30,241,31,24,31,24,30,24,29,140,31,143,31,64,31,111,31,111,30,244,31,198,31,114,31,11,31,76,31,82,31,106,31,219,31,219,30,25,31,180,31,180,30,180,29,157,31,157,30,109,31,140,31,139,31,124,31,36,31,142,31,134,31,152,31,73,31,15,31,175,31,60,31,60,30,21,31,149,31,109,31,83,31,7,31,7,30,225,31,141,31,187,31,187,30,238,31,208,31,112,31,161,31,161,30,93,31,93,30,46,31,18,31,18,30,198,31,143,31,205,31,164,31,80,31,92,31,25,31,25,30,25,29,150,31,150,30,150,29,224,31,224,30,224,29,31,31,31,30,21,31,203,31,203,30,176,31,158,31,41,31,73,31,55,31,55,30,36,31,227,31,153,31,200,31,156,31,42,31,43,31,150,31,160,31,160,30,131,31,129,31,24,31,130,31,86,31,114,31,114,30,119,31,66,31,123,31,59,31,168,31,181,31,45,31,36,31,36,30,140,31,232,31,194,31,105,31,205,31,89,31,240,31,104,31,84,31,183,31,36,31,104,31,231,31,59,31,130,31,130,30,130,29,223,31,223,30,39,31,255,31,43,31,43,30,145,31,147,31,147,30,35,31,180,31,249,31,27,31,27,30,27,29,183,31,251,31,117,31,87,31,3,31,3,30,37,31,37,30,124,31,219,31,193,31,56,31,56,30,56,29,114,31,93,31,122,31,132,31,169,31,169,30,28,31,28,30,205,31,56,31,28,31,28,30,28,29,251,31,217,31,43,31,156,31,36,31,33,31,35,31,22,31,163,31,187,31,219,31,81,31,84,31,84,30,210,31,135,31,91,31,144,31,144,30,202,31,15,31,176,31,164,31,164,30,48,31,158,31,89,31,67,31,67,30,67,29,113,31,195,31,172,31,172,30,172,29,220,31,220,30,162,31,103,31,58,31,69,31,129,31,136,31,20,31,178,31,210,31,216,31,143,31,134,31,142,31,170,31,92,31,14,31,14,30,121,31,121,30,94,31,94,30,30,31,217,31,189,31,168,31,249,31,54,31,54,30,215,31,36,31,171,31,39,31,207,31,28,31,158,31,53,31,160,31,45,31,51,31,214,31,60,31,60,30,23,31,76,31,177,31,177,30,177,29,197,31,242,31,124,31,136,31,136,30,91,31,6,31,42,31,42,30,23,31,108,31,108,30,142,31,142,30,152,31,189,31,153,31,153,30,80,31,105,31,73,31,13,31,54,31,24,31,128,31,128,30,161,31,161,30,161,29,3,31,3,30,177,31,46,31,58,31,58,30,103,31,103,30,230,31,182,31,182,30,141,31,118,31,36,31,191,31,233,31,191,31,254,31,176,31,123,31,123,30,243,31,189,31,41,31,218,31,218,30,131,31,131,30,251,31,88,31,114,31,114,30,114,29,69,31,69,30,69,29,123,31,123,30,154,31,192,31,29,31,29,30,17,31,154,31,154,30,103,31,103,30,152,31,226,31,223,31,205,31,85,31,136,31,205,31,209,31,35,31,26,31,26,30,26,29,106,31,197,31,197,30,197,29,39,31,213,31,116,31,74,31,95,31,174,31,174,30,146,31,186,31,186,30,186,29,89,31,89,30,191,31,191,30,171,31,181,31,131,31,151,31,41,31,249,31,249,30,249,29,132,31,178,31,71,31,71,30,127,31,159,31,31,31,40,31,29,31,163,31,187,31,173,31,106,31,241,31,218,31,4,31,225,31,134,31,64,31,154,31,178,31,137,31,136,31,136,30,151,31,39,31,82,31,32,31,32,30,10,31,161,31,32,31,170,31,104,31,104,30,104,29,161,31,113,31,67,31,253,31,23,31,121,31,20,31,20,30,68,31,70,31,47,31,82,31,82,30,250,31,109,31,58,31,225,31,78,31,160,31,55,31,55,30,170,31,119,31,119,30,39,31,125,31,125,30,11,31,206,31,206,30,63,31,154,31,172,31,241,31,129,31,129,30,189,31,184,31,99,31,1,31,1,30,90,31,90,30,90,29,20,31,20,30,91,31,4,31,92,31,92,30,196,31,35,31,167,31,167,30,40,31,150,31,42,31,216,31,13,31,232,31,210,31,228,31,128,31,41,31,38,31,53,31,12,31,216,31,216,30,17,31,125,31,59,31,147,31,109,31,190,31,149,31,175,31,65,31,186,31,83,31,131,31,91,31,139,31,201,31,169,31,255,31,169,31,23,31,227,31,227,30,151,31,223,31,110,31,110,30,110,29,7,31,7,30,244,31,219,31,159,31,159,30,116,31,187,31,187,30,169,31,163,31,184,31,220,31,242,31,184,31,221,31,225,31,216,31,213,31,245,31,150,31,38,31,191,31,191,30,196,31,196,30,64,31,101,31,170,31,217,31,156,31,135,31,47,31,121,31,169,31,27,31,157,31,214,31,121,31,121,30,121,29,41,31,181,31,38,31,184,31,135,31,126,31,139,31,139,30,108,31,147,31,140,31,140,30,35,31,35,30,159,31,71,31,71,30,58,31,249,31,159,31,3,31,12,31,98,31,115,31,17,31,17,30,17,29,218,31,236,31,222,31,61,31,188,31,188,30,82,31,255,31,255,30,86,31,86,30,154,31,212,31,247,31,86,31,6,31,232,31,79,31,115,31,154,31,154,30,243,31,121,31,15,31,209,31,39,31,119,31,119,30,112,31,112,30,170,31,185,31,185,30,140,31,162,31,1,31,238,31,72,31,72,30,107,31,107,30,22,31,75,31,39,31,185,31,53,31,140,31,140,30,12,31,12,30,152,31,105,31,105,30,178,31,178,30,148,31,174,31,174,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
