-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 216;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (94,0,89,0,0,0,139,0,119,0,131,0,210,0,62,0,232,0,88,0,76,0,216,0,183,0,160,0,41,0,51,0,0,0,125,0,217,0,47,0,236,0,243,0,249,0,0,0,47,0,184,0,116,0,130,0,121,0,173,0,164,0,243,0,56,0,144,0,136,0,19,0,0,0,117,0,0,0,0,0,0,0,0,0,18,0,204,0,0,0,50,0,211,0,39,0,85,0,88,0,58,0,127,0,0,0,0,0,67,0,132,0,234,0,68,0,0,0,4,0,158,0,104,0,0,0,9,0,105,0,150,0,109,0,131,0,186,0,58,0,94,0,67,0,0,0,0,0,240,0,113,0,155,0,148,0,0,0,232,0,108,0,39,0,0,0,129,0,27,0,180,0,201,0,118,0,0,0,0,0,24,0,224,0,156,0,0,0,143,0,0,0,0,0,83,0,163,0,36,0,5,0,122,0,0,0,160,0,160,0,0,0,0,0,113,0,142,0,44,0,254,0,198,0,205,0,98,0,90,0,108,0,235,0,194,0,76,0,87,0,246,0,214,0,158,0,175,0,137,0,23,0,0,0,0,0,85,0,162,0,54,0,0,0,106,0,0,0,41,0,113,0,0,0,122,0,123,0,32,0,0,0,0,0,171,0,20,0,170,0,0,0,67,0,63,0,111,0,37,0,147,0,119,0,0,0,0,0,90,0,247,0,228,0,98,0,171,0,12,0,0,0,108,0,245,0,249,0,167,0,255,0,13,0,10,0,225,0,21,0,134,0,142,0,175,0,194,0,17,0,131,0,54,0,31,0,169,0,203,0,107,0,194,0,204,0,99,0,74,0,54,0,166,0,140,0,60,0,0,0,191,0,40,0,255,0,50,0,94,0,168,0,219,0,61,0,150,0,31,0,170,0,177,0,157,0,72,0,64,0,56,0,33,0,226,0,193,0,140,0,172,0,0,0,124,0,0,0,255,0,118,0);
signal scenario_full  : scenario_type := (94,31,89,31,89,30,139,31,119,31,131,31,210,31,62,31,232,31,88,31,76,31,216,31,183,31,160,31,41,31,51,31,51,30,125,31,217,31,47,31,236,31,243,31,249,31,249,30,47,31,184,31,116,31,130,31,121,31,173,31,164,31,243,31,56,31,144,31,136,31,19,31,19,30,117,31,117,30,117,29,117,28,117,27,18,31,204,31,204,30,50,31,211,31,39,31,85,31,88,31,58,31,127,31,127,30,127,29,67,31,132,31,234,31,68,31,68,30,4,31,158,31,104,31,104,30,9,31,105,31,150,31,109,31,131,31,186,31,58,31,94,31,67,31,67,30,67,29,240,31,113,31,155,31,148,31,148,30,232,31,108,31,39,31,39,30,129,31,27,31,180,31,201,31,118,31,118,30,118,29,24,31,224,31,156,31,156,30,143,31,143,30,143,29,83,31,163,31,36,31,5,31,122,31,122,30,160,31,160,31,160,30,160,29,113,31,142,31,44,31,254,31,198,31,205,31,98,31,90,31,108,31,235,31,194,31,76,31,87,31,246,31,214,31,158,31,175,31,137,31,23,31,23,30,23,29,85,31,162,31,54,31,54,30,106,31,106,30,41,31,113,31,113,30,122,31,123,31,32,31,32,30,32,29,171,31,20,31,170,31,170,30,67,31,63,31,111,31,37,31,147,31,119,31,119,30,119,29,90,31,247,31,228,31,98,31,171,31,12,31,12,30,108,31,245,31,249,31,167,31,255,31,13,31,10,31,225,31,21,31,134,31,142,31,175,31,194,31,17,31,131,31,54,31,31,31,169,31,203,31,107,31,194,31,204,31,99,31,74,31,54,31,166,31,140,31,60,31,60,30,191,31,40,31,255,31,50,31,94,31,168,31,219,31,61,31,150,31,31,31,170,31,177,31,157,31,72,31,64,31,56,31,33,31,226,31,193,31,140,31,172,31,172,30,124,31,124,30,255,31,118,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
