-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 790;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (108,0,105,0,161,0,0,0,77,0,0,0,104,0,0,0,182,0,0,0,43,0,66,0,0,0,103,0,141,0,0,0,252,0,129,0,49,0,0,0,207,0,213,0,0,0,0,0,151,0,215,0,61,0,61,0,61,0,70,0,93,0,0,0,0,0,102,0,64,0,215,0,68,0,0,0,0,0,191,0,197,0,0,0,111,0,68,0,224,0,12,0,67,0,147,0,0,0,29,0,0,0,75,0,241,0,152,0,10,0,171,0,4,0,107,0,211,0,91,0,127,0,33,0,49,0,125,0,88,0,243,0,0,0,202,0,156,0,77,0,198,0,225,0,65,0,139,0,214,0,0,0,232,0,180,0,67,0,201,0,0,0,0,0,130,0,241,0,190,0,160,0,0,0,0,0,0,0,0,0,0,0,0,0,77,0,0,0,105,0,81,0,236,0,26,0,161,0,246,0,40,0,200,0,106,0,0,0,239,0,114,0,19,0,69,0,0,0,134,0,0,0,76,0,0,0,124,0,0,0,59,0,56,0,84,0,227,0,147,0,0,0,0,0,177,0,120,0,101,0,97,0,43,0,226,0,206,0,148,0,98,0,134,0,0,0,0,0,183,0,0,0,0,0,66,0,57,0,0,0,214,0,255,0,129,0,0,0,248,0,134,0,126,0,0,0,165,0,0,0,0,0,111,0,193,0,213,0,123,0,94,0,192,0,0,0,120,0,73,0,5,0,0,0,227,0,137,0,82,0,10,0,176,0,167,0,49,0,246,0,30,0,0,0,102,0,0,0,123,0,176,0,122,0,20,0,30,0,176,0,40,0,25,0,105,0,0,0,175,0,28,0,176,0,166,0,100,0,5,0,145,0,130,0,163,0,34,0,0,0,37,0,49,0,78,0,0,0,0,0,232,0,85,0,0,0,19,0,89,0,0,0,111,0,154,0,88,0,0,0,8,0,160,0,141,0,51,0,46,0,0,0,165,0,0,0,27,0,236,0,83,0,225,0,0,0,217,0,50,0,216,0,0,0,40,0,159,0,107,0,0,0,109,0,90,0,127,0,0,0,230,0,0,0,0,0,0,0,0,0,144,0,106,0,65,0,149,0,194,0,21,0,215,0,13,0,156,0,46,0,183,0,98,0,222,0,0,0,0,0,0,0,133,0,209,0,223,0,0,0,149,0,80,0,49,0,42,0,120,0,0,0,203,0,0,0,54,0,9,0,216,0,148,0,251,0,250,0,147,0,31,0,165,0,0,0,165,0,94,0,160,0,84,0,105,0,240,0,0,0,133,0,105,0,62,0,126,0,0,0,48,0,64,0,88,0,226,0,28,0,0,0,17,0,24,0,69,0,7,0,0,0,0,0,0,0,233,0,0,0,0,0,211,0,0,0,60,0,116,0,0,0,21,0,142,0,235,0,32,0,49,0,109,0,0,0,173,0,114,0,42,0,193,0,0,0,220,0,0,0,47,0,221,0,102,0,196,0,30,0,15,0,117,0,0,0,95,0,170,0,0,0,0,0,62,0,237,0,0,0,41,0,122,0,5,0,71,0,110,0,37,0,116,0,151,0,114,0,219,0,24,0,105,0,249,0,230,0,0,0,246,0,215,0,0,0,80,0,246,0,195,0,107,0,197,0,0,0,127,0,75,0,224,0,58,0,248,0,176,0,111,0,0,0,191,0,42,0,0,0,144,0,62,0,0,0,29,0,156,0,223,0,253,0,63,0,53,0,129,0,231,0,82,0,150,0,0,0,0,0,21,0,188,0,83,0,0,0,137,0,241,0,170,0,230,0,25,0,197,0,113,0,0,0,139,0,0,0,196,0,202,0,170,0,0,0,180,0,0,0,0,0,87,0,176,0,204,0,0,0,233,0,103,0,131,0,0,0,94,0,109,0,0,0,43,0,153,0,124,0,4,0,245,0,251,0,0,0,131,0,228,0,0,0,147,0,0,0,123,0,31,0,65,0,13,0,155,0,148,0,44,0,0,0,0,0,135,0,237,0,218,0,0,0,0,0,30,0,140,0,37,0,43,0,40,0,122,0,0,0,51,0,9,0,30,0,98,0,83,0,94,0,51,0,0,0,226,0,58,0,96,0,49,0,206,0,208,0,40,0,0,0,218,0,217,0,171,0,14,0,225,0,0,0,0,0,230,0,57,0,124,0,206,0,21,0,35,0,0,0,127,0,24,0,144,0,53,0,198,0,76,0,0,0,38,0,214,0,0,0,78,0,87,0,149,0,199,0,69,0,147,0,162,0,200,0,0,0,216,0,163,0,0,0,215,0,19,0,233,0,0,0,218,0,97,0,199,0,108,0,0,0,144,0,4,0,104,0,91,0,0,0,0,0,40,0,206,0,0,0,78,0,113,0,238,0,35,0,88,0,157,0,107,0,52,0,79,0,0,0,96,0,8,0,99,0,57,0,0,0,238,0,16,0,35,0,0,0,206,0,8,0,12,0,173,0,0,0,224,0,104,0,4,0,78,0,92,0,189,0,205,0,22,0,92,0,0,0,23,0,0,0,0,0,164,0,207,0,118,0,39,0,190,0,238,0,0,0,91,0,250,0,189,0,225,0,145,0,242,0,0,0,0,0,174,0,145,0,231,0,8,0,0,0,203,0,237,0,82,0,26,0,0,0,235,0,154,0,190,0,14,0,193,0,86,0,203,0,182,0,120,0,154,0,0,0,0,0,40,0,200,0,0,0,153,0,212,0,0,0,0,0,0,0,65,0,114,0,46,0,66,0,0,0,213,0,0,0,0,0,74,0,0,0,0,0,206,0,244,0,185,0,204,0,148,0,0,0,0,0,111,0,177,0,174,0,83,0,176,0,40,0,0,0,119,0,18,0,0,0,122,0,23,0,190,0,220,0,178,0,222,0,76,0,35,0,98,0,219,0,153,0,177,0,50,0,0,0,0,0,210,0,13,0,252,0,117,0,202,0,145,0,235,0,0,0,0,0,38,0,133,0,226,0,68,0,73,0,0,0,118,0,201,0,109,0,12,0,0,0,46,0,203,0,0,0,87,0,147,0,0,0,232,0,178,0,23,0,61,0,0,0,130,0,92,0,0,0,110,0,207,0,0,0,0,0,72,0,234,0,0,0,0,0,77,0,78,0,0,0,0,0,0,0,22,0,187,0,122,0,10,0,171,0,57,0,138,0,67,0,56,0,0,0,0,0,0,0,61,0,0,0,103,0,0,0,57,0,132,0,144,0,194,0,27,0,0,0,17,0,5,0,92,0,173,0,195,0,2,0,218,0,109,0,26,0,0,0,73,0,48,0,63,0,119,0,67,0,70,0,171,0,208,0,8,0,15,0,58,0,5,0,0,0,217,0,211,0,0,0,69,0,84,0,0,0,231,0,118,0,71,0,242,0,129,0,0,0,155,0,150,0,41,0,228,0,250,0,73,0,227,0,39,0,92,0,238,0,11,0,41,0,212,0,212,0,0,0,0,0,134,0,75,0,0,0,197,0,14,0,139,0,103,0,0,0,240,0,1,0,36,0,123,0,0,0,8,0,1,0,0,0,212,0,24,0,10,0,201,0);
signal scenario_full  : scenario_type := (108,31,105,31,161,31,161,30,77,31,77,30,104,31,104,30,182,31,182,30,43,31,66,31,66,30,103,31,141,31,141,30,252,31,129,31,49,31,49,30,207,31,213,31,213,30,213,29,151,31,215,31,61,31,61,31,61,31,70,31,93,31,93,30,93,29,102,31,64,31,215,31,68,31,68,30,68,29,191,31,197,31,197,30,111,31,68,31,224,31,12,31,67,31,147,31,147,30,29,31,29,30,75,31,241,31,152,31,10,31,171,31,4,31,107,31,211,31,91,31,127,31,33,31,49,31,125,31,88,31,243,31,243,30,202,31,156,31,77,31,198,31,225,31,65,31,139,31,214,31,214,30,232,31,180,31,67,31,201,31,201,30,201,29,130,31,241,31,190,31,160,31,160,30,160,29,160,28,160,27,160,26,160,25,77,31,77,30,105,31,81,31,236,31,26,31,161,31,246,31,40,31,200,31,106,31,106,30,239,31,114,31,19,31,69,31,69,30,134,31,134,30,76,31,76,30,124,31,124,30,59,31,56,31,84,31,227,31,147,31,147,30,147,29,177,31,120,31,101,31,97,31,43,31,226,31,206,31,148,31,98,31,134,31,134,30,134,29,183,31,183,30,183,29,66,31,57,31,57,30,214,31,255,31,129,31,129,30,248,31,134,31,126,31,126,30,165,31,165,30,165,29,111,31,193,31,213,31,123,31,94,31,192,31,192,30,120,31,73,31,5,31,5,30,227,31,137,31,82,31,10,31,176,31,167,31,49,31,246,31,30,31,30,30,102,31,102,30,123,31,176,31,122,31,20,31,30,31,176,31,40,31,25,31,105,31,105,30,175,31,28,31,176,31,166,31,100,31,5,31,145,31,130,31,163,31,34,31,34,30,37,31,49,31,78,31,78,30,78,29,232,31,85,31,85,30,19,31,89,31,89,30,111,31,154,31,88,31,88,30,8,31,160,31,141,31,51,31,46,31,46,30,165,31,165,30,27,31,236,31,83,31,225,31,225,30,217,31,50,31,216,31,216,30,40,31,159,31,107,31,107,30,109,31,90,31,127,31,127,30,230,31,230,30,230,29,230,28,230,27,144,31,106,31,65,31,149,31,194,31,21,31,215,31,13,31,156,31,46,31,183,31,98,31,222,31,222,30,222,29,222,28,133,31,209,31,223,31,223,30,149,31,80,31,49,31,42,31,120,31,120,30,203,31,203,30,54,31,9,31,216,31,148,31,251,31,250,31,147,31,31,31,165,31,165,30,165,31,94,31,160,31,84,31,105,31,240,31,240,30,133,31,105,31,62,31,126,31,126,30,48,31,64,31,88,31,226,31,28,31,28,30,17,31,24,31,69,31,7,31,7,30,7,29,7,28,233,31,233,30,233,29,211,31,211,30,60,31,116,31,116,30,21,31,142,31,235,31,32,31,49,31,109,31,109,30,173,31,114,31,42,31,193,31,193,30,220,31,220,30,47,31,221,31,102,31,196,31,30,31,15,31,117,31,117,30,95,31,170,31,170,30,170,29,62,31,237,31,237,30,41,31,122,31,5,31,71,31,110,31,37,31,116,31,151,31,114,31,219,31,24,31,105,31,249,31,230,31,230,30,246,31,215,31,215,30,80,31,246,31,195,31,107,31,197,31,197,30,127,31,75,31,224,31,58,31,248,31,176,31,111,31,111,30,191,31,42,31,42,30,144,31,62,31,62,30,29,31,156,31,223,31,253,31,63,31,53,31,129,31,231,31,82,31,150,31,150,30,150,29,21,31,188,31,83,31,83,30,137,31,241,31,170,31,230,31,25,31,197,31,113,31,113,30,139,31,139,30,196,31,202,31,170,31,170,30,180,31,180,30,180,29,87,31,176,31,204,31,204,30,233,31,103,31,131,31,131,30,94,31,109,31,109,30,43,31,153,31,124,31,4,31,245,31,251,31,251,30,131,31,228,31,228,30,147,31,147,30,123,31,31,31,65,31,13,31,155,31,148,31,44,31,44,30,44,29,135,31,237,31,218,31,218,30,218,29,30,31,140,31,37,31,43,31,40,31,122,31,122,30,51,31,9,31,30,31,98,31,83,31,94,31,51,31,51,30,226,31,58,31,96,31,49,31,206,31,208,31,40,31,40,30,218,31,217,31,171,31,14,31,225,31,225,30,225,29,230,31,57,31,124,31,206,31,21,31,35,31,35,30,127,31,24,31,144,31,53,31,198,31,76,31,76,30,38,31,214,31,214,30,78,31,87,31,149,31,199,31,69,31,147,31,162,31,200,31,200,30,216,31,163,31,163,30,215,31,19,31,233,31,233,30,218,31,97,31,199,31,108,31,108,30,144,31,4,31,104,31,91,31,91,30,91,29,40,31,206,31,206,30,78,31,113,31,238,31,35,31,88,31,157,31,107,31,52,31,79,31,79,30,96,31,8,31,99,31,57,31,57,30,238,31,16,31,35,31,35,30,206,31,8,31,12,31,173,31,173,30,224,31,104,31,4,31,78,31,92,31,189,31,205,31,22,31,92,31,92,30,23,31,23,30,23,29,164,31,207,31,118,31,39,31,190,31,238,31,238,30,91,31,250,31,189,31,225,31,145,31,242,31,242,30,242,29,174,31,145,31,231,31,8,31,8,30,203,31,237,31,82,31,26,31,26,30,235,31,154,31,190,31,14,31,193,31,86,31,203,31,182,31,120,31,154,31,154,30,154,29,40,31,200,31,200,30,153,31,212,31,212,30,212,29,212,28,65,31,114,31,46,31,66,31,66,30,213,31,213,30,213,29,74,31,74,30,74,29,206,31,244,31,185,31,204,31,148,31,148,30,148,29,111,31,177,31,174,31,83,31,176,31,40,31,40,30,119,31,18,31,18,30,122,31,23,31,190,31,220,31,178,31,222,31,76,31,35,31,98,31,219,31,153,31,177,31,50,31,50,30,50,29,210,31,13,31,252,31,117,31,202,31,145,31,235,31,235,30,235,29,38,31,133,31,226,31,68,31,73,31,73,30,118,31,201,31,109,31,12,31,12,30,46,31,203,31,203,30,87,31,147,31,147,30,232,31,178,31,23,31,61,31,61,30,130,31,92,31,92,30,110,31,207,31,207,30,207,29,72,31,234,31,234,30,234,29,77,31,78,31,78,30,78,29,78,28,22,31,187,31,122,31,10,31,171,31,57,31,138,31,67,31,56,31,56,30,56,29,56,28,61,31,61,30,103,31,103,30,57,31,132,31,144,31,194,31,27,31,27,30,17,31,5,31,92,31,173,31,195,31,2,31,218,31,109,31,26,31,26,30,73,31,48,31,63,31,119,31,67,31,70,31,171,31,208,31,8,31,15,31,58,31,5,31,5,30,217,31,211,31,211,30,69,31,84,31,84,30,231,31,118,31,71,31,242,31,129,31,129,30,155,31,150,31,41,31,228,31,250,31,73,31,227,31,39,31,92,31,238,31,11,31,41,31,212,31,212,31,212,30,212,29,134,31,75,31,75,30,197,31,14,31,139,31,103,31,103,30,240,31,1,31,36,31,123,31,123,30,8,31,1,31,1,30,212,31,24,31,10,31,201,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
