-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 365;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,56,0,186,0,92,0,6,0,10,0,169,0,4,0,140,0,0,0,36,0,0,0,250,0,161,0,223,0,0,0,225,0,74,0,195,0,35,0,229,0,34,0,155,0,228,0,173,0,202,0,89,0,238,0,118,0,0,0,230,0,190,0,142,0,0,0,0,0,120,0,34,0,23,0,35,0,171,0,150,0,8,0,6,0,85,0,95,0,80,0,163,0,0,0,94,0,0,0,19,0,212,0,79,0,0,0,209,0,0,0,171,0,108,0,222,0,115,0,159,0,131,0,20,0,93,0,171,0,139,0,53,0,0,0,29,0,183,0,0,0,246,0,51,0,9,0,9,0,49,0,160,0,100,0,0,0,62,0,18,0,121,0,42,0,0,0,31,0,45,0,0,0,232,0,0,0,190,0,192,0,16,0,0,0,0,0,223,0,199,0,151,0,48,0,61,0,0,0,206,0,0,0,115,0,189,0,0,0,234,0,186,0,1,0,203,0,78,0,0,0,0,0,0,0,22,0,196,0,236,0,109,0,91,0,0,0,198,0,0,0,0,0,98,0,187,0,70,0,71,0,162,0,225,0,228,0,100,0,197,0,64,0,0,0,124,0,41,0,250,0,9,0,0,0,50,0,120,0,0,0,225,0,71,0,67,0,133,0,39,0,78,0,234,0,253,0,163,0,9,0,119,0,0,0,0,0,0,0,32,0,198,0,0,0,63,0,77,0,142,0,73,0,145,0,212,0,89,0,79,0,174,0,183,0,152,0,54,0,236,0,200,0,57,0,213,0,175,0,221,0,49,0,249,0,19,0,220,0,22,0,254,0,155,0,215,0,0,0,220,0,0,0,142,0,174,0,89,0,0,0,62,0,128,0,123,0,196,0,200,0,0,0,0,0,10,0,0,0,0,0,216,0,225,0,192,0,152,0,239,0,245,0,0,0,27,0,0,0,139,0,167,0,52,0,0,0,100,0,236,0,107,0,107,0,174,0,32,0,0,0,0,0,0,0,158,0,53,0,241,0,189,0,89,0,194,0,239,0,75,0,17,0,233,0,233,0,143,0,155,0,0,0,0,0,213,0,8,0,31,0,19,0,252,0,0,0,197,0,128,0,97,0,209,0,108,0,190,0,168,0,199,0,138,0,97,0,0,0,240,0,109,0,0,0,0,0,15,0,0,0,0,0,67,0,85,0,90,0,133,0,0,0,80,0,115,0,181,0,227,0,26,0,165,0,217,0,39,0,0,0,227,0,229,0,192,0,155,0,0,0,115,0,212,0,14,0,186,0,131,0,50,0,122,0,219,0,75,0,0,0,155,0,49,0,133,0,199,0,0,0,0,0,251,0,0,0,145,0,0,0,142,0,0,0,131,0,211,0,132,0,0,0,151,0,187,0,59,0,127,0,81,0,245,0,231,0,23,0,158,0,0,0,241,0,155,0,128,0,198,0,0,0,0,0,87,0,7,0,22,0,205,0,27,0,0,0,0,0,81,0,61,0,214,0,25,0,198,0,151,0,32,0,122,0,101,0,0,0,141,0,7,0,161,0,236,0,44,0,242,0,217,0,13,0,71,0,0,0,208,0,254,0,209,0,189,0,247,0,145,0,198,0,35,0,123,0,206,0,69,0,125,0,217,0,0,0,62,0);
signal scenario_full  : scenario_type := (0,0,56,31,186,31,92,31,6,31,10,31,169,31,4,31,140,31,140,30,36,31,36,30,250,31,161,31,223,31,223,30,225,31,74,31,195,31,35,31,229,31,34,31,155,31,228,31,173,31,202,31,89,31,238,31,118,31,118,30,230,31,190,31,142,31,142,30,142,29,120,31,34,31,23,31,35,31,171,31,150,31,8,31,6,31,85,31,95,31,80,31,163,31,163,30,94,31,94,30,19,31,212,31,79,31,79,30,209,31,209,30,171,31,108,31,222,31,115,31,159,31,131,31,20,31,93,31,171,31,139,31,53,31,53,30,29,31,183,31,183,30,246,31,51,31,9,31,9,31,49,31,160,31,100,31,100,30,62,31,18,31,121,31,42,31,42,30,31,31,45,31,45,30,232,31,232,30,190,31,192,31,16,31,16,30,16,29,223,31,199,31,151,31,48,31,61,31,61,30,206,31,206,30,115,31,189,31,189,30,234,31,186,31,1,31,203,31,78,31,78,30,78,29,78,28,22,31,196,31,236,31,109,31,91,31,91,30,198,31,198,30,198,29,98,31,187,31,70,31,71,31,162,31,225,31,228,31,100,31,197,31,64,31,64,30,124,31,41,31,250,31,9,31,9,30,50,31,120,31,120,30,225,31,71,31,67,31,133,31,39,31,78,31,234,31,253,31,163,31,9,31,119,31,119,30,119,29,119,28,32,31,198,31,198,30,63,31,77,31,142,31,73,31,145,31,212,31,89,31,79,31,174,31,183,31,152,31,54,31,236,31,200,31,57,31,213,31,175,31,221,31,49,31,249,31,19,31,220,31,22,31,254,31,155,31,215,31,215,30,220,31,220,30,142,31,174,31,89,31,89,30,62,31,128,31,123,31,196,31,200,31,200,30,200,29,10,31,10,30,10,29,216,31,225,31,192,31,152,31,239,31,245,31,245,30,27,31,27,30,139,31,167,31,52,31,52,30,100,31,236,31,107,31,107,31,174,31,32,31,32,30,32,29,32,28,158,31,53,31,241,31,189,31,89,31,194,31,239,31,75,31,17,31,233,31,233,31,143,31,155,31,155,30,155,29,213,31,8,31,31,31,19,31,252,31,252,30,197,31,128,31,97,31,209,31,108,31,190,31,168,31,199,31,138,31,97,31,97,30,240,31,109,31,109,30,109,29,15,31,15,30,15,29,67,31,85,31,90,31,133,31,133,30,80,31,115,31,181,31,227,31,26,31,165,31,217,31,39,31,39,30,227,31,229,31,192,31,155,31,155,30,115,31,212,31,14,31,186,31,131,31,50,31,122,31,219,31,75,31,75,30,155,31,49,31,133,31,199,31,199,30,199,29,251,31,251,30,145,31,145,30,142,31,142,30,131,31,211,31,132,31,132,30,151,31,187,31,59,31,127,31,81,31,245,31,231,31,23,31,158,31,158,30,241,31,155,31,128,31,198,31,198,30,198,29,87,31,7,31,22,31,205,31,27,31,27,30,27,29,81,31,61,31,214,31,25,31,198,31,151,31,32,31,122,31,101,31,101,30,141,31,7,31,161,31,236,31,44,31,242,31,217,31,13,31,71,31,71,30,208,31,254,31,209,31,189,31,247,31,145,31,198,31,35,31,123,31,206,31,69,31,125,31,217,31,217,30,62,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
