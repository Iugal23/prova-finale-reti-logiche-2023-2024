-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_747 is
end project_tb_747;

architecture project_tb_arch_747 of project_tb_747 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 779;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (156,0,81,0,54,0,105,0,152,0,0,0,251,0,14,0,148,0,118,0,218,0,5,0,248,0,176,0,0,0,143,0,0,0,209,0,234,0,139,0,194,0,84,0,192,0,196,0,141,0,69,0,195,0,50,0,122,0,5,0,58,0,203,0,0,0,168,0,118,0,234,0,141,0,211,0,17,0,0,0,126,0,202,0,0,0,31,0,21,0,139,0,0,0,0,0,216,0,161,0,219,0,213,0,44,0,0,0,124,0,253,0,162,0,180,0,240,0,0,0,88,0,198,0,103,0,203,0,49,0,213,0,247,0,36,0,154,0,0,0,98,0,0,0,232,0,57,0,28,0,0,0,255,0,77,0,0,0,0,0,119,0,150,0,209,0,98,0,205,0,0,0,181,0,186,0,79,0,29,0,0,0,66,0,0,0,250,0,208,0,160,0,68,0,45,0,87,0,62,0,72,0,58,0,64,0,224,0,53,0,148,0,44,0,214,0,51,0,182,0,0,0,13,0,10,0,0,0,170,0,0,0,229,0,213,0,190,0,21,0,190,0,0,0,34,0,127,0,0,0,0,0,97,0,0,0,19,0,223,0,40,0,69,0,0,0,207,0,167,0,148,0,84,0,214,0,46,0,36,0,143,0,175,0,62,0,235,0,12,0,0,0,0,0,118,0,0,0,0,0,215,0,33,0,114,0,130,0,0,0,50,0,148,0,152,0,136,0,151,0,0,0,33,0,0,0,199,0,182,0,184,0,0,0,54,0,0,0,24,0,13,0,145,0,40,0,214,0,243,0,177,0,187,0,120,0,127,0,222,0,0,0,21,0,101,0,31,0,0,0,189,0,174,0,0,0,107,0,22,0,138,0,158,0,253,0,39,0,111,0,8,0,40,0,95,0,28,0,200,0,27,0,173,0,0,0,166,0,90,0,56,0,0,0,121,0,73,0,43,0,0,0,99,0,47,0,90,0,168,0,0,0,0,0,237,0,86,0,0,0,251,0,77,0,99,0,194,0,112,0,0,0,19,0,0,0,140,0,14,0,197,0,173,0,159,0,0,0,0,0,225,0,120,0,90,0,21,0,205,0,0,0,108,0,10,0,179,0,251,0,171,0,31,0,94,0,21,0,149,0,135,0,0,0,159,0,0,0,218,0,65,0,153,0,211,0,209,0,233,0,197,0,110,0,78,0,97,0,0,0,63,0,207,0,161,0,145,0,247,0,68,0,211,0,44,0,205,0,155,0,121,0,8,0,81,0,207,0,0,0,133,0,78,0,168,0,0,0,0,0,0,0,0,0,0,0,0,0,0,0,208,0,8,0,245,0,142,0,104,0,0,0,0,0,140,0,179,0,197,0,13,0,180,0,0,0,205,0,28,0,0,0,220,0,66,0,64,0,23,0,159,0,0,0,0,0,147,0,23,0,82,0,188,0,133,0,95,0,0,0,21,0,4,0,77,0,119,0,0,0,118,0,16,0,0,0,61,0,15,0,0,0,79,0,232,0,93,0,0,0,95,0,67,0,203,0,166,0,130,0,144,0,50,0,187,0,248,0,97,0,235,0,203,0,122,0,0,0,145,0,84,0,22,0,0,0,208,0,76,0,92,0,57,0,0,0,132,0,90,0,225,0,54,0,121,0,54,0,0,0,192,0,192,0,246,0,0,0,83,0,0,0,199,0,196,0,50,0,0,0,65,0,207,0,0,0,174,0,246,0,25,0,163,0,31,0,0,0,137,0,245,0,92,0,162,0,159,0,228,0,0,0,104,0,86,0,12,0,35,0,24,0,171,0,87,0,208,0,230,0,104,0,122,0,33,0,188,0,63,0,147,0,248,0,28,0,0,0,29,0,0,0,161,0,133,0,98,0,205,0,0,0,40,0,11,0,188,0,0,0,83,0,195,0,0,0,0,0,228,0,0,0,166,0,49,0,200,0,68,0,42,0,20,0,47,0,238,0,226,0,0,0,151,0,0,0,0,0,0,0,46,0,144,0,121,0,44,0,236,0,180,0,75,0,0,0,0,0,165,0,64,0,181,0,144,0,0,0,207,0,85,0,172,0,77,0,168,0,12,0,12,0,0,0,218,0,83,0,152,0,85,0,14,0,224,0,114,0,225,0,7,0,107,0,104,0,234,0,245,0,85,0,75,0,65,0,0,0,36,0,0,0,53,0,236,0,121,0,228,0,78,0,39,0,0,0,0,0,98,0,108,0,181,0,205,0,0,0,0,0,84,0,208,0,61,0,0,0,133,0,29,0,201,0,37,0,120,0,69,0,85,0,113,0,140,0,0,0,253,0,118,0,169,0,112,0,54,0,18,0,96,0,129,0,0,0,61,0,0,0,0,0,133,0,113,0,0,0,0,0,75,0,0,0,245,0,0,0,237,0,118,0,130,0,0,0,168,0,231,0,226,0,216,0,24,0,22,0,175,0,0,0,117,0,239,0,48,0,226,0,248,0,78,0,202,0,214,0,198,0,5,0,0,0,0,0,71,0,51,0,10,0,195,0,75,0,128,0,160,0,0,0,144,0,233,0,87,0,159,0,197,0,87,0,164,0,167,0,148,0,240,0,0,0,142,0,78,0,29,0,29,0,0,0,180,0,138,0,11,0,0,0,0,0,24,0,249,0,102,0,224,0,72,0,133,0,0,0,0,0,240,0,204,0,230,0,29,0,78,0,201,0,137,0,224,0,244,0,36,0,101,0,133,0,180,0,48,0,68,0,0,0,0,0,34,0,176,0,0,0,76,0,183,0,0,0,209,0,46,0,217,0,196,0,169,0,126,0,130,0,180,0,62,0,0,0,184,0,82,0,199,0,165,0,0,0,93,0,173,0,153,0,0,0,117,0,134,0,0,0,170,0,0,0,185,0,42,0,230,0,253,0,182,0,56,0,209,0,0,0,222,0,252,0,151,0,50,0,179,0,0,0,93,0,161,0,21,0,0,0,89,0,147,0,215,0,250,0,197,0,0,0,137,0,156,0,154,0,0,0,59,0,23,0,124,0,0,0,0,0,231,0,0,0,221,0,112,0,69,0,25,0,167,0,0,0,202,0,0,0,101,0,70,0,0,0,0,0,233,0,0,0,107,0,180,0,0,0,7,0,33,0,125,0,0,0,0,0,0,0,0,0,0,0,0,0,156,0,0,0,74,0,145,0,179,0,80,0,196,0,177,0,60,0,99,0,0,0,159,0,117,0,150,0,67,0,210,0,166,0,0,0,60,0,0,0,92,0,183,0,172,0,26,0,45,0,80,0,0,0,172,0,153,0,107,0,214,0,0,0,130,0,142,0,116,0,0,0,228,0,173,0,203,0,39,0,62,0,116,0,2,0,0,0,141,0,47,0,245,0,229,0,7,0,194,0,6,0,0,0,3,0,167,0,156,0,247,0,172,0,255,0,56,0,130,0,53,0,214,0,45,0,16,0,0,0,0,0,150,0,46,0,111,0,203,0,37,0,96,0,235,0,133,0,4,0,171,0,33,0,0,0,147,0,88,0,14,0);
signal scenario_full  : scenario_type := (156,31,81,31,54,31,105,31,152,31,152,30,251,31,14,31,148,31,118,31,218,31,5,31,248,31,176,31,176,30,143,31,143,30,209,31,234,31,139,31,194,31,84,31,192,31,196,31,141,31,69,31,195,31,50,31,122,31,5,31,58,31,203,31,203,30,168,31,118,31,234,31,141,31,211,31,17,31,17,30,126,31,202,31,202,30,31,31,21,31,139,31,139,30,139,29,216,31,161,31,219,31,213,31,44,31,44,30,124,31,253,31,162,31,180,31,240,31,240,30,88,31,198,31,103,31,203,31,49,31,213,31,247,31,36,31,154,31,154,30,98,31,98,30,232,31,57,31,28,31,28,30,255,31,77,31,77,30,77,29,119,31,150,31,209,31,98,31,205,31,205,30,181,31,186,31,79,31,29,31,29,30,66,31,66,30,250,31,208,31,160,31,68,31,45,31,87,31,62,31,72,31,58,31,64,31,224,31,53,31,148,31,44,31,214,31,51,31,182,31,182,30,13,31,10,31,10,30,170,31,170,30,229,31,213,31,190,31,21,31,190,31,190,30,34,31,127,31,127,30,127,29,97,31,97,30,19,31,223,31,40,31,69,31,69,30,207,31,167,31,148,31,84,31,214,31,46,31,36,31,143,31,175,31,62,31,235,31,12,31,12,30,12,29,118,31,118,30,118,29,215,31,33,31,114,31,130,31,130,30,50,31,148,31,152,31,136,31,151,31,151,30,33,31,33,30,199,31,182,31,184,31,184,30,54,31,54,30,24,31,13,31,145,31,40,31,214,31,243,31,177,31,187,31,120,31,127,31,222,31,222,30,21,31,101,31,31,31,31,30,189,31,174,31,174,30,107,31,22,31,138,31,158,31,253,31,39,31,111,31,8,31,40,31,95,31,28,31,200,31,27,31,173,31,173,30,166,31,90,31,56,31,56,30,121,31,73,31,43,31,43,30,99,31,47,31,90,31,168,31,168,30,168,29,237,31,86,31,86,30,251,31,77,31,99,31,194,31,112,31,112,30,19,31,19,30,140,31,14,31,197,31,173,31,159,31,159,30,159,29,225,31,120,31,90,31,21,31,205,31,205,30,108,31,10,31,179,31,251,31,171,31,31,31,94,31,21,31,149,31,135,31,135,30,159,31,159,30,218,31,65,31,153,31,211,31,209,31,233,31,197,31,110,31,78,31,97,31,97,30,63,31,207,31,161,31,145,31,247,31,68,31,211,31,44,31,205,31,155,31,121,31,8,31,81,31,207,31,207,30,133,31,78,31,168,31,168,30,168,29,168,28,168,27,168,26,168,25,168,24,208,31,8,31,245,31,142,31,104,31,104,30,104,29,140,31,179,31,197,31,13,31,180,31,180,30,205,31,28,31,28,30,220,31,66,31,64,31,23,31,159,31,159,30,159,29,147,31,23,31,82,31,188,31,133,31,95,31,95,30,21,31,4,31,77,31,119,31,119,30,118,31,16,31,16,30,61,31,15,31,15,30,79,31,232,31,93,31,93,30,95,31,67,31,203,31,166,31,130,31,144,31,50,31,187,31,248,31,97,31,235,31,203,31,122,31,122,30,145,31,84,31,22,31,22,30,208,31,76,31,92,31,57,31,57,30,132,31,90,31,225,31,54,31,121,31,54,31,54,30,192,31,192,31,246,31,246,30,83,31,83,30,199,31,196,31,50,31,50,30,65,31,207,31,207,30,174,31,246,31,25,31,163,31,31,31,31,30,137,31,245,31,92,31,162,31,159,31,228,31,228,30,104,31,86,31,12,31,35,31,24,31,171,31,87,31,208,31,230,31,104,31,122,31,33,31,188,31,63,31,147,31,248,31,28,31,28,30,29,31,29,30,161,31,133,31,98,31,205,31,205,30,40,31,11,31,188,31,188,30,83,31,195,31,195,30,195,29,228,31,228,30,166,31,49,31,200,31,68,31,42,31,20,31,47,31,238,31,226,31,226,30,151,31,151,30,151,29,151,28,46,31,144,31,121,31,44,31,236,31,180,31,75,31,75,30,75,29,165,31,64,31,181,31,144,31,144,30,207,31,85,31,172,31,77,31,168,31,12,31,12,31,12,30,218,31,83,31,152,31,85,31,14,31,224,31,114,31,225,31,7,31,107,31,104,31,234,31,245,31,85,31,75,31,65,31,65,30,36,31,36,30,53,31,236,31,121,31,228,31,78,31,39,31,39,30,39,29,98,31,108,31,181,31,205,31,205,30,205,29,84,31,208,31,61,31,61,30,133,31,29,31,201,31,37,31,120,31,69,31,85,31,113,31,140,31,140,30,253,31,118,31,169,31,112,31,54,31,18,31,96,31,129,31,129,30,61,31,61,30,61,29,133,31,113,31,113,30,113,29,75,31,75,30,245,31,245,30,237,31,118,31,130,31,130,30,168,31,231,31,226,31,216,31,24,31,22,31,175,31,175,30,117,31,239,31,48,31,226,31,248,31,78,31,202,31,214,31,198,31,5,31,5,30,5,29,71,31,51,31,10,31,195,31,75,31,128,31,160,31,160,30,144,31,233,31,87,31,159,31,197,31,87,31,164,31,167,31,148,31,240,31,240,30,142,31,78,31,29,31,29,31,29,30,180,31,138,31,11,31,11,30,11,29,24,31,249,31,102,31,224,31,72,31,133,31,133,30,133,29,240,31,204,31,230,31,29,31,78,31,201,31,137,31,224,31,244,31,36,31,101,31,133,31,180,31,48,31,68,31,68,30,68,29,34,31,176,31,176,30,76,31,183,31,183,30,209,31,46,31,217,31,196,31,169,31,126,31,130,31,180,31,62,31,62,30,184,31,82,31,199,31,165,31,165,30,93,31,173,31,153,31,153,30,117,31,134,31,134,30,170,31,170,30,185,31,42,31,230,31,253,31,182,31,56,31,209,31,209,30,222,31,252,31,151,31,50,31,179,31,179,30,93,31,161,31,21,31,21,30,89,31,147,31,215,31,250,31,197,31,197,30,137,31,156,31,154,31,154,30,59,31,23,31,124,31,124,30,124,29,231,31,231,30,221,31,112,31,69,31,25,31,167,31,167,30,202,31,202,30,101,31,70,31,70,30,70,29,233,31,233,30,107,31,180,31,180,30,7,31,33,31,125,31,125,30,125,29,125,28,125,27,125,26,125,25,156,31,156,30,74,31,145,31,179,31,80,31,196,31,177,31,60,31,99,31,99,30,159,31,117,31,150,31,67,31,210,31,166,31,166,30,60,31,60,30,92,31,183,31,172,31,26,31,45,31,80,31,80,30,172,31,153,31,107,31,214,31,214,30,130,31,142,31,116,31,116,30,228,31,173,31,203,31,39,31,62,31,116,31,2,31,2,30,141,31,47,31,245,31,229,31,7,31,194,31,6,31,6,30,3,31,167,31,156,31,247,31,172,31,255,31,56,31,130,31,53,31,214,31,45,31,16,31,16,30,16,29,150,31,46,31,111,31,203,31,37,31,96,31,235,31,133,31,4,31,171,31,33,31,33,30,147,31,88,31,14,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
