-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 212;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (74,0,80,0,0,0,57,0,0,0,85,0,40,0,83,0,85,0,15,0,0,0,0,0,102,0,0,0,0,0,0,0,80,0,164,0,124,0,232,0,119,0,125,0,0,0,86,0,22,0,246,0,240,0,44,0,0,0,0,0,0,0,127,0,238,0,113,0,0,0,190,0,80,0,127,0,234,0,248,0,151,0,160,0,154,0,152,0,165,0,180,0,32,0,176,0,208,0,223,0,96,0,185,0,236,0,186,0,63,0,0,0,88,0,0,0,61,0,13,0,0,0,0,0,90,0,0,0,91,0,180,0,235,0,25,0,0,0,85,0,151,0,234,0,0,0,66,0,105,0,6,0,14,0,14,0,63,0,213,0,187,0,0,0,236,0,141,0,136,0,2,0,89,0,0,0,231,0,127,0,63,0,75,0,0,0,234,0,236,0,0,0,90,0,103,0,126,0,0,0,0,0,0,0,101,0,0,0,128,0,138,0,3,0,0,0,6,0,119,0,255,0,163,0,233,0,0,0,231,0,24,0,225,0,7,0,69,0,214,0,0,0,63,0,32,0,36,0,195,0,137,0,46,0,86,0,159,0,148,0,32,0,225,0,216,0,64,0,196,0,194,0,231,0,151,0,204,0,42,0,93,0,150,0,251,0,73,0,241,0,23,0,145,0,87,0,49,0,81,0,223,0,87,0,206,0,86,0,0,0,104,0,26,0,0,0,95,0,213,0,185,0,0,0,77,0,150,0,0,0,37,0,131,0,52,0,0,0,135,0,165,0,19,0,0,0,62,0,40,0,189,0,82,0,70,0,173,0,254,0,60,0,199,0,0,0,147,0,105,0,214,0,0,0,0,0,201,0,113,0,207,0,0,0,97,0,0,0,190,0,48,0,251,0,207,0,45,0,228,0,138,0,0,0,0,0,118,0,234,0,228,0,14,0,217,0,0,0,42,0,0,0,73,0);
signal scenario_full  : scenario_type := (74,31,80,31,80,30,57,31,57,30,85,31,40,31,83,31,85,31,15,31,15,30,15,29,102,31,102,30,102,29,102,28,80,31,164,31,124,31,232,31,119,31,125,31,125,30,86,31,22,31,246,31,240,31,44,31,44,30,44,29,44,28,127,31,238,31,113,31,113,30,190,31,80,31,127,31,234,31,248,31,151,31,160,31,154,31,152,31,165,31,180,31,32,31,176,31,208,31,223,31,96,31,185,31,236,31,186,31,63,31,63,30,88,31,88,30,61,31,13,31,13,30,13,29,90,31,90,30,91,31,180,31,235,31,25,31,25,30,85,31,151,31,234,31,234,30,66,31,105,31,6,31,14,31,14,31,63,31,213,31,187,31,187,30,236,31,141,31,136,31,2,31,89,31,89,30,231,31,127,31,63,31,75,31,75,30,234,31,236,31,236,30,90,31,103,31,126,31,126,30,126,29,126,28,101,31,101,30,128,31,138,31,3,31,3,30,6,31,119,31,255,31,163,31,233,31,233,30,231,31,24,31,225,31,7,31,69,31,214,31,214,30,63,31,32,31,36,31,195,31,137,31,46,31,86,31,159,31,148,31,32,31,225,31,216,31,64,31,196,31,194,31,231,31,151,31,204,31,42,31,93,31,150,31,251,31,73,31,241,31,23,31,145,31,87,31,49,31,81,31,223,31,87,31,206,31,86,31,86,30,104,31,26,31,26,30,95,31,213,31,185,31,185,30,77,31,150,31,150,30,37,31,131,31,52,31,52,30,135,31,165,31,19,31,19,30,62,31,40,31,189,31,82,31,70,31,173,31,254,31,60,31,199,31,199,30,147,31,105,31,214,31,214,30,214,29,201,31,113,31,207,31,207,30,97,31,97,30,190,31,48,31,251,31,207,31,45,31,228,31,138,31,138,30,138,29,118,31,234,31,228,31,14,31,217,31,217,30,42,31,42,30,73,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
