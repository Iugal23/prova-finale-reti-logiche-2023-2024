-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 784;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,196,0,120,0,24,0,203,0,0,0,214,0,158,0,92,0,13,0,144,0,139,0,154,0,46,0,47,0,150,0,231,0,0,0,168,0,29,0,0,0,139,0,245,0,105,0,0,0,0,0,28,0,234,0,103,0,0,0,0,0,171,0,179,0,0,0,118,0,33,0,188,0,0,0,0,0,239,0,0,0,128,0,2,0,6,0,213,0,127,0,0,0,99,0,0,0,218,0,118,0,246,0,0,0,28,0,72,0,213,0,197,0,170,0,78,0,0,0,223,0,102,0,174,0,0,0,63,0,135,0,158,0,81,0,199,0,8,0,0,0,183,0,141,0,0,0,0,0,90,0,42,0,0,0,207,0,132,0,210,0,0,0,167,0,250,0,152,0,239,0,192,0,91,0,0,0,179,0,18,0,158,0,216,0,22,0,75,0,2,0,138,0,0,0,0,0,188,0,118,0,173,0,33,0,216,0,210,0,164,0,45,0,65,0,0,0,193,0,84,0,93,0,215,0,208,0,62,0,40,0,0,0,234,0,199,0,0,0,86,0,0,0,120,0,0,0,0,0,93,0,240,0,164,0,167,0,0,0,227,0,71,0,244,0,120,0,56,0,0,0,235,0,0,0,255,0,250,0,49,0,41,0,181,0,0,0,66,0,238,0,110,0,73,0,0,0,247,0,145,0,149,0,4,0,202,0,99,0,139,0,164,0,173,0,0,0,16,0,151,0,4,0,178,0,241,0,127,0,129,0,230,0,239,0,175,0,0,0,47,0,0,0,169,0,10,0,83,0,0,0,140,0,72,0,13,0,0,0,48,0,0,0,23,0,0,0,77,0,131,0,0,0,224,0,82,0,164,0,255,0,252,0,3,0,0,0,163,0,218,0,0,0,11,0,245,0,216,0,232,0,116,0,8,0,47,0,42,0,124,0,193,0,37,0,0,0,64,0,7,0,1,0,240,0,57,0,223,0,215,0,0,0,12,0,125,0,202,0,0,0,0,0,108,0,68,0,184,0,219,0,45,0,146,0,223,0,225,0,0,0,0,0,0,0,69,0,106,0,103,0,216,0,0,0,209,0,48,0,153,0,0,0,192,0,149,0,188,0,67,0,85,0,204,0,250,0,185,0,147,0,116,0,242,0,0,0,165,0,103,0,215,0,5,0,0,0,141,0,253,0,154,0,164,0,14,0,9,0,222,0,0,0,129,0,142,0,0,0,0,0,180,0,0,0,201,0,13,0,240,0,40,0,252,0,26,0,122,0,245,0,139,0,128,0,0,0,128,0,139,0,64,0,253,0,81,0,216,0,0,0,18,0,199,0,81,0,107,0,46,0,0,0,23,0,0,0,154,0,201,0,95,0,120,0,148,0,26,0,51,0,0,0,36,0,21,0,14,0,0,0,218,0,14,0,201,0,0,0,144,0,0,0,196,0,104,0,0,0,231,0,216,0,179,0,96,0,63,0,41,0,87,0,0,0,60,0,239,0,197,0,253,0,92,0,249,0,103,0,205,0,101,0,30,0,184,0,0,0,73,0,98,0,14,0,42,0,254,0,129,0,248,0,199,0,30,0,249,0,17,0,189,0,188,0,0,0,0,0,168,0,0,0,0,0,55,0,185,0,67,0,73,0,101,0,0,0,242,0,94,0,0,0,0,0,46,0,55,0,133,0,32,0,235,0,111,0,7,0,156,0,199,0,245,0,73,0,253,0,0,0,0,0,207,0,115,0,209,0,53,0,23,0,15,0,0,0,73,0,156,0,114,0,66,0,41,0,102,0,8,0,0,0,66,0,230,0,151,0,199,0,0,0,54,0,69,0,0,0,108,0,170,0,146,0,83,0,207,0,205,0,230,0,252,0,0,0,210,0,31,0,165,0,153,0,243,0,0,0,20,0,243,0,0,0,77,0,122,0,68,0,0,0,0,0,15,0,227,0,68,0,250,0,22,0,145,0,0,0,61,0,104,0,220,0,241,0,98,0,0,0,0,0,0,0,0,0,0,0,153,0,0,0,199,0,125,0,84,0,174,0,236,0,208,0,245,0,129,0,0,0,149,0,65,0,82,0,83,0,179,0,123,0,192,0,14,0,0,0,199,0,85,0,144,0,233,0,111,0,90,0,0,0,46,0,93,0,49,0,12,0,225,0,239,0,125,0,171,0,214,0,82,0,137,0,30,0,204,0,0,0,15,0,182,0,51,0,25,0,129,0,182,0,135,0,163,0,0,0,20,0,130,0,117,0,39,0,119,0,198,0,153,0,34,0,235,0,6,0,0,0,36,0,0,0,70,0,159,0,215,0,0,0,19,0,0,0,187,0,2,0,0,0,99,0,176,0,91,0,0,0,0,0,255,0,172,0,0,0,181,0,207,0,191,0,206,0,95,0,185,0,1,0,10,0,245,0,108,0,231,0,255,0,177,0,132,0,117,0,105,0,242,0,216,0,0,0,0,0,0,0,0,0,204,0,136,0,242,0,241,0,165,0,198,0,0,0,144,0,143,0,149,0,84,0,73,0,250,0,51,0,134,0,139,0,205,0,206,0,253,0,0,0,233,0,7,0,0,0,0,0,174,0,0,0,0,0,248,0,212,0,100,0,30,0,146,0,0,0,0,0,235,0,23,0,52,0,8,0,0,0,0,0,74,0,210,0,162,0,206,0,175,0,203,0,110,0,124,0,0,0,155,0,223,0,225,0,141,0,105,0,227,0,142,0,177,0,220,0,197,0,177,0,0,0,128,0,77,0,0,0,127,0,0,0,0,0,39,0,151,0,88,0,98,0,0,0,191,0,0,0,14,0,23,0,250,0,0,0,0,0,120,0,0,0,0,0,220,0,154,0,0,0,249,0,234,0,179,0,180,0,104,0,0,0,0,0,13,0,124,0,135,0,48,0,78,0,0,0,0,0,72,0,242,0,150,0,158,0,193,0,182,0,0,0,191,0,0,0,98,0,2,0,130,0,70,0,177,0,238,0,111,0,140,0,89,0,91,0,0,0,162,0,90,0,0,0,0,0,169,0,120,0,37,0,133,0,153,0,142,0,241,0,37,0,232,0,28,0,245,0,147,0,54,0,245,0,207,0,192,0,221,0,55,0,129,0,118,0,221,0,83,0,99,0,0,0,49,0,142,0,241,0,95,0,145,0,75,0,137,0,173,0,0,0,223,0,181,0,208,0,118,0,195,0,41,0,202,0,152,0,137,0,80,0,67,0,34,0,129,0,3,0,11,0,255,0,57,0,85,0,0,0,124,0,157,0,0,0,145,0,7,0,174,0,145,0,129,0,216,0,172,0,60,0,227,0,0,0,216,0,173,0,49,0,207,0,140,0,225,0,50,0,0,0,0,0,28,0,98,0,208,0,236,0,240,0,192,0,182,0,232,0,67,0,145,0,129,0,247,0,19,0,208,0,16,0,114,0,75,0,74,0,133,0,32,0,165,0,0,0,132,0,249,0,120,0,4,0,227,0,188,0,228,0,189,0,0,0,0,0,76,0,60,0,105,0,134,0,104,0,172,0,137,0,252,0);
signal scenario_full  : scenario_type := (0,0,196,31,120,31,24,31,203,31,203,30,214,31,158,31,92,31,13,31,144,31,139,31,154,31,46,31,47,31,150,31,231,31,231,30,168,31,29,31,29,30,139,31,245,31,105,31,105,30,105,29,28,31,234,31,103,31,103,30,103,29,171,31,179,31,179,30,118,31,33,31,188,31,188,30,188,29,239,31,239,30,128,31,2,31,6,31,213,31,127,31,127,30,99,31,99,30,218,31,118,31,246,31,246,30,28,31,72,31,213,31,197,31,170,31,78,31,78,30,223,31,102,31,174,31,174,30,63,31,135,31,158,31,81,31,199,31,8,31,8,30,183,31,141,31,141,30,141,29,90,31,42,31,42,30,207,31,132,31,210,31,210,30,167,31,250,31,152,31,239,31,192,31,91,31,91,30,179,31,18,31,158,31,216,31,22,31,75,31,2,31,138,31,138,30,138,29,188,31,118,31,173,31,33,31,216,31,210,31,164,31,45,31,65,31,65,30,193,31,84,31,93,31,215,31,208,31,62,31,40,31,40,30,234,31,199,31,199,30,86,31,86,30,120,31,120,30,120,29,93,31,240,31,164,31,167,31,167,30,227,31,71,31,244,31,120,31,56,31,56,30,235,31,235,30,255,31,250,31,49,31,41,31,181,31,181,30,66,31,238,31,110,31,73,31,73,30,247,31,145,31,149,31,4,31,202,31,99,31,139,31,164,31,173,31,173,30,16,31,151,31,4,31,178,31,241,31,127,31,129,31,230,31,239,31,175,31,175,30,47,31,47,30,169,31,10,31,83,31,83,30,140,31,72,31,13,31,13,30,48,31,48,30,23,31,23,30,77,31,131,31,131,30,224,31,82,31,164,31,255,31,252,31,3,31,3,30,163,31,218,31,218,30,11,31,245,31,216,31,232,31,116,31,8,31,47,31,42,31,124,31,193,31,37,31,37,30,64,31,7,31,1,31,240,31,57,31,223,31,215,31,215,30,12,31,125,31,202,31,202,30,202,29,108,31,68,31,184,31,219,31,45,31,146,31,223,31,225,31,225,30,225,29,225,28,69,31,106,31,103,31,216,31,216,30,209,31,48,31,153,31,153,30,192,31,149,31,188,31,67,31,85,31,204,31,250,31,185,31,147,31,116,31,242,31,242,30,165,31,103,31,215,31,5,31,5,30,141,31,253,31,154,31,164,31,14,31,9,31,222,31,222,30,129,31,142,31,142,30,142,29,180,31,180,30,201,31,13,31,240,31,40,31,252,31,26,31,122,31,245,31,139,31,128,31,128,30,128,31,139,31,64,31,253,31,81,31,216,31,216,30,18,31,199,31,81,31,107,31,46,31,46,30,23,31,23,30,154,31,201,31,95,31,120,31,148,31,26,31,51,31,51,30,36,31,21,31,14,31,14,30,218,31,14,31,201,31,201,30,144,31,144,30,196,31,104,31,104,30,231,31,216,31,179,31,96,31,63,31,41,31,87,31,87,30,60,31,239,31,197,31,253,31,92,31,249,31,103,31,205,31,101,31,30,31,184,31,184,30,73,31,98,31,14,31,42,31,254,31,129,31,248,31,199,31,30,31,249,31,17,31,189,31,188,31,188,30,188,29,168,31,168,30,168,29,55,31,185,31,67,31,73,31,101,31,101,30,242,31,94,31,94,30,94,29,46,31,55,31,133,31,32,31,235,31,111,31,7,31,156,31,199,31,245,31,73,31,253,31,253,30,253,29,207,31,115,31,209,31,53,31,23,31,15,31,15,30,73,31,156,31,114,31,66,31,41,31,102,31,8,31,8,30,66,31,230,31,151,31,199,31,199,30,54,31,69,31,69,30,108,31,170,31,146,31,83,31,207,31,205,31,230,31,252,31,252,30,210,31,31,31,165,31,153,31,243,31,243,30,20,31,243,31,243,30,77,31,122,31,68,31,68,30,68,29,15,31,227,31,68,31,250,31,22,31,145,31,145,30,61,31,104,31,220,31,241,31,98,31,98,30,98,29,98,28,98,27,98,26,153,31,153,30,199,31,125,31,84,31,174,31,236,31,208,31,245,31,129,31,129,30,149,31,65,31,82,31,83,31,179,31,123,31,192,31,14,31,14,30,199,31,85,31,144,31,233,31,111,31,90,31,90,30,46,31,93,31,49,31,12,31,225,31,239,31,125,31,171,31,214,31,82,31,137,31,30,31,204,31,204,30,15,31,182,31,51,31,25,31,129,31,182,31,135,31,163,31,163,30,20,31,130,31,117,31,39,31,119,31,198,31,153,31,34,31,235,31,6,31,6,30,36,31,36,30,70,31,159,31,215,31,215,30,19,31,19,30,187,31,2,31,2,30,99,31,176,31,91,31,91,30,91,29,255,31,172,31,172,30,181,31,207,31,191,31,206,31,95,31,185,31,1,31,10,31,245,31,108,31,231,31,255,31,177,31,132,31,117,31,105,31,242,31,216,31,216,30,216,29,216,28,216,27,204,31,136,31,242,31,241,31,165,31,198,31,198,30,144,31,143,31,149,31,84,31,73,31,250,31,51,31,134,31,139,31,205,31,206,31,253,31,253,30,233,31,7,31,7,30,7,29,174,31,174,30,174,29,248,31,212,31,100,31,30,31,146,31,146,30,146,29,235,31,23,31,52,31,8,31,8,30,8,29,74,31,210,31,162,31,206,31,175,31,203,31,110,31,124,31,124,30,155,31,223,31,225,31,141,31,105,31,227,31,142,31,177,31,220,31,197,31,177,31,177,30,128,31,77,31,77,30,127,31,127,30,127,29,39,31,151,31,88,31,98,31,98,30,191,31,191,30,14,31,23,31,250,31,250,30,250,29,120,31,120,30,120,29,220,31,154,31,154,30,249,31,234,31,179,31,180,31,104,31,104,30,104,29,13,31,124,31,135,31,48,31,78,31,78,30,78,29,72,31,242,31,150,31,158,31,193,31,182,31,182,30,191,31,191,30,98,31,2,31,130,31,70,31,177,31,238,31,111,31,140,31,89,31,91,31,91,30,162,31,90,31,90,30,90,29,169,31,120,31,37,31,133,31,153,31,142,31,241,31,37,31,232,31,28,31,245,31,147,31,54,31,245,31,207,31,192,31,221,31,55,31,129,31,118,31,221,31,83,31,99,31,99,30,49,31,142,31,241,31,95,31,145,31,75,31,137,31,173,31,173,30,223,31,181,31,208,31,118,31,195,31,41,31,202,31,152,31,137,31,80,31,67,31,34,31,129,31,3,31,11,31,255,31,57,31,85,31,85,30,124,31,157,31,157,30,145,31,7,31,174,31,145,31,129,31,216,31,172,31,60,31,227,31,227,30,216,31,173,31,49,31,207,31,140,31,225,31,50,31,50,30,50,29,28,31,98,31,208,31,236,31,240,31,192,31,182,31,232,31,67,31,145,31,129,31,247,31,19,31,208,31,16,31,114,31,75,31,74,31,133,31,32,31,165,31,165,30,132,31,249,31,120,31,4,31,227,31,188,31,228,31,189,31,189,30,189,29,76,31,60,31,105,31,134,31,104,31,172,31,137,31,252,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
