-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_380 is
end project_tb_380;

architecture project_tb_arch_380 of project_tb_380 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 711;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (87,0,189,0,77,0,160,0,217,0,16,0,179,0,86,0,246,0,77,0,0,0,227,0,0,0,158,0,6,0,0,0,199,0,67,0,222,0,0,0,0,0,78,0,156,0,207,0,137,0,0,0,96,0,173,0,0,0,112,0,81,0,0,0,148,0,103,0,0,0,136,0,12,0,41,0,169,0,48,0,242,0,231,0,23,0,0,0,165,0,0,0,113,0,146,0,0,0,180,0,135,0,243,0,88,0,244,0,32,0,0,0,22,0,252,0,169,0,217,0,239,0,0,0,0,0,229,0,132,0,229,0,230,0,208,0,192,0,4,0,39,0,0,0,0,0,77,0,6,0,231,0,0,0,6,0,86,0,10,0,13,0,182,0,61,0,239,0,210,0,42,0,117,0,217,0,58,0,92,0,7,0,0,0,212,0,4,0,96,0,38,0,0,0,46,0,12,0,0,0,206,0,180,0,171,0,175,0,250,0,190,0,92,0,3,0,211,0,79,0,0,0,212,0,193,0,201,0,222,0,74,0,227,0,0,0,247,0,11,0,242,0,4,0,101,0,0,0,88,0,0,0,237,0,10,0,97,0,241,0,129,0,76,0,192,0,231,0,235,0,253,0,12,0,249,0,245,0,0,0,139,0,165,0,186,0,0,0,0,0,134,0,180,0,0,0,0,0,88,0,25,0,189,0,237,0,0,0,169,0,65,0,142,0,5,0,0,0,0,0,56,0,0,0,0,0,35,0,184,0,248,0,0,0,0,0,253,0,134,0,0,0,222,0,210,0,64,0,43,0,0,0,162,0,177,0,3,0,153,0,196,0,118,0,0,0,174,0,189,0,125,0,90,0,175,0,189,0,73,0,91,0,223,0,58,0,0,0,136,0,0,0,157,0,101,0,56,0,0,0,123,0,177,0,230,0,6,0,0,0,149,0,0,0,104,0,249,0,70,0,242,0,244,0,207,0,176,0,210,0,197,0,46,0,104,0,44,0,131,0,155,0,75,0,0,0,110,0,137,0,192,0,253,0,181,0,108,0,0,0,91,0,113,0,164,0,0,0,0,0,116,0,139,0,0,0,45,0,105,0,196,0,204,0,41,0,0,0,102,0,0,0,156,0,112,0,29,0,0,0,3,0,178,0,0,0,0,0,200,0,18,0,214,0,24,0,0,0,195,0,191,0,140,0,143,0,42,0,154,0,0,0,0,0,95,0,243,0,11,0,61,0,224,0,34,0,249,0,230,0,75,0,0,0,236,0,0,0,11,0,81,0,161,0,230,0,0,0,121,0,154,0,62,0,0,0,201,0,132,0,92,0,97,0,0,0,133,0,127,0,114,0,0,0,107,0,190,0,117,0,94,0,40,0,6,0,1,0,63,0,7,0,141,0,56,0,187,0,42,0,93,0,8,0,90,0,0,0,155,0,49,0,51,0,242,0,5,0,0,0,168,0,0,0,208,0,113,0,147,0,0,0,255,0,121,0,38,0,169,0,168,0,158,0,0,0,157,0,92,0,11,0,202,0,106,0,222,0,27,0,236,0,42,0,72,0,0,0,127,0,103,0,51,0,62,0,88,0,175,0,72,0,153,0,0,0,0,0,59,0,92,0,91,0,64,0,201,0,80,0,209,0,193,0,148,0,0,0,192,0,104,0,87,0,153,0,103,0,151,0,0,0,16,0,191,0,157,0,82,0,115,0,182,0,0,0,166,0,0,0,71,0,168,0,3,0,42,0,0,0,239,0,80,0,0,0,255,0,224,0,64,0,153,0,113,0,218,0,141,0,110,0,0,0,39,0,0,0,28,0,0,0,209,0,23,0,0,0,234,0,105,0,84,0,62,0,189,0,40,0,0,0,120,0,150,0,0,0,212,0,131,0,2,0,177,0,0,0,151,0,0,0,176,0,195,0,152,0,166,0,133,0,201,0,0,0,240,0,155,0,46,0,0,0,19,0,234,0,26,0,200,0,44,0,104,0,0,0,129,0,28,0,41,0,167,0,0,0,0,0,0,0,41,0,226,0,29,0,151,0,163,0,48,0,38,0,67,0,0,0,0,0,134,0,0,0,0,0,178,0,141,0,67,0,0,0,0,0,230,0,49,0,62,0,11,0,31,0,244,0,0,0,0,0,187,0,34,0,0,0,0,0,0,0,216,0,177,0,0,0,116,0,199,0,101,0,125,0,237,0,8,0,59,0,15,0,174,0,207,0,0,0,206,0,78,0,0,0,86,0,153,0,100,0,133,0,80,0,67,0,118,0,49,0,157,0,35,0,113,0,68,0,0,0,118,0,0,0,97,0,131,0,59,0,42,0,0,0,70,0,54,0,0,0,47,0,187,0,95,0,64,0,43,0,180,0,0,0,92,0,168,0,0,0,155,0,221,0,0,0,160,0,165,0,39,0,0,0,64,0,165,0,232,0,20,0,27,0,77,0,98,0,28,0,174,0,55,0,0,0,49,0,10,0,145,0,140,0,113,0,117,0,169,0,56,0,79,0,0,0,38,0,17,0,175,0,0,0,16,0,30,0,179,0,199,0,97,0,181,0,246,0,146,0,158,0,176,0,0,0,0,0,75,0,239,0,187,0,243,0,59,0,0,0,0,0,81,0,15,0,119,0,194,0,129,0,28,0,234,0,0,0,51,0,192,0,89,0,178,0,0,0,206,0,173,0,184,0,253,0,127,0,241,0,243,0,65,0,175,0,131,0,51,0,193,0,0,0,0,0,2,0,209,0,6,0,84,0,0,0,0,0,8,0,48,0,78,0,19,0,37,0,237,0,42,0,9,0,126,0,40,0,250,0,181,0,208,0,224,0,222,0,64,0,20,0,184,0,173,0,38,0,105,0,179,0,44,0,215,0,0,0,153,0,239,0,186,0,28,0,0,0,223,0,0,0,135,0,35,0,85,0,167,0,252,0,17,0,9,0,169,0,126,0,47,0,0,0,103,0,203,0,205,0,108,0,143,0,0,0,209,0,117,0,35,0,210,0,85,0,0,0,168,0,161,0,69,0,240,0,244,0,54,0,174,0,0,0,234,0,214,0,135,0,188,0,5,0,17,0,40,0,106,0,0,0,232,0,0,0,167,0,77,0,192,0,167,0,193,0,243,0,0,0,168,0,111,0,0,0,129,0,4,0,174,0,0,0,211,0,219,0,203,0,204,0,0,0,0,0,130,0,144,0,141,0,0,0,68,0,20,0);
signal scenario_full  : scenario_type := (87,31,189,31,77,31,160,31,217,31,16,31,179,31,86,31,246,31,77,31,77,30,227,31,227,30,158,31,6,31,6,30,199,31,67,31,222,31,222,30,222,29,78,31,156,31,207,31,137,31,137,30,96,31,173,31,173,30,112,31,81,31,81,30,148,31,103,31,103,30,136,31,12,31,41,31,169,31,48,31,242,31,231,31,23,31,23,30,165,31,165,30,113,31,146,31,146,30,180,31,135,31,243,31,88,31,244,31,32,31,32,30,22,31,252,31,169,31,217,31,239,31,239,30,239,29,229,31,132,31,229,31,230,31,208,31,192,31,4,31,39,31,39,30,39,29,77,31,6,31,231,31,231,30,6,31,86,31,10,31,13,31,182,31,61,31,239,31,210,31,42,31,117,31,217,31,58,31,92,31,7,31,7,30,212,31,4,31,96,31,38,31,38,30,46,31,12,31,12,30,206,31,180,31,171,31,175,31,250,31,190,31,92,31,3,31,211,31,79,31,79,30,212,31,193,31,201,31,222,31,74,31,227,31,227,30,247,31,11,31,242,31,4,31,101,31,101,30,88,31,88,30,237,31,10,31,97,31,241,31,129,31,76,31,192,31,231,31,235,31,253,31,12,31,249,31,245,31,245,30,139,31,165,31,186,31,186,30,186,29,134,31,180,31,180,30,180,29,88,31,25,31,189,31,237,31,237,30,169,31,65,31,142,31,5,31,5,30,5,29,56,31,56,30,56,29,35,31,184,31,248,31,248,30,248,29,253,31,134,31,134,30,222,31,210,31,64,31,43,31,43,30,162,31,177,31,3,31,153,31,196,31,118,31,118,30,174,31,189,31,125,31,90,31,175,31,189,31,73,31,91,31,223,31,58,31,58,30,136,31,136,30,157,31,101,31,56,31,56,30,123,31,177,31,230,31,6,31,6,30,149,31,149,30,104,31,249,31,70,31,242,31,244,31,207,31,176,31,210,31,197,31,46,31,104,31,44,31,131,31,155,31,75,31,75,30,110,31,137,31,192,31,253,31,181,31,108,31,108,30,91,31,113,31,164,31,164,30,164,29,116,31,139,31,139,30,45,31,105,31,196,31,204,31,41,31,41,30,102,31,102,30,156,31,112,31,29,31,29,30,3,31,178,31,178,30,178,29,200,31,18,31,214,31,24,31,24,30,195,31,191,31,140,31,143,31,42,31,154,31,154,30,154,29,95,31,243,31,11,31,61,31,224,31,34,31,249,31,230,31,75,31,75,30,236,31,236,30,11,31,81,31,161,31,230,31,230,30,121,31,154,31,62,31,62,30,201,31,132,31,92,31,97,31,97,30,133,31,127,31,114,31,114,30,107,31,190,31,117,31,94,31,40,31,6,31,1,31,63,31,7,31,141,31,56,31,187,31,42,31,93,31,8,31,90,31,90,30,155,31,49,31,51,31,242,31,5,31,5,30,168,31,168,30,208,31,113,31,147,31,147,30,255,31,121,31,38,31,169,31,168,31,158,31,158,30,157,31,92,31,11,31,202,31,106,31,222,31,27,31,236,31,42,31,72,31,72,30,127,31,103,31,51,31,62,31,88,31,175,31,72,31,153,31,153,30,153,29,59,31,92,31,91,31,64,31,201,31,80,31,209,31,193,31,148,31,148,30,192,31,104,31,87,31,153,31,103,31,151,31,151,30,16,31,191,31,157,31,82,31,115,31,182,31,182,30,166,31,166,30,71,31,168,31,3,31,42,31,42,30,239,31,80,31,80,30,255,31,224,31,64,31,153,31,113,31,218,31,141,31,110,31,110,30,39,31,39,30,28,31,28,30,209,31,23,31,23,30,234,31,105,31,84,31,62,31,189,31,40,31,40,30,120,31,150,31,150,30,212,31,131,31,2,31,177,31,177,30,151,31,151,30,176,31,195,31,152,31,166,31,133,31,201,31,201,30,240,31,155,31,46,31,46,30,19,31,234,31,26,31,200,31,44,31,104,31,104,30,129,31,28,31,41,31,167,31,167,30,167,29,167,28,41,31,226,31,29,31,151,31,163,31,48,31,38,31,67,31,67,30,67,29,134,31,134,30,134,29,178,31,141,31,67,31,67,30,67,29,230,31,49,31,62,31,11,31,31,31,244,31,244,30,244,29,187,31,34,31,34,30,34,29,34,28,216,31,177,31,177,30,116,31,199,31,101,31,125,31,237,31,8,31,59,31,15,31,174,31,207,31,207,30,206,31,78,31,78,30,86,31,153,31,100,31,133,31,80,31,67,31,118,31,49,31,157,31,35,31,113,31,68,31,68,30,118,31,118,30,97,31,131,31,59,31,42,31,42,30,70,31,54,31,54,30,47,31,187,31,95,31,64,31,43,31,180,31,180,30,92,31,168,31,168,30,155,31,221,31,221,30,160,31,165,31,39,31,39,30,64,31,165,31,232,31,20,31,27,31,77,31,98,31,28,31,174,31,55,31,55,30,49,31,10,31,145,31,140,31,113,31,117,31,169,31,56,31,79,31,79,30,38,31,17,31,175,31,175,30,16,31,30,31,179,31,199,31,97,31,181,31,246,31,146,31,158,31,176,31,176,30,176,29,75,31,239,31,187,31,243,31,59,31,59,30,59,29,81,31,15,31,119,31,194,31,129,31,28,31,234,31,234,30,51,31,192,31,89,31,178,31,178,30,206,31,173,31,184,31,253,31,127,31,241,31,243,31,65,31,175,31,131,31,51,31,193,31,193,30,193,29,2,31,209,31,6,31,84,31,84,30,84,29,8,31,48,31,78,31,19,31,37,31,237,31,42,31,9,31,126,31,40,31,250,31,181,31,208,31,224,31,222,31,64,31,20,31,184,31,173,31,38,31,105,31,179,31,44,31,215,31,215,30,153,31,239,31,186,31,28,31,28,30,223,31,223,30,135,31,35,31,85,31,167,31,252,31,17,31,9,31,169,31,126,31,47,31,47,30,103,31,203,31,205,31,108,31,143,31,143,30,209,31,117,31,35,31,210,31,85,31,85,30,168,31,161,31,69,31,240,31,244,31,54,31,174,31,174,30,234,31,214,31,135,31,188,31,5,31,17,31,40,31,106,31,106,30,232,31,232,30,167,31,77,31,192,31,167,31,193,31,243,31,243,30,168,31,111,31,111,30,129,31,4,31,174,31,174,30,211,31,219,31,203,31,204,31,204,30,204,29,130,31,144,31,141,31,141,30,68,31,20,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
