-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 974;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,187,0,0,0,205,0,195,0,140,0,22,0,52,0,196,0,207,0,222,0,182,0,90,0,0,0,78,0,193,0,225,0,39,0,226,0,162,0,0,0,0,0,77,0,66,0,56,0,159,0,75,0,116,0,126,0,135,0,120,0,227,0,0,0,100,0,0,0,32,0,9,0,53,0,190,0,97,0,157,0,40,0,195,0,19,0,39,0,133,0,90,0,0,0,207,0,60,0,251,0,115,0,172,0,199,0,66,0,190,0,0,0,109,0,200,0,98,0,0,0,231,0,204,0,240,0,181,0,213,0,60,0,24,0,92,0,0,0,82,0,53,0,0,0,0,0,0,0,167,0,60,0,177,0,0,0,197,0,32,0,112,0,49,0,132,0,137,0,8,0,70,0,35,0,215,0,164,0,67,0,179,0,59,0,54,0,158,0,110,0,45,0,23,0,0,0,107,0,250,0,219,0,217,0,197,0,90,0,103,0,179,0,129,0,108,0,178,0,170,0,121,0,193,0,93,0,128,0,219,0,0,0,127,0,105,0,185,0,131,0,80,0,248,0,85,0,177,0,137,0,110,0,78,0,138,0,0,0,107,0,186,0,175,0,1,0,168,0,114,0,66,0,19,0,248,0,0,0,249,0,146,0,68,0,30,0,120,0,246,0,82,0,0,0,105,0,15,0,142,0,0,0,32,0,132,0,34,0,203,0,0,0,130,0,216,0,88,0,225,0,131,0,55,0,132,0,0,0,0,0,225,0,54,0,225,0,58,0,234,0,216,0,144,0,197,0,0,0,50,0,123,0,0,0,10,0,0,0,0,0,0,0,202,0,0,0,71,0,0,0,205,0,80,0,136,0,0,0,39,0,0,0,0,0,190,0,0,0,216,0,244,0,23,0,241,0,184,0,227,0,0,0,12,0,20,0,0,0,91,0,230,0,33,0,170,0,79,0,0,0,9,0,193,0,152,0,0,0,101,0,0,0,186,0,90,0,212,0,191,0,83,0,8,0,0,0,97,0,176,0,204,0,0,0,173,0,243,0,197,0,83,0,0,0,195,0,182,0,0,0,163,0,0,0,225,0,207,0,51,0,11,0,17,0,103,0,95,0,233,0,0,0,232,0,137,0,60,0,43,0,0,0,0,0,192,0,0,0,49,0,226,0,240,0,255,0,248,0,115,0,232,0,32,0,210,0,214,0,47,0,47,0,149,0,27,0,73,0,128,0,24,0,0,0,252,0,209,0,0,0,116,0,0,0,178,0,0,0,205,0,113,0,0,0,241,0,98,0,219,0,227,0,194,0,131,0,117,0,0,0,127,0,128,0,0,0,50,0,44,0,201,0,176,0,0,0,0,0,153,0,117,0,133,0,144,0,237,0,23,0,14,0,143,0,235,0,53,0,27,0,0,0,208,0,239,0,49,0,0,0,64,0,44,0,219,0,206,0,18,0,2,0,24,0,0,0,100,0,167,0,176,0,0,0,215,0,78,0,0,0,0,0,85,0,25,0,24,0,36,0,88,0,17,0,134,0,47,0,0,0,252,0,217,0,73,0,175,0,58,0,0,0,90,0,39,0,186,0,0,0,3,0,0,0,117,0,0,0,101,0,150,0,192,0,169,0,3,0,151,0,11,0,5,0,251,0,19,0,0,0,83,0,63,0,153,0,188,0,110,0,198,0,0,0,107,0,239,0,20,0,209,0,0,0,93,0,190,0,0,0,34,0,66,0,231,0,210,0,125,0,0,0,97,0,89,0,132,0,170,0,30,0,83,0,11,0,172,0,168,0,17,0,77,0,117,0,180,0,174,0,24,0,206,0,164,0,233,0,232,0,219,0,225,0,198,0,219,0,183,0,69,0,0,0,0,0,88,0,241,0,101,0,235,0,226,0,0,0,90,0,146,0,68,0,205,0,0,0,0,0,18,0,21,0,201,0,175,0,211,0,0,0,40,0,70,0,21,0,2,0,59,0,198,0,29,0,92,0,0,0,207,0,48,0,39,0,62,0,167,0,160,0,0,0,88,0,0,0,195,0,184,0,91,0,95,0,128,0,158,0,155,0,0,0,0,0,0,0,35,0,0,0,208,0,117,0,0,0,22,0,171,0,93,0,94,0,218,0,228,0,0,0,13,0,73,0,221,0,0,0,215,0,180,0,145,0,102,0,44,0,33,0,0,0,29,0,200,0,172,0,187,0,109,0,0,0,187,0,0,0,143,0,89,0,241,0,232,0,116,0,116,0,210,0,144,0,74,0,217,0,130,0,0,0,31,0,55,0,240,0,186,0,3,0,246,0,0,0,55,0,65,0,187,0,0,0,162,0,68,0,0,0,15,0,18,0,136,0,137,0,239,0,182,0,165,0,112,0,80,0,0,0,0,0,99,0,106,0,44,0,45,0,142,0,10,0,117,0,198,0,44,0,66,0,0,0,59,0,116,0,164,0,254,0,246,0,0,0,171,0,0,0,0,0,87,0,0,0,131,0,222,0,0,0,88,0,13,0,126,0,114,0,58,0,45,0,237,0,139,0,0,0,33,0,100,0,16,0,128,0,3,0,146,0,255,0,47,0,0,0,232,0,31,0,169,0,95,0,102,0,235,0,24,0,139,0,230,0,169,0,154,0,222,0,224,0,0,0,93,0,103,0,182,0,117,0,62,0,77,0,254,0,33,0,121,0,0,0,178,0,62,0,0,0,0,0,188,0,0,0,226,0,225,0,0,0,197,0,149,0,72,0,156,0,126,0,194,0,0,0,31,0,16,0,0,0,236,0,185,0,63,0,200,0,153,0,57,0,153,0,1,0,11,0,180,0,255,0,0,0,0,0,0,0,41,0,147,0,96,0,0,0,0,0,0,0,106,0,104,0,97,0,75,0,203,0,89,0,0,0,109,0,0,0,133,0,13,0,219,0,25,0,203,0,250,0,9,0,167,0,93,0,76,0,152,0,191,0,154,0,111,0,184,0,100,0,0,0,0,0,0,0,198,0,78,0,37,0,207,0,0,0,75,0,237,0,208,0,2,0,182,0,118,0,193,0,72,0,0,0,34,0,153,0,71,0,0,0,0,0,40,0,9,0,162,0,77,0,9,0,222,0,210,0,153,0,131,0,73,0,126,0,53,0,107,0,242,0,0,0,127,0,182,0,246,0,198,0,144,0,75,0,180,0,43,0,137,0,72,0,0,0,233,0,230,0,11,0,0,0,0,0,41,0,3,0,27,0,237,0,19,0,3,0,0,0,152,0,90,0,112,0,120,0,100,0,70,0,168,0,80,0,0,0,218,0,128,0,156,0,42,0,209,0,34,0,0,0,71,0,0,0,43,0,127,0,10,0,199,0,22,0,10,0,0,0,27,0,129,0,167,0,36,0,1,0,204,0,47,0,68,0,51,0,0,0,110,0,213,0,97,0,145,0,152,0,144,0,34,0,195,0,0,0,233,0,224,0,0,0,0,0,219,0,6,0,0,0,0,0,0,0,155,0,0,0,105,0,204,0,39,0,93,0,65,0,32,0,203,0,88,0,0,0,251,0,185,0,179,0,197,0,101,0,71,0,0,0,206,0,27,0,198,0,222,0,39,0,146,0,75,0,122,0,0,0,0,0,135,0,21,0,100,0,162,0,0,0,247,0,49,0,77,0,171,0,0,0,0,0,201,0,243,0,0,0,199,0,39,0,77,0,201,0,163,0,149,0,33,0,164,0,159,0,4,0,47,0,208,0,199,0,222,0,63,0,164,0,53,0,158,0,89,0,31,0,166,0,0,0,52,0,217,0,157,0,171,0,79,0,174,0,97,0,0,0,211,0,0,0,18,0,129,0,156,0,169,0,183,0,0,0,26,0,0,0,250,0,185,0,17,0,70,0,0,0,28,0,100,0,62,0,179,0,181,0,122,0,196,0,116,0,0,0,0,0,108,0,202,0,152,0,51,0,252,0,75,0,142,0,0,0,140,0,219,0,185,0,162,0,75,0,208,0,60,0,55,0,0,0,107,0,228,0,72,0,60,0,215,0,11,0,0,0,138,0,0,0,37,0,52,0,221,0,226,0,49,0,0,0,66,0,0,0,101,0,6,0,191,0,159,0,0,0,1,0,17,0,149,0,236,0,108,0,23,0,96,0,179,0,62,0,90,0,0,0,144,0,162,0,0,0,0,0,0,0,24,0,34,0,128,0,29,0,0,0,0,0,0,0,0,0,0,0,9,0,0,0,78,0,51,0,0,0,0,0,213,0,192,0,161,0,193,0,39,0,237,0,0,0,77,0,174,0,23,0,40,0,46,0,39,0,254,0,109,0,80,0,62,0,0,0,125,0,0,0,161,0,222,0,0,0,105,0,73,0,85,0,46,0,248,0,62,0,92,0,141,0,94,0,0,0,82,0);
signal scenario_full  : scenario_type := (0,0,0,0,187,31,187,30,205,31,195,31,140,31,22,31,52,31,196,31,207,31,222,31,182,31,90,31,90,30,78,31,193,31,225,31,39,31,226,31,162,31,162,30,162,29,77,31,66,31,56,31,159,31,75,31,116,31,126,31,135,31,120,31,227,31,227,30,100,31,100,30,32,31,9,31,53,31,190,31,97,31,157,31,40,31,195,31,19,31,39,31,133,31,90,31,90,30,207,31,60,31,251,31,115,31,172,31,199,31,66,31,190,31,190,30,109,31,200,31,98,31,98,30,231,31,204,31,240,31,181,31,213,31,60,31,24,31,92,31,92,30,82,31,53,31,53,30,53,29,53,28,167,31,60,31,177,31,177,30,197,31,32,31,112,31,49,31,132,31,137,31,8,31,70,31,35,31,215,31,164,31,67,31,179,31,59,31,54,31,158,31,110,31,45,31,23,31,23,30,107,31,250,31,219,31,217,31,197,31,90,31,103,31,179,31,129,31,108,31,178,31,170,31,121,31,193,31,93,31,128,31,219,31,219,30,127,31,105,31,185,31,131,31,80,31,248,31,85,31,177,31,137,31,110,31,78,31,138,31,138,30,107,31,186,31,175,31,1,31,168,31,114,31,66,31,19,31,248,31,248,30,249,31,146,31,68,31,30,31,120,31,246,31,82,31,82,30,105,31,15,31,142,31,142,30,32,31,132,31,34,31,203,31,203,30,130,31,216,31,88,31,225,31,131,31,55,31,132,31,132,30,132,29,225,31,54,31,225,31,58,31,234,31,216,31,144,31,197,31,197,30,50,31,123,31,123,30,10,31,10,30,10,29,10,28,202,31,202,30,71,31,71,30,205,31,80,31,136,31,136,30,39,31,39,30,39,29,190,31,190,30,216,31,244,31,23,31,241,31,184,31,227,31,227,30,12,31,20,31,20,30,91,31,230,31,33,31,170,31,79,31,79,30,9,31,193,31,152,31,152,30,101,31,101,30,186,31,90,31,212,31,191,31,83,31,8,31,8,30,97,31,176,31,204,31,204,30,173,31,243,31,197,31,83,31,83,30,195,31,182,31,182,30,163,31,163,30,225,31,207,31,51,31,11,31,17,31,103,31,95,31,233,31,233,30,232,31,137,31,60,31,43,31,43,30,43,29,192,31,192,30,49,31,226,31,240,31,255,31,248,31,115,31,232,31,32,31,210,31,214,31,47,31,47,31,149,31,27,31,73,31,128,31,24,31,24,30,252,31,209,31,209,30,116,31,116,30,178,31,178,30,205,31,113,31,113,30,241,31,98,31,219,31,227,31,194,31,131,31,117,31,117,30,127,31,128,31,128,30,50,31,44,31,201,31,176,31,176,30,176,29,153,31,117,31,133,31,144,31,237,31,23,31,14,31,143,31,235,31,53,31,27,31,27,30,208,31,239,31,49,31,49,30,64,31,44,31,219,31,206,31,18,31,2,31,24,31,24,30,100,31,167,31,176,31,176,30,215,31,78,31,78,30,78,29,85,31,25,31,24,31,36,31,88,31,17,31,134,31,47,31,47,30,252,31,217,31,73,31,175,31,58,31,58,30,90,31,39,31,186,31,186,30,3,31,3,30,117,31,117,30,101,31,150,31,192,31,169,31,3,31,151,31,11,31,5,31,251,31,19,31,19,30,83,31,63,31,153,31,188,31,110,31,198,31,198,30,107,31,239,31,20,31,209,31,209,30,93,31,190,31,190,30,34,31,66,31,231,31,210,31,125,31,125,30,97,31,89,31,132,31,170,31,30,31,83,31,11,31,172,31,168,31,17,31,77,31,117,31,180,31,174,31,24,31,206,31,164,31,233,31,232,31,219,31,225,31,198,31,219,31,183,31,69,31,69,30,69,29,88,31,241,31,101,31,235,31,226,31,226,30,90,31,146,31,68,31,205,31,205,30,205,29,18,31,21,31,201,31,175,31,211,31,211,30,40,31,70,31,21,31,2,31,59,31,198,31,29,31,92,31,92,30,207,31,48,31,39,31,62,31,167,31,160,31,160,30,88,31,88,30,195,31,184,31,91,31,95,31,128,31,158,31,155,31,155,30,155,29,155,28,35,31,35,30,208,31,117,31,117,30,22,31,171,31,93,31,94,31,218,31,228,31,228,30,13,31,73,31,221,31,221,30,215,31,180,31,145,31,102,31,44,31,33,31,33,30,29,31,200,31,172,31,187,31,109,31,109,30,187,31,187,30,143,31,89,31,241,31,232,31,116,31,116,31,210,31,144,31,74,31,217,31,130,31,130,30,31,31,55,31,240,31,186,31,3,31,246,31,246,30,55,31,65,31,187,31,187,30,162,31,68,31,68,30,15,31,18,31,136,31,137,31,239,31,182,31,165,31,112,31,80,31,80,30,80,29,99,31,106,31,44,31,45,31,142,31,10,31,117,31,198,31,44,31,66,31,66,30,59,31,116,31,164,31,254,31,246,31,246,30,171,31,171,30,171,29,87,31,87,30,131,31,222,31,222,30,88,31,13,31,126,31,114,31,58,31,45,31,237,31,139,31,139,30,33,31,100,31,16,31,128,31,3,31,146,31,255,31,47,31,47,30,232,31,31,31,169,31,95,31,102,31,235,31,24,31,139,31,230,31,169,31,154,31,222,31,224,31,224,30,93,31,103,31,182,31,117,31,62,31,77,31,254,31,33,31,121,31,121,30,178,31,62,31,62,30,62,29,188,31,188,30,226,31,225,31,225,30,197,31,149,31,72,31,156,31,126,31,194,31,194,30,31,31,16,31,16,30,236,31,185,31,63,31,200,31,153,31,57,31,153,31,1,31,11,31,180,31,255,31,255,30,255,29,255,28,41,31,147,31,96,31,96,30,96,29,96,28,106,31,104,31,97,31,75,31,203,31,89,31,89,30,109,31,109,30,133,31,13,31,219,31,25,31,203,31,250,31,9,31,167,31,93,31,76,31,152,31,191,31,154,31,111,31,184,31,100,31,100,30,100,29,100,28,198,31,78,31,37,31,207,31,207,30,75,31,237,31,208,31,2,31,182,31,118,31,193,31,72,31,72,30,34,31,153,31,71,31,71,30,71,29,40,31,9,31,162,31,77,31,9,31,222,31,210,31,153,31,131,31,73,31,126,31,53,31,107,31,242,31,242,30,127,31,182,31,246,31,198,31,144,31,75,31,180,31,43,31,137,31,72,31,72,30,233,31,230,31,11,31,11,30,11,29,41,31,3,31,27,31,237,31,19,31,3,31,3,30,152,31,90,31,112,31,120,31,100,31,70,31,168,31,80,31,80,30,218,31,128,31,156,31,42,31,209,31,34,31,34,30,71,31,71,30,43,31,127,31,10,31,199,31,22,31,10,31,10,30,27,31,129,31,167,31,36,31,1,31,204,31,47,31,68,31,51,31,51,30,110,31,213,31,97,31,145,31,152,31,144,31,34,31,195,31,195,30,233,31,224,31,224,30,224,29,219,31,6,31,6,30,6,29,6,28,155,31,155,30,105,31,204,31,39,31,93,31,65,31,32,31,203,31,88,31,88,30,251,31,185,31,179,31,197,31,101,31,71,31,71,30,206,31,27,31,198,31,222,31,39,31,146,31,75,31,122,31,122,30,122,29,135,31,21,31,100,31,162,31,162,30,247,31,49,31,77,31,171,31,171,30,171,29,201,31,243,31,243,30,199,31,39,31,77,31,201,31,163,31,149,31,33,31,164,31,159,31,4,31,47,31,208,31,199,31,222,31,63,31,164,31,53,31,158,31,89,31,31,31,166,31,166,30,52,31,217,31,157,31,171,31,79,31,174,31,97,31,97,30,211,31,211,30,18,31,129,31,156,31,169,31,183,31,183,30,26,31,26,30,250,31,185,31,17,31,70,31,70,30,28,31,100,31,62,31,179,31,181,31,122,31,196,31,116,31,116,30,116,29,108,31,202,31,152,31,51,31,252,31,75,31,142,31,142,30,140,31,219,31,185,31,162,31,75,31,208,31,60,31,55,31,55,30,107,31,228,31,72,31,60,31,215,31,11,31,11,30,138,31,138,30,37,31,52,31,221,31,226,31,49,31,49,30,66,31,66,30,101,31,6,31,191,31,159,31,159,30,1,31,17,31,149,31,236,31,108,31,23,31,96,31,179,31,62,31,90,31,90,30,144,31,162,31,162,30,162,29,162,28,24,31,34,31,128,31,29,31,29,30,29,29,29,28,29,27,29,26,9,31,9,30,78,31,51,31,51,30,51,29,213,31,192,31,161,31,193,31,39,31,237,31,237,30,77,31,174,31,23,31,40,31,46,31,39,31,254,31,109,31,80,31,62,31,62,30,125,31,125,30,161,31,222,31,222,30,105,31,73,31,85,31,46,31,248,31,62,31,92,31,141,31,94,31,94,30,82,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
