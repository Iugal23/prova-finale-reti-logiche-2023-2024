-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_799 is
end project_tb_799;

architecture project_tb_arch_799 of project_tb_799 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 759;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (71,0,38,0,1,0,1,0,216,0,131,0,58,0,0,0,153,0,76,0,225,0,0,0,147,0,173,0,0,0,0,0,89,0,111,0,224,0,70,0,60,0,221,0,0,0,34,0,0,0,36,0,182,0,218,0,216,0,169,0,87,0,41,0,238,0,0,0,61,0,0,0,72,0,174,0,15,0,113,0,59,0,225,0,143,0,170,0,146,0,107,0,0,0,201,0,213,0,144,0,0,0,243,0,92,0,87,0,96,0,241,0,43,0,0,0,0,0,0,0,208,0,230,0,200,0,226,0,27,0,0,0,51,0,0,0,0,0,47,0,0,0,136,0,75,0,33,0,103,0,75,0,193,0,66,0,12,0,0,0,223,0,247,0,0,0,0,0,88,0,191,0,79,0,144,0,153,0,0,0,191,0,0,0,0,0,176,0,72,0,0,0,172,0,50,0,0,0,0,0,20,0,0,0,227,0,0,0,0,0,203,0,26,0,193,0,207,0,160,0,0,0,163,0,151,0,24,0,199,0,217,0,203,0,0,0,182,0,61,0,104,0,180,0,86,0,41,0,57,0,234,0,0,0,39,0,185,0,157,0,110,0,26,0,107,0,94,0,76,0,26,0,18,0,235,0,207,0,58,0,150,0,189,0,0,0,0,0,0,0,98,0,7,0,213,0,0,0,0,0,225,0,252,0,158,0,135,0,118,0,96,0,143,0,50,0,21,0,159,0,245,0,215,0,199,0,142,0,0,0,99,0,78,0,91,0,103,0,48,0,106,0,0,0,0,0,34,0,0,0,115,0,0,0,53,0,0,0,37,0,223,0,6,0,34,0,0,0,193,0,134,0,0,0,139,0,37,0,133,0,173,0,115,0,5,0,181,0,0,0,23,0,9,0,0,0,69,0,92,0,86,0,138,0,184,0,49,0,236,0,76,0,147,0,59,0,185,0,246,0,205,0,14,0,0,0,15,0,0,0,235,0,37,0,0,0,0,0,0,0,210,0,13,0,0,0,0,0,109,0,146,0,200,0,14,0,0,0,208,0,19,0,0,0,111,0,3,0,27,0,106,0,66,0,0,0,232,0,160,0,165,0,81,0,0,0,189,0,63,0,152,0,230,0,64,0,222,0,206,0,217,0,127,0,233,0,0,0,0,0,200,0,87,0,91,0,139,0,45,0,34,0,0,0,157,0,116,0,102,0,243,0,237,0,224,0,30,0,156,0,147,0,159,0,0,0,233,0,17,0,75,0,222,0,26,0,202,0,0,0,127,0,171,0,87,0,49,0,0,0,0,0,117,0,60,0,136,0,46,0,0,0,172,0,84,0,36,0,142,0,157,0,248,0,144,0,13,0,194,0,29,0,152,0,26,0,205,0,241,0,0,0,248,0,23,0,209,0,67,0,237,0,0,0,240,0,0,0,190,0,77,0,0,0,73,0,114,0,173,0,61,0,143,0,10,0,242,0,0,0,0,0,255,0,12,0,223,0,219,0,217,0,0,0,79,0,186,0,0,0,0,0,37,0,86,0,191,0,230,0,54,0,0,0,255,0,140,0,26,0,104,0,214,0,174,0,249,0,45,0,203,0,0,0,210,0,65,0,93,0,30,0,162,0,0,0,47,0,239,0,0,0,34,0,102,0,0,0,226,0,195,0,104,0,0,0,209,0,95,0,234,0,2,0,12,0,0,0,218,0,77,0,53,0,117,0,38,0,107,0,93,0,9,0,251,0,73,0,79,0,170,0,145,0,248,0,197,0,78,0,88,0,116,0,0,0,157,0,220,0,65,0,86,0,168,0,19,0,235,0,204,0,0,0,195,0,113,0,135,0,165,0,0,0,0,0,67,0,126,0,109,0,25,0,250,0,217,0,195,0,128,0,0,0,23,0,122,0,209,0,71,0,140,0,0,0,102,0,131,0,0,0,0,0,97,0,0,0,74,0,0,0,209,0,82,0,205,0,4,0,46,0,155,0,8,0,0,0,248,0,35,0,204,0,0,0,221,0,135,0,0,0,193,0,155,0,36,0,0,0,0,0,0,0,236,0,10,0,123,0,83,0,233,0,54,0,0,0,196,0,224,0,218,0,180,0,0,0,123,0,76,0,219,0,126,0,0,0,30,0,190,0,0,0,152,0,66,0,235,0,191,0,0,0,231,0,165,0,254,0,173,0,22,0,244,0,59,0,91,0,71,0,195,0,0,0,164,0,3,0,0,0,125,0,0,0,0,0,80,0,88,0,92,0,72,0,84,0,46,0,80,0,189,0,158,0,222,0,0,0,29,0,248,0,146,0,30,0,251,0,49,0,157,0,18,0,75,0,0,0,0,0,93,0,0,0,239,0,98,0,111,0,120,0,134,0,116,0,108,0,10,0,159,0,0,0,92,0,46,0,0,0,135,0,0,0,0,0,0,0,132,0,75,0,180,0,54,0,0,0,60,0,14,0,82,0,0,0,0,0,4,0,172,0,101,0,0,0,104,0,231,0,0,0,189,0,0,0,0,0,50,0,162,0,126,0,0,0,212,0,108,0,0,0,174,0,215,0,177,0,192,0,0,0,232,0,65,0,0,0,0,0,0,0,0,0,62,0,201,0,118,0,0,0,0,0,0,0,0,0,0,0,6,0,32,0,0,0,8,0,0,0,40,0,203,0,124,0,9,0,29,0,199,0,0,0,191,0,32,0,177,0,22,0,124,0,110,0,243,0,26,0,140,0,11,0,123,0,46,0,0,0,11,0,202,0,37,0,0,0,160,0,254,0,124,0,0,0,186,0,0,0,193,0,185,0,230,0,129,0,194,0,250,0,12,0,47,0,0,0,225,0,18,0,0,0,125,0,138,0,203,0,0,0,0,0,121,0,0,0,140,0,0,0,182,0,60,0,37,0,228,0,82,0,218,0,69,0,17,0,247,0,67,0,118,0,0,0,110,0,123,0,0,0,228,0,0,0,99,0,0,0,0,0,33,0,215,0,101,0,88,0,134,0,192,0,99,0,0,0,2,0,0,0,109,0,22,0,221,0,138,0,0,0,79,0,34,0,158,0,128,0,212,0,104,0,123,0,228,0,65,0,45,0,69,0,192,0,0,0,0,0,223,0,0,0,72,0,45,0,127,0,235,0,151,0,64,0,91,0,134,0,225,0,19,0,48,0,199,0,160,0,17,0,7,0,0,0,0,0,184,0,133,0,0,0,154,0,118,0,182,0,174,0,0,0,212,0,142,0,6,0,0,0,57,0,130,0,212,0,157,0,69,0,7,0,10,0,0,0,221,0,32,0,221,0,255,0,248,0,25,0,84,0,63,0,244,0,170,0,30,0,0,0,0,0,100,0,136,0,199,0,69,0,17,0,45,0,205,0,199,0,117,0,0,0,65,0,0,0,238,0,8,0,0,0,0,0,0,0,232,0,46,0,0,0,128,0);
signal scenario_full  : scenario_type := (71,31,38,31,1,31,1,31,216,31,131,31,58,31,58,30,153,31,76,31,225,31,225,30,147,31,173,31,173,30,173,29,89,31,111,31,224,31,70,31,60,31,221,31,221,30,34,31,34,30,36,31,182,31,218,31,216,31,169,31,87,31,41,31,238,31,238,30,61,31,61,30,72,31,174,31,15,31,113,31,59,31,225,31,143,31,170,31,146,31,107,31,107,30,201,31,213,31,144,31,144,30,243,31,92,31,87,31,96,31,241,31,43,31,43,30,43,29,43,28,208,31,230,31,200,31,226,31,27,31,27,30,51,31,51,30,51,29,47,31,47,30,136,31,75,31,33,31,103,31,75,31,193,31,66,31,12,31,12,30,223,31,247,31,247,30,247,29,88,31,191,31,79,31,144,31,153,31,153,30,191,31,191,30,191,29,176,31,72,31,72,30,172,31,50,31,50,30,50,29,20,31,20,30,227,31,227,30,227,29,203,31,26,31,193,31,207,31,160,31,160,30,163,31,151,31,24,31,199,31,217,31,203,31,203,30,182,31,61,31,104,31,180,31,86,31,41,31,57,31,234,31,234,30,39,31,185,31,157,31,110,31,26,31,107,31,94,31,76,31,26,31,18,31,235,31,207,31,58,31,150,31,189,31,189,30,189,29,189,28,98,31,7,31,213,31,213,30,213,29,225,31,252,31,158,31,135,31,118,31,96,31,143,31,50,31,21,31,159,31,245,31,215,31,199,31,142,31,142,30,99,31,78,31,91,31,103,31,48,31,106,31,106,30,106,29,34,31,34,30,115,31,115,30,53,31,53,30,37,31,223,31,6,31,34,31,34,30,193,31,134,31,134,30,139,31,37,31,133,31,173,31,115,31,5,31,181,31,181,30,23,31,9,31,9,30,69,31,92,31,86,31,138,31,184,31,49,31,236,31,76,31,147,31,59,31,185,31,246,31,205,31,14,31,14,30,15,31,15,30,235,31,37,31,37,30,37,29,37,28,210,31,13,31,13,30,13,29,109,31,146,31,200,31,14,31,14,30,208,31,19,31,19,30,111,31,3,31,27,31,106,31,66,31,66,30,232,31,160,31,165,31,81,31,81,30,189,31,63,31,152,31,230,31,64,31,222,31,206,31,217,31,127,31,233,31,233,30,233,29,200,31,87,31,91,31,139,31,45,31,34,31,34,30,157,31,116,31,102,31,243,31,237,31,224,31,30,31,156,31,147,31,159,31,159,30,233,31,17,31,75,31,222,31,26,31,202,31,202,30,127,31,171,31,87,31,49,31,49,30,49,29,117,31,60,31,136,31,46,31,46,30,172,31,84,31,36,31,142,31,157,31,248,31,144,31,13,31,194,31,29,31,152,31,26,31,205,31,241,31,241,30,248,31,23,31,209,31,67,31,237,31,237,30,240,31,240,30,190,31,77,31,77,30,73,31,114,31,173,31,61,31,143,31,10,31,242,31,242,30,242,29,255,31,12,31,223,31,219,31,217,31,217,30,79,31,186,31,186,30,186,29,37,31,86,31,191,31,230,31,54,31,54,30,255,31,140,31,26,31,104,31,214,31,174,31,249,31,45,31,203,31,203,30,210,31,65,31,93,31,30,31,162,31,162,30,47,31,239,31,239,30,34,31,102,31,102,30,226,31,195,31,104,31,104,30,209,31,95,31,234,31,2,31,12,31,12,30,218,31,77,31,53,31,117,31,38,31,107,31,93,31,9,31,251,31,73,31,79,31,170,31,145,31,248,31,197,31,78,31,88,31,116,31,116,30,157,31,220,31,65,31,86,31,168,31,19,31,235,31,204,31,204,30,195,31,113,31,135,31,165,31,165,30,165,29,67,31,126,31,109,31,25,31,250,31,217,31,195,31,128,31,128,30,23,31,122,31,209,31,71,31,140,31,140,30,102,31,131,31,131,30,131,29,97,31,97,30,74,31,74,30,209,31,82,31,205,31,4,31,46,31,155,31,8,31,8,30,248,31,35,31,204,31,204,30,221,31,135,31,135,30,193,31,155,31,36,31,36,30,36,29,36,28,236,31,10,31,123,31,83,31,233,31,54,31,54,30,196,31,224,31,218,31,180,31,180,30,123,31,76,31,219,31,126,31,126,30,30,31,190,31,190,30,152,31,66,31,235,31,191,31,191,30,231,31,165,31,254,31,173,31,22,31,244,31,59,31,91,31,71,31,195,31,195,30,164,31,3,31,3,30,125,31,125,30,125,29,80,31,88,31,92,31,72,31,84,31,46,31,80,31,189,31,158,31,222,31,222,30,29,31,248,31,146,31,30,31,251,31,49,31,157,31,18,31,75,31,75,30,75,29,93,31,93,30,239,31,98,31,111,31,120,31,134,31,116,31,108,31,10,31,159,31,159,30,92,31,46,31,46,30,135,31,135,30,135,29,135,28,132,31,75,31,180,31,54,31,54,30,60,31,14,31,82,31,82,30,82,29,4,31,172,31,101,31,101,30,104,31,231,31,231,30,189,31,189,30,189,29,50,31,162,31,126,31,126,30,212,31,108,31,108,30,174,31,215,31,177,31,192,31,192,30,232,31,65,31,65,30,65,29,65,28,65,27,62,31,201,31,118,31,118,30,118,29,118,28,118,27,118,26,6,31,32,31,32,30,8,31,8,30,40,31,203,31,124,31,9,31,29,31,199,31,199,30,191,31,32,31,177,31,22,31,124,31,110,31,243,31,26,31,140,31,11,31,123,31,46,31,46,30,11,31,202,31,37,31,37,30,160,31,254,31,124,31,124,30,186,31,186,30,193,31,185,31,230,31,129,31,194,31,250,31,12,31,47,31,47,30,225,31,18,31,18,30,125,31,138,31,203,31,203,30,203,29,121,31,121,30,140,31,140,30,182,31,60,31,37,31,228,31,82,31,218,31,69,31,17,31,247,31,67,31,118,31,118,30,110,31,123,31,123,30,228,31,228,30,99,31,99,30,99,29,33,31,215,31,101,31,88,31,134,31,192,31,99,31,99,30,2,31,2,30,109,31,22,31,221,31,138,31,138,30,79,31,34,31,158,31,128,31,212,31,104,31,123,31,228,31,65,31,45,31,69,31,192,31,192,30,192,29,223,31,223,30,72,31,45,31,127,31,235,31,151,31,64,31,91,31,134,31,225,31,19,31,48,31,199,31,160,31,17,31,7,31,7,30,7,29,184,31,133,31,133,30,154,31,118,31,182,31,174,31,174,30,212,31,142,31,6,31,6,30,57,31,130,31,212,31,157,31,69,31,7,31,10,31,10,30,221,31,32,31,221,31,255,31,248,31,25,31,84,31,63,31,244,31,170,31,30,31,30,30,30,29,100,31,136,31,199,31,69,31,17,31,45,31,205,31,199,31,117,31,117,30,65,31,65,30,238,31,8,31,8,30,8,29,8,28,232,31,46,31,46,30,128,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
