-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_264 is
end project_tb_264;

architecture project_tb_arch_264 of project_tb_264 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 916;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (217,0,24,0,170,0,0,0,89,0,0,0,134,0,173,0,83,0,145,0,0,0,89,0,163,0,231,0,149,0,130,0,57,0,31,0,151,0,4,0,0,0,144,0,119,0,0,0,60,0,157,0,108,0,52,0,181,0,0,0,0,0,177,0,138,0,21,0,120,0,0,0,151,0,247,0,198,0,122,0,189,0,17,0,0,0,238,0,119,0,88,0,102,0,0,0,115,0,81,0,84,0,45,0,64,0,20,0,79,0,120,0,44,0,76,0,219,0,103,0,102,0,101,0,0,0,133,0,0,0,80,0,193,0,95,0,11,0,103,0,62,0,235,0,194,0,66,0,23,0,244,0,1,0,244,0,210,0,4,0,210,0,212,0,242,0,0,0,112,0,99,0,0,0,26,0,104,0,39,0,0,0,191,0,184,0,128,0,220,0,227,0,0,0,123,0,163,0,178,0,209,0,190,0,0,0,0,0,247,0,173,0,156,0,24,0,246,0,7,0,0,0,0,0,237,0,104,0,201,0,229,0,0,0,127,0,183,0,6,0,212,0,255,0,172,0,245,0,19,0,43,0,0,0,0,0,17,0,244,0,3,0,131,0,59,0,75,0,136,0,162,0,202,0,128,0,133,0,9,0,164,0,253,0,191,0,15,0,0,0,77,0,103,0,167,0,66,0,0,0,128,0,116,0,222,0,68,0,155,0,109,0,0,0,8,0,10,0,25,0,41,0,37,0,145,0,0,0,164,0,217,0,16,0,26,0,0,0,218,0,42,0,0,0,0,0,0,0,213,0,0,0,43,0,144,0,49,0,72,0,68,0,197,0,172,0,29,0,233,0,201,0,227,0,202,0,21,0,101,0,133,0,133,0,188,0,73,0,0,0,135,0,164,0,0,0,38,0,0,0,240,0,0,0,184,0,82,0,221,0,107,0,74,0,180,0,0,0,0,0,179,0,0,0,78,0,215,0,110,0,135,0,228,0,15,0,225,0,140,0,202,0,251,0,222,0,0,0,0,0,25,0,5,0,241,0,0,0,97,0,4,0,54,0,118,0,134,0,217,0,190,0,245,0,121,0,215,0,147,0,122,0,156,0,80,0,99,0,0,0,35,0,170,0,175,0,5,0,0,0,199,0,162,0,139,0,0,0,163,0,147,0,101,0,90,0,94,0,0,0,253,0,189,0,0,0,77,0,243,0,156,0,0,0,0,0,64,0,0,0,34,0,0,0,155,0,236,0,0,0,52,0,0,0,92,0,0,0,0,0,0,0,44,0,70,0,49,0,162,0,232,0,232,0,160,0,12,0,0,0,217,0,145,0,103,0,215,0,248,0,52,0,0,0,74,0,0,0,0,0,253,0,255,0,0,0,92,0,168,0,0,0,21,0,33,0,131,0,0,0,249,0,186,0,229,0,0,0,221,0,0,0,181,0,250,0,0,0,0,0,84,0,184,0,156,0,32,0,115,0,41,0,235,0,99,0,96,0,0,0,54,0,104,0,0,0,142,0,249,0,240,0,191,0,183,0,48,0,177,0,186,0,11,0,166,0,124,0,229,0,5,0,136,0,224,0,110,0,0,0,68,0,98,0,0,0,250,0,206,0,0,0,125,0,0,0,91,0,133,0,40,0,78,0,0,0,138,0,200,0,9,0,71,0,13,0,120,0,232,0,96,0,214,0,73,0,87,0,60,0,129,0,42,0,0,0,0,0,188,0,31,0,131,0,94,0,67,0,45,0,96,0,76,0,191,0,84,0,0,0,0,0,12,0,25,0,42,0,246,0,58,0,68,0,242,0,194,0,89,0,64,0,190,0,0,0,48,0,77,0,100,0,88,0,94,0,121,0,23,0,181,0,137,0,3,0,29,0,0,0,187,0,91,0,99,0,28,0,0,0,0,0,184,0,112,0,119,0,172,0,199,0,140,0,0,0,0,0,33,0,235,0,61,0,96,0,223,0,66,0,178,0,254,0,144,0,135,0,164,0,141,0,152,0,223,0,216,0,76,0,167,0,207,0,220,0,71,0,151,0,0,0,37,0,194,0,0,0,152,0,0,0,208,0,165,0,27,0,102,0,74,0,48,0,231,0,0,0,250,0,82,0,134,0,0,0,0,0,0,0,0,0,152,0,205,0,0,0,0,0,0,0,207,0,144,0,236,0,28,0,168,0,0,0,43,0,184,0,70,0,85,0,0,0,0,0,1,0,244,0,51,0,0,0,136,0,255,0,156,0,162,0,23,0,232,0,0,0,121,0,25,0,22,0,199,0,0,0,88,0,215,0,198,0,0,0,0,0,152,0,159,0,0,0,0,0,56,0,0,0,90,0,0,0,204,0,0,0,85,0,13,0,212,0,91,0,225,0,0,0,0,0,186,0,128,0,186,0,97,0,200,0,0,0,205,0,0,0,147,0,70,0,106,0,0,0,134,0,234,0,0,0,87,0,103,0,200,0,0,0,54,0,93,0,182,0,158,0,219,0,89,0,9,0,0,0,51,0,53,0,21,0,0,0,151,0,49,0,0,0,0,0,59,0,194,0,166,0,212,0,32,0,18,0,58,0,205,0,0,0,0,0,87,0,0,0,175,0,52,0,0,0,111,0,0,0,126,0,229,0,236,0,175,0,115,0,162,0,198,0,158,0,243,0,0,0,188,0,117,0,25,0,85,0,160,0,29,0,69,0,0,0,15,0,131,0,239,0,193,0,49,0,0,0,73,0,69,0,212,0,199,0,43,0,135,0,0,0,0,0,0,0,0,0,0,0,83,0,255,0,0,0,1,0,135,0,223,0,85,0,107,0,0,0,58,0,237,0,3,0,189,0,153,0,181,0,203,0,126,0,52,0,138,0,3,0,0,0,95,0,211,0,39,0,154,0,26,0,165,0,60,0,177,0,250,0,0,0,0,0,1,0,103,0,0,0,0,0,19,0,207,0,194,0,0,0,0,0,162,0,130,0,146,0,159,0,0,0,33,0,242,0,72,0,228,0,148,0,34,0,68,0,169,0,77,0,0,0,11,0,0,0,38,0,193,0,196,0,55,0,241,0,254,0,218,0,0,0,0,0,22,0,35,0,112,0,51,0,0,0,152,0,21,0,244,0,58,0,76,0,0,0,0,0,59,0,180,0,139,0,221,0,149,0,74,0,90,0,73,0,130,0,200,0,0,0,0,0,249,0,161,0,0,0,78,0,27,0,252,0,251,0,103,0,24,0,140,0,0,0,46,0,134,0,29,0,154,0,48,0,155,0,16,0,1,0,39,0,0,0,248,0,177,0,196,0,22,0,0,0,158,0,38,0,98,0,27,0,201,0,253,0,35,0,246,0,163,0,253,0,40,0,177,0,56,0,234,0,0,0,161,0,147,0,62,0,23,0,132,0,98,0,90,0,71,0,114,0,100,0,26,0,113,0,19,0,199,0,0,0,136,0,81,0,235,0,0,0,0,0,166,0,135,0,23,0,188,0,168,0,65,0,246,0,0,0,106,0,222,0,0,0,87,0,248,0,113,0,224,0,190,0,100,0,141,0,0,0,188,0,49,0,81,0,146,0,177,0,33,0,139,0,110,0,182,0,0,0,18,0,74,0,187,0,0,0,15,0,98,0,54,0,186,0,0,0,213,0,73,0,0,0,19,0,207,0,79,0,71,0,189,0,82,0,65,0,17,0,0,0,55,0,28,0,123,0,225,0,165,0,62,0,219,0,82,0,13,0,0,0,163,0,0,0,0,0,139,0,231,0,0,0,0,0,222,0,225,0,50,0,253,0,0,0,0,0,112,0,12,0,104,0,127,0,40,0,78,0,7,0,0,0,112,0,240,0,0,0,146,0,0,0,173,0,84,0,112,0,122,0,5,0,167,0,79,0,58,0,116,0,3,0,128,0,53,0,0,0,119,0,0,0,124,0,154,0,103,0,109,0,211,0,100,0,148,0,157,0,236,0,0,0,104,0,34,0,226,0,140,0,0,0,16,0,232,0,209,0,150,0,95,0,161,0,0,0,0,0,0,0,75,0,117,0,150,0,164,0,106,0,191,0,0,0,0,0,157,0,22,0,102,0,0,0,116,0,157,0,199,0,251,0,0,0,94,0,216,0,210,0,204,0,0,0,0,0,235,0,139,0,27,0);
signal scenario_full  : scenario_type := (217,31,24,31,170,31,170,30,89,31,89,30,134,31,173,31,83,31,145,31,145,30,89,31,163,31,231,31,149,31,130,31,57,31,31,31,151,31,4,31,4,30,144,31,119,31,119,30,60,31,157,31,108,31,52,31,181,31,181,30,181,29,177,31,138,31,21,31,120,31,120,30,151,31,247,31,198,31,122,31,189,31,17,31,17,30,238,31,119,31,88,31,102,31,102,30,115,31,81,31,84,31,45,31,64,31,20,31,79,31,120,31,44,31,76,31,219,31,103,31,102,31,101,31,101,30,133,31,133,30,80,31,193,31,95,31,11,31,103,31,62,31,235,31,194,31,66,31,23,31,244,31,1,31,244,31,210,31,4,31,210,31,212,31,242,31,242,30,112,31,99,31,99,30,26,31,104,31,39,31,39,30,191,31,184,31,128,31,220,31,227,31,227,30,123,31,163,31,178,31,209,31,190,31,190,30,190,29,247,31,173,31,156,31,24,31,246,31,7,31,7,30,7,29,237,31,104,31,201,31,229,31,229,30,127,31,183,31,6,31,212,31,255,31,172,31,245,31,19,31,43,31,43,30,43,29,17,31,244,31,3,31,131,31,59,31,75,31,136,31,162,31,202,31,128,31,133,31,9,31,164,31,253,31,191,31,15,31,15,30,77,31,103,31,167,31,66,31,66,30,128,31,116,31,222,31,68,31,155,31,109,31,109,30,8,31,10,31,25,31,41,31,37,31,145,31,145,30,164,31,217,31,16,31,26,31,26,30,218,31,42,31,42,30,42,29,42,28,213,31,213,30,43,31,144,31,49,31,72,31,68,31,197,31,172,31,29,31,233,31,201,31,227,31,202,31,21,31,101,31,133,31,133,31,188,31,73,31,73,30,135,31,164,31,164,30,38,31,38,30,240,31,240,30,184,31,82,31,221,31,107,31,74,31,180,31,180,30,180,29,179,31,179,30,78,31,215,31,110,31,135,31,228,31,15,31,225,31,140,31,202,31,251,31,222,31,222,30,222,29,25,31,5,31,241,31,241,30,97,31,4,31,54,31,118,31,134,31,217,31,190,31,245,31,121,31,215,31,147,31,122,31,156,31,80,31,99,31,99,30,35,31,170,31,175,31,5,31,5,30,199,31,162,31,139,31,139,30,163,31,147,31,101,31,90,31,94,31,94,30,253,31,189,31,189,30,77,31,243,31,156,31,156,30,156,29,64,31,64,30,34,31,34,30,155,31,236,31,236,30,52,31,52,30,92,31,92,30,92,29,92,28,44,31,70,31,49,31,162,31,232,31,232,31,160,31,12,31,12,30,217,31,145,31,103,31,215,31,248,31,52,31,52,30,74,31,74,30,74,29,253,31,255,31,255,30,92,31,168,31,168,30,21,31,33,31,131,31,131,30,249,31,186,31,229,31,229,30,221,31,221,30,181,31,250,31,250,30,250,29,84,31,184,31,156,31,32,31,115,31,41,31,235,31,99,31,96,31,96,30,54,31,104,31,104,30,142,31,249,31,240,31,191,31,183,31,48,31,177,31,186,31,11,31,166,31,124,31,229,31,5,31,136,31,224,31,110,31,110,30,68,31,98,31,98,30,250,31,206,31,206,30,125,31,125,30,91,31,133,31,40,31,78,31,78,30,138,31,200,31,9,31,71,31,13,31,120,31,232,31,96,31,214,31,73,31,87,31,60,31,129,31,42,31,42,30,42,29,188,31,31,31,131,31,94,31,67,31,45,31,96,31,76,31,191,31,84,31,84,30,84,29,12,31,25,31,42,31,246,31,58,31,68,31,242,31,194,31,89,31,64,31,190,31,190,30,48,31,77,31,100,31,88,31,94,31,121,31,23,31,181,31,137,31,3,31,29,31,29,30,187,31,91,31,99,31,28,31,28,30,28,29,184,31,112,31,119,31,172,31,199,31,140,31,140,30,140,29,33,31,235,31,61,31,96,31,223,31,66,31,178,31,254,31,144,31,135,31,164,31,141,31,152,31,223,31,216,31,76,31,167,31,207,31,220,31,71,31,151,31,151,30,37,31,194,31,194,30,152,31,152,30,208,31,165,31,27,31,102,31,74,31,48,31,231,31,231,30,250,31,82,31,134,31,134,30,134,29,134,28,134,27,152,31,205,31,205,30,205,29,205,28,207,31,144,31,236,31,28,31,168,31,168,30,43,31,184,31,70,31,85,31,85,30,85,29,1,31,244,31,51,31,51,30,136,31,255,31,156,31,162,31,23,31,232,31,232,30,121,31,25,31,22,31,199,31,199,30,88,31,215,31,198,31,198,30,198,29,152,31,159,31,159,30,159,29,56,31,56,30,90,31,90,30,204,31,204,30,85,31,13,31,212,31,91,31,225,31,225,30,225,29,186,31,128,31,186,31,97,31,200,31,200,30,205,31,205,30,147,31,70,31,106,31,106,30,134,31,234,31,234,30,87,31,103,31,200,31,200,30,54,31,93,31,182,31,158,31,219,31,89,31,9,31,9,30,51,31,53,31,21,31,21,30,151,31,49,31,49,30,49,29,59,31,194,31,166,31,212,31,32,31,18,31,58,31,205,31,205,30,205,29,87,31,87,30,175,31,52,31,52,30,111,31,111,30,126,31,229,31,236,31,175,31,115,31,162,31,198,31,158,31,243,31,243,30,188,31,117,31,25,31,85,31,160,31,29,31,69,31,69,30,15,31,131,31,239,31,193,31,49,31,49,30,73,31,69,31,212,31,199,31,43,31,135,31,135,30,135,29,135,28,135,27,135,26,83,31,255,31,255,30,1,31,135,31,223,31,85,31,107,31,107,30,58,31,237,31,3,31,189,31,153,31,181,31,203,31,126,31,52,31,138,31,3,31,3,30,95,31,211,31,39,31,154,31,26,31,165,31,60,31,177,31,250,31,250,30,250,29,1,31,103,31,103,30,103,29,19,31,207,31,194,31,194,30,194,29,162,31,130,31,146,31,159,31,159,30,33,31,242,31,72,31,228,31,148,31,34,31,68,31,169,31,77,31,77,30,11,31,11,30,38,31,193,31,196,31,55,31,241,31,254,31,218,31,218,30,218,29,22,31,35,31,112,31,51,31,51,30,152,31,21,31,244,31,58,31,76,31,76,30,76,29,59,31,180,31,139,31,221,31,149,31,74,31,90,31,73,31,130,31,200,31,200,30,200,29,249,31,161,31,161,30,78,31,27,31,252,31,251,31,103,31,24,31,140,31,140,30,46,31,134,31,29,31,154,31,48,31,155,31,16,31,1,31,39,31,39,30,248,31,177,31,196,31,22,31,22,30,158,31,38,31,98,31,27,31,201,31,253,31,35,31,246,31,163,31,253,31,40,31,177,31,56,31,234,31,234,30,161,31,147,31,62,31,23,31,132,31,98,31,90,31,71,31,114,31,100,31,26,31,113,31,19,31,199,31,199,30,136,31,81,31,235,31,235,30,235,29,166,31,135,31,23,31,188,31,168,31,65,31,246,31,246,30,106,31,222,31,222,30,87,31,248,31,113,31,224,31,190,31,100,31,141,31,141,30,188,31,49,31,81,31,146,31,177,31,33,31,139,31,110,31,182,31,182,30,18,31,74,31,187,31,187,30,15,31,98,31,54,31,186,31,186,30,213,31,73,31,73,30,19,31,207,31,79,31,71,31,189,31,82,31,65,31,17,31,17,30,55,31,28,31,123,31,225,31,165,31,62,31,219,31,82,31,13,31,13,30,163,31,163,30,163,29,139,31,231,31,231,30,231,29,222,31,225,31,50,31,253,31,253,30,253,29,112,31,12,31,104,31,127,31,40,31,78,31,7,31,7,30,112,31,240,31,240,30,146,31,146,30,173,31,84,31,112,31,122,31,5,31,167,31,79,31,58,31,116,31,3,31,128,31,53,31,53,30,119,31,119,30,124,31,154,31,103,31,109,31,211,31,100,31,148,31,157,31,236,31,236,30,104,31,34,31,226,31,140,31,140,30,16,31,232,31,209,31,150,31,95,31,161,31,161,30,161,29,161,28,75,31,117,31,150,31,164,31,106,31,191,31,191,30,191,29,157,31,22,31,102,31,102,30,116,31,157,31,199,31,251,31,251,30,94,31,216,31,210,31,204,31,204,30,204,29,235,31,139,31,27,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
