-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 758;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (244,0,128,0,107,0,161,0,67,0,0,0,253,0,75,0,198,0,168,0,209,0,111,0,155,0,223,0,0,0,27,0,0,0,2,0,36,0,200,0,115,0,140,0,62,0,143,0,96,0,0,0,226,0,74,0,4,0,57,0,54,0,19,0,161,0,178,0,0,0,160,0,122,0,0,0,228,0,0,0,167,0,175,0,94,0,0,0,12,0,65,0,78,0,46,0,179,0,0,0,0,0,0,0,144,0,183,0,115,0,194,0,95,0,20,0,163,0,85,0,95,0,141,0,181,0,11,0,198,0,41,0,189,0,158,0,82,0,190,0,203,0,0,0,162,0,246,0,0,0,100,0,2,0,87,0,144,0,96,0,199,0,247,0,250,0,198,0,156,0,107,0,131,0,0,0,213,0,89,0,5,0,165,0,99,0,14,0,196,0,197,0,136,0,0,0,0,0,97,0,95,0,180,0,150,0,18,0,226,0,167,0,0,0,168,0,206,0,186,0,166,0,192,0,168,0,180,0,153,0,55,0,0,0,4,0,37,0,211,0,0,0,3,0,95,0,0,0,0,0,94,0,200,0,211,0,28,0,160,0,56,0,50,0,122,0,232,0,45,0,40,0,188,0,0,0,41,0,0,0,114,0,137,0,245,0,55,0,182,0,0,0,28,0,138,0,58,0,244,0,247,0,137,0,146,0,253,0,76,0,141,0,0,0,16,0,0,0,36,0,245,0,180,0,57,0,0,0,0,0,102,0,0,0,148,0,110,0,190,0,213,0,48,0,108,0,56,0,225,0,0,0,15,0,0,0,0,0,0,0,0,0,56,0,141,0,222,0,218,0,0,0,63,0,86,0,158,0,226,0,0,0,54,0,0,0,125,0,94,0,116,0,132,0,87,0,0,0,208,0,0,0,125,0,41,0,0,0,194,0,230,0,0,0,160,0,200,0,0,0,26,0,116,0,151,0,0,0,148,0,149,0,0,0,219,0,114,0,23,0,202,0,54,0,45,0,45,0,221,0,6,0,76,0,245,0,24,0,57,0,230,0,100,0,253,0,13,0,97,0,247,0,0,0,228,0,0,0,141,0,0,0,192,0,30,0,209,0,31,0,61,0,0,0,215,0,0,0,0,0,24,0,23,0,208,0,126,0,159,0,0,0,10,0,32,0,219,0,0,0,0,0,222,0,7,0,210,0,175,0,254,0,199,0,191,0,225,0,10,0,111,0,244,0,224,0,0,0,56,0,60,0,255,0,107,0,0,0,154,0,206,0,50,0,66,0,120,0,229,0,0,0,34,0,254,0,133,0,199,0,172,0,0,0,39,0,0,0,0,0,0,0,146,0,117,0,0,0,26,0,62,0,37,0,254,0,0,0,22,0,36,0,103,0,130,0,147,0,68,0,179,0,0,0,0,0,175,0,12,0,131,0,153,0,214,0,0,0,4,0,166,0,51,0,51,0,71,0,0,0,49,0,194,0,0,0,247,0,193,0,0,0,0,0,135,0,232,0,176,0,195,0,215,0,164,0,19,0,16,0,26,0,0,0,203,0,53,0,35,0,226,0,0,0,0,0,76,0,199,0,226,0,147,0,0,0,200,0,216,0,0,0,43,0,187,0,141,0,186,0,0,0,0,0,0,0,101,0,38,0,0,0,215,0,0,0,0,0,0,0,165,0,105,0,39,0,53,0,0,0,0,0,139,0,68,0,0,0,168,0,0,0,162,0,192,0,218,0,79,0,238,0,212,0,22,0,88,0,87,0,0,0,54,0,42,0,122,0,0,0,7,0,42,0,178,0,234,0,65,0,228,0,247,0,158,0,254,0,15,0,43,0,83,0,105,0,225,0,0,0,189,0,34,0,59,0,31,0,83,0,134,0,95,0,4,0,143,0,129,0,53,0,242,0,23,0,124,0,224,0,0,0,218,0,0,0,88,0,39,0,82,0,130,0,0,0,0,0,68,0,204,0,86,0,3,0,181,0,120,0,0,0,254,0,212,0,134,0,182,0,81,0,44,0,53,0,109,0,169,0,146,0,38,0,20,0,0,0,115,0,0,0,70,0,0,0,248,0,149,0,66,0,218,0,235,0,241,0,171,0,139,0,0,0,66,0,54,0,28,0,240,0,36,0,118,0,36,0,58,0,101,0,45,0,0,0,227,0,0,0,247,0,0,0,106,0,232,0,172,0,75,0,0,0,223,0,33,0,122,0,115,0,23,0,22,0,232,0,71,0,0,0,82,0,169,0,250,0,55,0,214,0,0,0,0,0,43,0,236,0,133,0,58,0,0,0,177,0,129,0,88,0,246,0,160,0,0,0,195,0,112,0,0,0,0,0,51,0,54,0,63,0,143,0,249,0,121,0,48,0,201,0,0,0,0,0,247,0,0,0,20,0,20,0,185,0,45,0,185,0,143,0,0,0,165,0,74,0,0,0,0,0,150,0,36,0,34,0,18,0,0,0,78,0,56,0,166,0,162,0,130,0,251,0,127,0,0,0,131,0,0,0,73,0,231,0,194,0,14,0,194,0,225,0,13,0,191,0,190,0,138,0,71,0,0,0,36,0,211,0,196,0,0,0,238,0,126,0,0,0,225,0,0,0,0,0,0,0,33,0,241,0,8,0,200,0,0,0,58,0,0,0,66,0,82,0,71,0,27,0,93,0,181,0,0,0,0,0,187,0,143,0,0,0,171,0,78,0,13,0,67,0,44,0,204,0,42,0,0,0,228,0,5,0,32,0,226,0,40,0,152,0,205,0,82,0,242,0,208,0,255,0,127,0,249,0,57,0,189,0,16,0,83,0,144,0,165,0,0,0,0,0,84,0,42,0,102,0,0,0,0,0,45,0,37,0,67,0,239,0,89,0,0,0,114,0,89,0,10,0,0,0,0,0,117,0,0,0,0,0,244,0,0,0,0,0,1,0,46,0,0,0,0,0,72,0,16,0,147,0,128,0,13,0,172,0,0,0,62,0,7,0,0,0,0,0,28,0,99,0,66,0,5,0,116,0,115,0,0,0,0,0,0,0,187,0,70,0,86,0,210,0,153,0,250,0,0,0,2,0,143,0,0,0,20,0,0,0,235,0,129,0,223,0,96,0,0,0,0,0,42,0,87,0,88,0,233,0,0,0,0,0,147,0,131,0,204,0,70,0,0,0,91,0,179,0,230,0,138,0,143,0,204,0,9,0,108,0,181,0,4,0,119,0,228,0,104,0,38,0,140,0,137,0,0,0,36,0,120,0,47,0,99,0,33,0,163,0,54,0,36,0,19,0,18,0,0,0,181,0,84,0,68,0,56,0,23,0,79,0,0,0,181,0,30,0,178,0,162,0,152,0,225,0,34,0,0,0,161,0,0,0,219,0,76,0,215,0,129,0,0,0,133,0,0,0,41,0,1,0,96,0,0,0,176,0);
signal scenario_full  : scenario_type := (244,31,128,31,107,31,161,31,67,31,67,30,253,31,75,31,198,31,168,31,209,31,111,31,155,31,223,31,223,30,27,31,27,30,2,31,36,31,200,31,115,31,140,31,62,31,143,31,96,31,96,30,226,31,74,31,4,31,57,31,54,31,19,31,161,31,178,31,178,30,160,31,122,31,122,30,228,31,228,30,167,31,175,31,94,31,94,30,12,31,65,31,78,31,46,31,179,31,179,30,179,29,179,28,144,31,183,31,115,31,194,31,95,31,20,31,163,31,85,31,95,31,141,31,181,31,11,31,198,31,41,31,189,31,158,31,82,31,190,31,203,31,203,30,162,31,246,31,246,30,100,31,2,31,87,31,144,31,96,31,199,31,247,31,250,31,198,31,156,31,107,31,131,31,131,30,213,31,89,31,5,31,165,31,99,31,14,31,196,31,197,31,136,31,136,30,136,29,97,31,95,31,180,31,150,31,18,31,226,31,167,31,167,30,168,31,206,31,186,31,166,31,192,31,168,31,180,31,153,31,55,31,55,30,4,31,37,31,211,31,211,30,3,31,95,31,95,30,95,29,94,31,200,31,211,31,28,31,160,31,56,31,50,31,122,31,232,31,45,31,40,31,188,31,188,30,41,31,41,30,114,31,137,31,245,31,55,31,182,31,182,30,28,31,138,31,58,31,244,31,247,31,137,31,146,31,253,31,76,31,141,31,141,30,16,31,16,30,36,31,245,31,180,31,57,31,57,30,57,29,102,31,102,30,148,31,110,31,190,31,213,31,48,31,108,31,56,31,225,31,225,30,15,31,15,30,15,29,15,28,15,27,56,31,141,31,222,31,218,31,218,30,63,31,86,31,158,31,226,31,226,30,54,31,54,30,125,31,94,31,116,31,132,31,87,31,87,30,208,31,208,30,125,31,41,31,41,30,194,31,230,31,230,30,160,31,200,31,200,30,26,31,116,31,151,31,151,30,148,31,149,31,149,30,219,31,114,31,23,31,202,31,54,31,45,31,45,31,221,31,6,31,76,31,245,31,24,31,57,31,230,31,100,31,253,31,13,31,97,31,247,31,247,30,228,31,228,30,141,31,141,30,192,31,30,31,209,31,31,31,61,31,61,30,215,31,215,30,215,29,24,31,23,31,208,31,126,31,159,31,159,30,10,31,32,31,219,31,219,30,219,29,222,31,7,31,210,31,175,31,254,31,199,31,191,31,225,31,10,31,111,31,244,31,224,31,224,30,56,31,60,31,255,31,107,31,107,30,154,31,206,31,50,31,66,31,120,31,229,31,229,30,34,31,254,31,133,31,199,31,172,31,172,30,39,31,39,30,39,29,39,28,146,31,117,31,117,30,26,31,62,31,37,31,254,31,254,30,22,31,36,31,103,31,130,31,147,31,68,31,179,31,179,30,179,29,175,31,12,31,131,31,153,31,214,31,214,30,4,31,166,31,51,31,51,31,71,31,71,30,49,31,194,31,194,30,247,31,193,31,193,30,193,29,135,31,232,31,176,31,195,31,215,31,164,31,19,31,16,31,26,31,26,30,203,31,53,31,35,31,226,31,226,30,226,29,76,31,199,31,226,31,147,31,147,30,200,31,216,31,216,30,43,31,187,31,141,31,186,31,186,30,186,29,186,28,101,31,38,31,38,30,215,31,215,30,215,29,215,28,165,31,105,31,39,31,53,31,53,30,53,29,139,31,68,31,68,30,168,31,168,30,162,31,192,31,218,31,79,31,238,31,212,31,22,31,88,31,87,31,87,30,54,31,42,31,122,31,122,30,7,31,42,31,178,31,234,31,65,31,228,31,247,31,158,31,254,31,15,31,43,31,83,31,105,31,225,31,225,30,189,31,34,31,59,31,31,31,83,31,134,31,95,31,4,31,143,31,129,31,53,31,242,31,23,31,124,31,224,31,224,30,218,31,218,30,88,31,39,31,82,31,130,31,130,30,130,29,68,31,204,31,86,31,3,31,181,31,120,31,120,30,254,31,212,31,134,31,182,31,81,31,44,31,53,31,109,31,169,31,146,31,38,31,20,31,20,30,115,31,115,30,70,31,70,30,248,31,149,31,66,31,218,31,235,31,241,31,171,31,139,31,139,30,66,31,54,31,28,31,240,31,36,31,118,31,36,31,58,31,101,31,45,31,45,30,227,31,227,30,247,31,247,30,106,31,232,31,172,31,75,31,75,30,223,31,33,31,122,31,115,31,23,31,22,31,232,31,71,31,71,30,82,31,169,31,250,31,55,31,214,31,214,30,214,29,43,31,236,31,133,31,58,31,58,30,177,31,129,31,88,31,246,31,160,31,160,30,195,31,112,31,112,30,112,29,51,31,54,31,63,31,143,31,249,31,121,31,48,31,201,31,201,30,201,29,247,31,247,30,20,31,20,31,185,31,45,31,185,31,143,31,143,30,165,31,74,31,74,30,74,29,150,31,36,31,34,31,18,31,18,30,78,31,56,31,166,31,162,31,130,31,251,31,127,31,127,30,131,31,131,30,73,31,231,31,194,31,14,31,194,31,225,31,13,31,191,31,190,31,138,31,71,31,71,30,36,31,211,31,196,31,196,30,238,31,126,31,126,30,225,31,225,30,225,29,225,28,33,31,241,31,8,31,200,31,200,30,58,31,58,30,66,31,82,31,71,31,27,31,93,31,181,31,181,30,181,29,187,31,143,31,143,30,171,31,78,31,13,31,67,31,44,31,204,31,42,31,42,30,228,31,5,31,32,31,226,31,40,31,152,31,205,31,82,31,242,31,208,31,255,31,127,31,249,31,57,31,189,31,16,31,83,31,144,31,165,31,165,30,165,29,84,31,42,31,102,31,102,30,102,29,45,31,37,31,67,31,239,31,89,31,89,30,114,31,89,31,10,31,10,30,10,29,117,31,117,30,117,29,244,31,244,30,244,29,1,31,46,31,46,30,46,29,72,31,16,31,147,31,128,31,13,31,172,31,172,30,62,31,7,31,7,30,7,29,28,31,99,31,66,31,5,31,116,31,115,31,115,30,115,29,115,28,187,31,70,31,86,31,210,31,153,31,250,31,250,30,2,31,143,31,143,30,20,31,20,30,235,31,129,31,223,31,96,31,96,30,96,29,42,31,87,31,88,31,233,31,233,30,233,29,147,31,131,31,204,31,70,31,70,30,91,31,179,31,230,31,138,31,143,31,204,31,9,31,108,31,181,31,4,31,119,31,228,31,104,31,38,31,140,31,137,31,137,30,36,31,120,31,47,31,99,31,33,31,163,31,54,31,36,31,19,31,18,31,18,30,181,31,84,31,68,31,56,31,23,31,79,31,79,30,181,31,30,31,178,31,162,31,152,31,225,31,34,31,34,30,161,31,161,30,219,31,76,31,215,31,129,31,129,30,133,31,133,30,41,31,1,31,96,31,96,30,176,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
