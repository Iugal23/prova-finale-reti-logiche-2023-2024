-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_15 is
end project_tb_15;

architecture project_tb_arch_15 of project_tb_15 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 281;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (39,0,160,0,50,0,169,0,70,0,0,0,12,0,155,0,194,0,178,0,0,0,216,0,171,0,89,0,30,0,247,0,67,0,57,0,73,0,27,0,190,0,36,0,234,0,82,0,227,0,0,0,175,0,28,0,28,0,59,0,180,0,213,0,124,0,0,0,138,0,232,0,234,0,217,0,130,0,49,0,233,0,53,0,138,0,199,0,36,0,0,0,157,0,35,0,0,0,194,0,97,0,66,0,0,0,28,0,178,0,148,0,246,0,0,0,79,0,0,0,115,0,190,0,120,0,0,0,171,0,181,0,0,0,67,0,154,0,147,0,59,0,0,0,181,0,134,0,0,0,0,0,0,0,90,0,14,0,15,0,237,0,82,0,11,0,209,0,0,0,0,0,33,0,0,0,0,0,163,0,65,0,88,0,207,0,155,0,203,0,131,0,169,0,0,0,60,0,117,0,71,0,146,0,109,0,213,0,0,0,0,0,146,0,1,0,197,0,148,0,231,0,72,0,86,0,42,0,160,0,241,0,14,0,0,0,116,0,207,0,0,0,111,0,58,0,164,0,46,0,3,0,157,0,114,0,88,0,121,0,252,0,116,0,95,0,9,0,253,0,193,0,111,0,191,0,13,0,68,0,28,0,26,0,0,0,223,0,172,0,226,0,250,0,82,0,105,0,186,0,185,0,140,0,0,0,242,0,5,0,172,0,0,0,2,0,117,0,11,0,73,0,6,0,114,0,118,0,175,0,0,0,224,0,110,0,0,0,207,0,12,0,0,0,24,0,57,0,96,0,0,0,0,0,169,0,176,0,59,0,245,0,102,0,105,0,128,0,0,0,231,0,66,0,0,0,60,0,42,0,0,0,239,0,179,0,202,0,108,0,214,0,229,0,105,0,182,0,0,0,0,0,177,0,45,0,249,0,108,0,159,0,164,0,0,0,130,0,56,0,163,0,189,0,196,0,124,0,27,0,0,0,93,0,69,0,170,0,122,0,110,0,0,0,48,0,118,0,108,0,34,0,74,0,82,0,15,0,78,0,0,0,17,0,0,0,117,0,145,0,0,0,216,0,169,0,179,0,0,0,234,0,176,0,88,0,18,0,246,0,150,0,51,0,177,0,0,0,145,0,145,0,13,0,234,0,50,0,6,0,64,0,38,0,65,0,50,0,36,0,16,0,0,0,0,0,252,0,228,0,115,0,108,0,219,0,142,0,65,0,173,0,194,0,9,0,0,0,233,0,209,0,102,0,100,0,0,0,110,0,0,0);
signal scenario_full  : scenario_type := (39,31,160,31,50,31,169,31,70,31,70,30,12,31,155,31,194,31,178,31,178,30,216,31,171,31,89,31,30,31,247,31,67,31,57,31,73,31,27,31,190,31,36,31,234,31,82,31,227,31,227,30,175,31,28,31,28,31,59,31,180,31,213,31,124,31,124,30,138,31,232,31,234,31,217,31,130,31,49,31,233,31,53,31,138,31,199,31,36,31,36,30,157,31,35,31,35,30,194,31,97,31,66,31,66,30,28,31,178,31,148,31,246,31,246,30,79,31,79,30,115,31,190,31,120,31,120,30,171,31,181,31,181,30,67,31,154,31,147,31,59,31,59,30,181,31,134,31,134,30,134,29,134,28,90,31,14,31,15,31,237,31,82,31,11,31,209,31,209,30,209,29,33,31,33,30,33,29,163,31,65,31,88,31,207,31,155,31,203,31,131,31,169,31,169,30,60,31,117,31,71,31,146,31,109,31,213,31,213,30,213,29,146,31,1,31,197,31,148,31,231,31,72,31,86,31,42,31,160,31,241,31,14,31,14,30,116,31,207,31,207,30,111,31,58,31,164,31,46,31,3,31,157,31,114,31,88,31,121,31,252,31,116,31,95,31,9,31,253,31,193,31,111,31,191,31,13,31,68,31,28,31,26,31,26,30,223,31,172,31,226,31,250,31,82,31,105,31,186,31,185,31,140,31,140,30,242,31,5,31,172,31,172,30,2,31,117,31,11,31,73,31,6,31,114,31,118,31,175,31,175,30,224,31,110,31,110,30,207,31,12,31,12,30,24,31,57,31,96,31,96,30,96,29,169,31,176,31,59,31,245,31,102,31,105,31,128,31,128,30,231,31,66,31,66,30,60,31,42,31,42,30,239,31,179,31,202,31,108,31,214,31,229,31,105,31,182,31,182,30,182,29,177,31,45,31,249,31,108,31,159,31,164,31,164,30,130,31,56,31,163,31,189,31,196,31,124,31,27,31,27,30,93,31,69,31,170,31,122,31,110,31,110,30,48,31,118,31,108,31,34,31,74,31,82,31,15,31,78,31,78,30,17,31,17,30,117,31,145,31,145,30,216,31,169,31,179,31,179,30,234,31,176,31,88,31,18,31,246,31,150,31,51,31,177,31,177,30,145,31,145,31,13,31,234,31,50,31,6,31,64,31,38,31,65,31,50,31,36,31,16,31,16,30,16,29,252,31,228,31,115,31,108,31,219,31,142,31,65,31,173,31,194,31,9,31,9,30,233,31,209,31,102,31,100,31,100,30,110,31,110,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
