-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 759;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,38,0,243,0,128,0,52,0,191,0,0,0,151,0,195,0,53,0,81,0,236,0,227,0,91,0,108,0,72,0,16,0,142,0,184,0,0,0,226,0,0,0,125,0,0,0,43,0,65,0,80,0,74,0,38,0,75,0,0,0,135,0,194,0,204,0,240,0,155,0,243,0,0,0,2,0,0,0,70,0,37,0,91,0,0,0,115,0,0,0,173,0,145,0,172,0,21,0,187,0,174,0,170,0,58,0,18,0,127,0,102,0,97,0,255,0,18,0,136,0,34,0,69,0,213,0,60,0,137,0,22,0,255,0,232,0,75,0,0,0,217,0,0,0,103,0,87,0,193,0,0,0,237,0,74,0,179,0,116,0,112,0,50,0,23,0,74,0,126,0,124,0,0,0,0,0,50,0,0,0,240,0,22,0,36,0,11,0,2,0,0,0,216,0,0,0,67,0,202,0,184,0,120,0,66,0,1,0,39,0,0,0,18,0,196,0,0,0,12,0,0,0,112,0,254,0,148,0,172,0,135,0,89,0,170,0,43,0,0,0,200,0,225,0,188,0,213,0,53,0,50,0,183,0,7,0,181,0,125,0,200,0,0,0,201,0,43,0,144,0,3,0,116,0,199,0,102,0,130,0,22,0,200,0,62,0,174,0,11,0,50,0,0,0,46,0,57,0,0,0,0,0,0,0,198,0,247,0,255,0,80,0,155,0,15,0,214,0,46,0,111,0,172,0,31,0,112,0,0,0,15,0,182,0,166,0,72,0,229,0,48,0,91,0,150,0,47,0,36,0,0,0,120,0,0,0,0,0,70,0,141,0,238,0,44,0,23,0,136,0,169,0,27,0,245,0,0,0,132,0,119,0,0,0,113,0,185,0,0,0,0,0,56,0,0,0,165,0,24,0,0,0,0,0,0,0,110,0,100,0,1,0,76,0,255,0,118,0,248,0,0,0,221,0,0,0,0,0,48,0,228,0,0,0,231,0,140,0,199,0,169,0,0,0,0,0,10,0,147,0,61,0,128,0,133,0,142,0,112,0,65,0,243,0,99,0,0,0,3,0,0,0,0,0,201,0,215,0,154,0,240,0,141,0,174,0,0,0,15,0,11,0,194,0,0,0,0,0,0,0,0,0,221,0,203,0,243,0,0,0,114,0,150,0,11,0,157,0,180,0,74,0,245,0,55,0,0,0,161,0,0,0,158,0,0,0,0,0,186,0,177,0,156,0,0,0,165,0,30,0,104,0,101,0,0,0,99,0,0,0,225,0,63,0,148,0,44,0,249,0,0,0,5,0,172,0,177,0,251,0,98,0,0,0,186,0,199,0,0,0,79,0,220,0,122,0,121,0,76,0,239,0,92,0,172,0,0,0,32,0,0,0,192,0,15,0,0,0,206,0,22,0,86,0,56,0,227,0,231,0,218,0,50,0,174,0,238,0,197,0,238,0,0,0,186,0,60,0,152,0,171,0,13,0,0,0,176,0,251,0,73,0,135,0,0,0,91,0,13,0,45,0,10,0,196,0,191,0,242,0,55,0,160,0,89,0,237,0,0,0,146,0,0,0,153,0,224,0,254,0,175,0,67,0,0,0,102,0,232,0,0,0,18,0,15,0,211,0,109,0,41,0,191,0,0,0,48,0,0,0,0,0,194,0,12,0,0,0,0,0,83,0,96,0,0,0,0,0,236,0,139,0,6,0,0,0,193,0,57,0,0,0,116,0,5,0,25,0,0,0,17,0,196,0,239,0,0,0,84,0,6,0,195,0,13,0,81,0,23,0,94,0,233,0,236,0,60,0,0,0,74,0,165,0,11,0,0,0,135,0,44,0,98,0,0,0,242,0,87,0,22,0,36,0,57,0,151,0,76,0,0,0,0,0,147,0,166,0,248,0,119,0,8,0,2,0,70,0,45,0,182,0,191,0,203,0,55,0,89,0,103,0,117,0,169,0,0,0,0,0,160,0,12,0,147,0,210,0,222,0,182,0,233,0,78,0,0,0,186,0,0,0,0,0,63,0,47,0,106,0,17,0,110,0,0,0,177,0,60,0,0,0,42,0,180,0,218,0,0,0,13,0,40,0,125,0,17,0,149,0,1,0,41,0,32,0,241,0,216,0,134,0,74,0,46,0,234,0,7,0,64,0,28,0,172,0,115,0,0,0,127,0,96,0,34,0,0,0,43,0,134,0,162,0,245,0,64,0,192,0,82,0,247,0,72,0,64,0,77,0,149,0,78,0,0,0,164,0,0,0,0,0,32,0,0,0,138,0,44,0,37,0,3,0,0,0,169,0,0,0,152,0,67,0,143,0,0,0,109,0,92,0,190,0,0,0,0,0,167,0,118,0,188,0,143,0,210,0,194,0,44,0,44,0,48,0,141,0,119,0,59,0,126,0,21,0,45,0,0,0,163,0,125,0,250,0,47,0,0,0,131,0,230,0,0,0,110,0,43,0,0,0,41,0,207,0,240,0,0,0,20,0,137,0,164,0,145,0,248,0,21,0,100,0,172,0,1,0,246,0,116,0,26,0,139,0,120,0,210,0,0,0,130,0,0,0,17,0,234,0,38,0,4,0,69,0,0,0,76,0,0,0,57,0,92,0,233,0,75,0,60,0,73,0,223,0,69,0,152,0,111,0,135,0,143,0,156,0,54,0,15,0,136,0,148,0,204,0,182,0,19,0,0,0,235,0,170,0,168,0,0,0,0,0,154,0,159,0,81,0,52,0,180,0,186,0,84,0,162,0,251,0,54,0,0,0,0,0,202,0,127,0,241,0,207,0,153,0,161,0,0,0,82,0,154,0,157,0,136,0,224,0,46,0,0,0,0,0,0,0,112,0,0,0,76,0,170,0,236,0,112,0,205,0,92,0,0,0,211,0,95,0,27,0,150,0,63,0,34,0,197,0,81,0,138,0,119,0,75,0,245,0,43,0,45,0,206,0,148,0,66,0,0,0,124,0,170,0,191,0,205,0,46,0,192,0,165,0,0,0,39,0,139,0,66,0,242,0,233,0,169,0,154,0,212,0,0,0,51,0,0,0,3,0,0,0,165,0,0,0,64,0,28,0,165,0,0,0,0,0,0,0,176,0,22,0,15,0,0,0,70,0,0,0,240,0,52,0,0,0,106,0,135,0,0,0,11,0,89,0,0,0,157,0,176,0,221,0,95,0,49,0,76,0,151,0,194,0,128,0,220,0,89,0,99,0,160,0,0,0,0,0,143,0,178,0,99,0,0,0,98,0,108,0,63,0,242,0,125,0,0,0,45,0,146,0,242,0,206,0,245,0,0,0,220,0,68,0,0,0,67,0,210,0,26,0,118,0,0,0,194,0,0,0,111,0,177,0,30,0,177,0,151,0,209,0,13,0,110,0,49,0,16,0,11,0,54,0,238,0,153,0,51,0,175,0);
signal scenario_full  : scenario_type := (0,0,38,31,243,31,128,31,52,31,191,31,191,30,151,31,195,31,53,31,81,31,236,31,227,31,91,31,108,31,72,31,16,31,142,31,184,31,184,30,226,31,226,30,125,31,125,30,43,31,65,31,80,31,74,31,38,31,75,31,75,30,135,31,194,31,204,31,240,31,155,31,243,31,243,30,2,31,2,30,70,31,37,31,91,31,91,30,115,31,115,30,173,31,145,31,172,31,21,31,187,31,174,31,170,31,58,31,18,31,127,31,102,31,97,31,255,31,18,31,136,31,34,31,69,31,213,31,60,31,137,31,22,31,255,31,232,31,75,31,75,30,217,31,217,30,103,31,87,31,193,31,193,30,237,31,74,31,179,31,116,31,112,31,50,31,23,31,74,31,126,31,124,31,124,30,124,29,50,31,50,30,240,31,22,31,36,31,11,31,2,31,2,30,216,31,216,30,67,31,202,31,184,31,120,31,66,31,1,31,39,31,39,30,18,31,196,31,196,30,12,31,12,30,112,31,254,31,148,31,172,31,135,31,89,31,170,31,43,31,43,30,200,31,225,31,188,31,213,31,53,31,50,31,183,31,7,31,181,31,125,31,200,31,200,30,201,31,43,31,144,31,3,31,116,31,199,31,102,31,130,31,22,31,200,31,62,31,174,31,11,31,50,31,50,30,46,31,57,31,57,30,57,29,57,28,198,31,247,31,255,31,80,31,155,31,15,31,214,31,46,31,111,31,172,31,31,31,112,31,112,30,15,31,182,31,166,31,72,31,229,31,48,31,91,31,150,31,47,31,36,31,36,30,120,31,120,30,120,29,70,31,141,31,238,31,44,31,23,31,136,31,169,31,27,31,245,31,245,30,132,31,119,31,119,30,113,31,185,31,185,30,185,29,56,31,56,30,165,31,24,31,24,30,24,29,24,28,110,31,100,31,1,31,76,31,255,31,118,31,248,31,248,30,221,31,221,30,221,29,48,31,228,31,228,30,231,31,140,31,199,31,169,31,169,30,169,29,10,31,147,31,61,31,128,31,133,31,142,31,112,31,65,31,243,31,99,31,99,30,3,31,3,30,3,29,201,31,215,31,154,31,240,31,141,31,174,31,174,30,15,31,11,31,194,31,194,30,194,29,194,28,194,27,221,31,203,31,243,31,243,30,114,31,150,31,11,31,157,31,180,31,74,31,245,31,55,31,55,30,161,31,161,30,158,31,158,30,158,29,186,31,177,31,156,31,156,30,165,31,30,31,104,31,101,31,101,30,99,31,99,30,225,31,63,31,148,31,44,31,249,31,249,30,5,31,172,31,177,31,251,31,98,31,98,30,186,31,199,31,199,30,79,31,220,31,122,31,121,31,76,31,239,31,92,31,172,31,172,30,32,31,32,30,192,31,15,31,15,30,206,31,22,31,86,31,56,31,227,31,231,31,218,31,50,31,174,31,238,31,197,31,238,31,238,30,186,31,60,31,152,31,171,31,13,31,13,30,176,31,251,31,73,31,135,31,135,30,91,31,13,31,45,31,10,31,196,31,191,31,242,31,55,31,160,31,89,31,237,31,237,30,146,31,146,30,153,31,224,31,254,31,175,31,67,31,67,30,102,31,232,31,232,30,18,31,15,31,211,31,109,31,41,31,191,31,191,30,48,31,48,30,48,29,194,31,12,31,12,30,12,29,83,31,96,31,96,30,96,29,236,31,139,31,6,31,6,30,193,31,57,31,57,30,116,31,5,31,25,31,25,30,17,31,196,31,239,31,239,30,84,31,6,31,195,31,13,31,81,31,23,31,94,31,233,31,236,31,60,31,60,30,74,31,165,31,11,31,11,30,135,31,44,31,98,31,98,30,242,31,87,31,22,31,36,31,57,31,151,31,76,31,76,30,76,29,147,31,166,31,248,31,119,31,8,31,2,31,70,31,45,31,182,31,191,31,203,31,55,31,89,31,103,31,117,31,169,31,169,30,169,29,160,31,12,31,147,31,210,31,222,31,182,31,233,31,78,31,78,30,186,31,186,30,186,29,63,31,47,31,106,31,17,31,110,31,110,30,177,31,60,31,60,30,42,31,180,31,218,31,218,30,13,31,40,31,125,31,17,31,149,31,1,31,41,31,32,31,241,31,216,31,134,31,74,31,46,31,234,31,7,31,64,31,28,31,172,31,115,31,115,30,127,31,96,31,34,31,34,30,43,31,134,31,162,31,245,31,64,31,192,31,82,31,247,31,72,31,64,31,77,31,149,31,78,31,78,30,164,31,164,30,164,29,32,31,32,30,138,31,44,31,37,31,3,31,3,30,169,31,169,30,152,31,67,31,143,31,143,30,109,31,92,31,190,31,190,30,190,29,167,31,118,31,188,31,143,31,210,31,194,31,44,31,44,31,48,31,141,31,119,31,59,31,126,31,21,31,45,31,45,30,163,31,125,31,250,31,47,31,47,30,131,31,230,31,230,30,110,31,43,31,43,30,41,31,207,31,240,31,240,30,20,31,137,31,164,31,145,31,248,31,21,31,100,31,172,31,1,31,246,31,116,31,26,31,139,31,120,31,210,31,210,30,130,31,130,30,17,31,234,31,38,31,4,31,69,31,69,30,76,31,76,30,57,31,92,31,233,31,75,31,60,31,73,31,223,31,69,31,152,31,111,31,135,31,143,31,156,31,54,31,15,31,136,31,148,31,204,31,182,31,19,31,19,30,235,31,170,31,168,31,168,30,168,29,154,31,159,31,81,31,52,31,180,31,186,31,84,31,162,31,251,31,54,31,54,30,54,29,202,31,127,31,241,31,207,31,153,31,161,31,161,30,82,31,154,31,157,31,136,31,224,31,46,31,46,30,46,29,46,28,112,31,112,30,76,31,170,31,236,31,112,31,205,31,92,31,92,30,211,31,95,31,27,31,150,31,63,31,34,31,197,31,81,31,138,31,119,31,75,31,245,31,43,31,45,31,206,31,148,31,66,31,66,30,124,31,170,31,191,31,205,31,46,31,192,31,165,31,165,30,39,31,139,31,66,31,242,31,233,31,169,31,154,31,212,31,212,30,51,31,51,30,3,31,3,30,165,31,165,30,64,31,28,31,165,31,165,30,165,29,165,28,176,31,22,31,15,31,15,30,70,31,70,30,240,31,52,31,52,30,106,31,135,31,135,30,11,31,89,31,89,30,157,31,176,31,221,31,95,31,49,31,76,31,151,31,194,31,128,31,220,31,89,31,99,31,160,31,160,30,160,29,143,31,178,31,99,31,99,30,98,31,108,31,63,31,242,31,125,31,125,30,45,31,146,31,242,31,206,31,245,31,245,30,220,31,68,31,68,30,67,31,210,31,26,31,118,31,118,30,194,31,194,30,111,31,177,31,30,31,177,31,151,31,209,31,13,31,110,31,49,31,16,31,11,31,54,31,238,31,153,31,51,31,175,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
