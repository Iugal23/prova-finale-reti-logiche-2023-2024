-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_579 is
end project_tb_579;

architecture project_tb_arch_579 of project_tb_579 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 809;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,0,0,28,0,214,0,45,0,57,0,144,0,180,0,167,0,0,0,247,0,0,0,199,0,129,0,99,0,185,0,52,0,0,0,180,0,186,0,169,0,175,0,80,0,0,0,67,0,243,0,239,0,223,0,44,0,240,0,122,0,65,0,34,0,40,0,169,0,249,0,108,0,0,0,78,0,17,0,117,0,0,0,94,0,185,0,226,0,201,0,24,0,27,0,210,0,207,0,187,0,0,0,0,0,236,0,0,0,138,0,73,0,142,0,195,0,57,0,111,0,0,0,0,0,66,0,116,0,1,0,84,0,233,0,238,0,146,0,0,0,65,0,211,0,34,0,30,0,0,0,111,0,26,0,0,0,137,0,13,0,152,0,135,0,225,0,194,0,219,0,2,0,116,0,66,0,179,0,214,0,167,0,241,0,185,0,0,0,0,0,0,0,112,0,0,0,49,0,208,0,179,0,0,0,3,0,15,0,211,0,6,0,0,0,179,0,97,0,78,0,0,0,142,0,0,0,203,0,187,0,138,0,131,0,0,0,133,0,246,0,73,0,0,0,192,0,5,0,71,0,146,0,0,0,75,0,43,0,238,0,186,0,181,0,5,0,0,0,27,0,156,0,0,0,149,0,222,0,0,0,230,0,98,0,39,0,83,0,32,0,156,0,0,0,35,0,112,0,201,0,19,0,0,0,247,0,153,0,140,0,168,0,0,0,74,0,203,0,232,0,200,0,54,0,195,0,11,0,0,0,77,0,0,0,170,0,146,0,190,0,235,0,163,0,62,0,0,0,188,0,2,0,156,0,127,0,83,0,162,0,124,0,148,0,102,0,0,0,216,0,87,0,9,0,0,0,0,0,191,0,84,0,66,0,185,0,0,0,219,0,0,0,218,0,20,0,197,0,53,0,193,0,20,0,122,0,0,0,144,0,164,0,63,0,85,0,170,0,119,0,0,0,160,0,14,0,218,0,145,0,251,0,235,0,102,0,163,0,4,0,61,0,188,0,154,0,0,0,0,0,182,0,8,0,116,0,181,0,40,0,0,0,151,0,235,0,183,0,41,0,217,0,92,0,121,0,34,0,161,0,0,0,105,0,0,0,167,0,207,0,183,0,0,0,29,0,154,0,95,0,16,0,0,0,0,0,38,0,66,0,122,0,213,0,100,0,0,0,176,0,0,0,241,0,0,0,26,0,213,0,216,0,0,0,0,0,0,0,253,0,0,0,45,0,152,0,194,0,170,0,70,0,87,0,8,0,179,0,196,0,21,0,121,0,59,0,187,0,47,0,81,0,209,0,20,0,230,0,1,0,19,0,72,0,210,0,165,0,19,0,191,0,158,0,215,0,0,0,0,0,69,0,0,0,0,0,145,0,200,0,13,0,0,0,0,0,188,0,0,0,237,0,0,0,233,0,28,0,0,0,222,0,24,0,79,0,71,0,0,0,0,0,25,0,132,0,71,0,96,0,185,0,203,0,192,0,133,0,67,0,37,0,183,0,147,0,0,0,83,0,0,0,170,0,51,0,0,0,108,0,211,0,237,0,145,0,0,0,79,0,0,0,88,0,94,0,54,0,160,0,120,0,191,0,254,0,68,0,78,0,169,0,0,0,203,0,0,0,125,0,222,0,0,0,152,0,162,0,0,0,234,0,9,0,9,0,0,0,0,0,0,0,0,0,11,0,5,0,194,0,186,0,156,0,55,0,226,0,0,0,244,0,0,0,34,0,0,0,19,0,95,0,0,0,109,0,96,0,153,0,197,0,0,0,246,0,221,0,29,0,104,0,217,0,232,0,250,0,112,0,71,0,0,0,163,0,68,0,164,0,117,0,25,0,241,0,180,0,168,0,195,0,0,0,4,0,130,0,209,0,141,0,185,0,45,0,163,0,0,0,228,0,0,0,12,0,0,0,106,0,0,0,233,0,226,0,150,0,60,0,89,0,233,0,182,0,113,0,201,0,191,0,9,0,163,0,109,0,195,0,122,0,145,0,236,0,56,0,43,0,0,0,60,0,147,0,0,0,14,0,145,0,137,0,0,0,151,0,0,0,152,0,18,0,21,0,138,0,231,0,65,0,85,0,0,0,137,0,0,0,107,0,69,0,227,0,177,0,195,0,249,0,202,0,183,0,166,0,20,0,22,0,243,0,164,0,159,0,199,0,0,0,0,0,223,0,66,0,98,0,38,0,11,0,27,0,62,0,161,0,84,0,245,0,143,0,50,0,63,0,130,0,155,0,0,0,204,0,138,0,166,0,179,0,119,0,0,0,150,0,3,0,10,0,106,0,139,0,54,0,0,0,121,0,117,0,0,0,78,0,112,0,92,0,132,0,201,0,147,0,233,0,233,0,121,0,22,0,65,0,232,0,109,0,0,0,0,0,231,0,120,0,193,0,45,0,197,0,81,0,160,0,0,0,0,0,88,0,229,0,163,0,78,0,0,0,86,0,11,0,218,0,79,0,0,0,0,0,239,0,43,0,0,0,126,0,73,0,251,0,149,0,122,0,230,0,108,0,127,0,7,0,124,0,233,0,0,0,0,0,27,0,179,0,64,0,251,0,0,0,194,0,0,0,24,0,155,0,230,0,28,0,0,0,24,0,205,0,0,0,241,0,71,0,249,0,157,0,4,0,225,0,53,0,217,0,145,0,133,0,0,0,236,0,163,0,249,0,0,0,174,0,246,0,115,0,2,0,2,0,122,0,182,0,0,0,0,0,183,0,158,0,0,0,23,0,101,0,144,0,71,0,13,0,206,0,45,0,0,0,159,0,24,0,140,0,30,0,47,0,137,0,62,0,245,0,132,0,194,0,134,0,220,0,13,0,147,0,0,0,125,0,224,0,226,0,161,0,0,0,119,0,0,0,223,0,22,0,152,0,0,0,67,0,250,0,0,0,0,0,0,0,101,0,89,0,0,0,0,0,35,0,247,0,233,0,0,0,0,0,15,0,48,0,65,0,249,0,190,0,99,0,209,0,50,0,102,0,50,0,112,0,120,0,0,0,47,0,50,0,85,0,0,0,240,0,0,0,200,0,13,0,202,0,209,0,0,0,196,0,203,0,0,0,112,0,156,0,0,0,223,0,0,0,238,0,201,0,241,0,105,0,47,0,0,0,54,0,181,0,84,0,158,0,0,0,71,0,102,0,121,0,184,0,26,0,0,0,60,0,0,0,98,0,0,0,144,0,152,0,124,0,29,0,126,0,64,0,221,0,61,0,239,0,131,0,0,0,191,0,94,0,228,0,10,0,51,0,0,0,0,0,120,0,0,0,3,0,15,0,0,0,32,0,175,0,40,0,0,0,247,0,33,0,14,0,255,0,67,0,100,0,92,0,128,0,0,0,159,0,16,0,150,0,70,0,43,0,108,0,0,0,237,0,232,0,0,0,109,0,134,0,196,0,0,0,0,0,58,0,0,0,80,0,208,0,92,0,0,0,229,0,0,0,98,0,44,0,0,0,0,0,0,0,104,0,150,0,149,0,232,0,183,0,90,0,29,0,155,0,156,0,47,0,36,0,214,0,197,0,37,0,158,0,15,0,43,0,0,0,105,0,90,0,157,0,160,0,234,0,0,0,207,0,105,0,0,0,104,0,159,0,0,0,143,0,253,0,157,0,82,0,185,0);
signal scenario_full  : scenario_type := (0,0,0,0,0,0,28,31,214,31,45,31,57,31,144,31,180,31,167,31,167,30,247,31,247,30,199,31,129,31,99,31,185,31,52,31,52,30,180,31,186,31,169,31,175,31,80,31,80,30,67,31,243,31,239,31,223,31,44,31,240,31,122,31,65,31,34,31,40,31,169,31,249,31,108,31,108,30,78,31,17,31,117,31,117,30,94,31,185,31,226,31,201,31,24,31,27,31,210,31,207,31,187,31,187,30,187,29,236,31,236,30,138,31,73,31,142,31,195,31,57,31,111,31,111,30,111,29,66,31,116,31,1,31,84,31,233,31,238,31,146,31,146,30,65,31,211,31,34,31,30,31,30,30,111,31,26,31,26,30,137,31,13,31,152,31,135,31,225,31,194,31,219,31,2,31,116,31,66,31,179,31,214,31,167,31,241,31,185,31,185,30,185,29,185,28,112,31,112,30,49,31,208,31,179,31,179,30,3,31,15,31,211,31,6,31,6,30,179,31,97,31,78,31,78,30,142,31,142,30,203,31,187,31,138,31,131,31,131,30,133,31,246,31,73,31,73,30,192,31,5,31,71,31,146,31,146,30,75,31,43,31,238,31,186,31,181,31,5,31,5,30,27,31,156,31,156,30,149,31,222,31,222,30,230,31,98,31,39,31,83,31,32,31,156,31,156,30,35,31,112,31,201,31,19,31,19,30,247,31,153,31,140,31,168,31,168,30,74,31,203,31,232,31,200,31,54,31,195,31,11,31,11,30,77,31,77,30,170,31,146,31,190,31,235,31,163,31,62,31,62,30,188,31,2,31,156,31,127,31,83,31,162,31,124,31,148,31,102,31,102,30,216,31,87,31,9,31,9,30,9,29,191,31,84,31,66,31,185,31,185,30,219,31,219,30,218,31,20,31,197,31,53,31,193,31,20,31,122,31,122,30,144,31,164,31,63,31,85,31,170,31,119,31,119,30,160,31,14,31,218,31,145,31,251,31,235,31,102,31,163,31,4,31,61,31,188,31,154,31,154,30,154,29,182,31,8,31,116,31,181,31,40,31,40,30,151,31,235,31,183,31,41,31,217,31,92,31,121,31,34,31,161,31,161,30,105,31,105,30,167,31,207,31,183,31,183,30,29,31,154,31,95,31,16,31,16,30,16,29,38,31,66,31,122,31,213,31,100,31,100,30,176,31,176,30,241,31,241,30,26,31,213,31,216,31,216,30,216,29,216,28,253,31,253,30,45,31,152,31,194,31,170,31,70,31,87,31,8,31,179,31,196,31,21,31,121,31,59,31,187,31,47,31,81,31,209,31,20,31,230,31,1,31,19,31,72,31,210,31,165,31,19,31,191,31,158,31,215,31,215,30,215,29,69,31,69,30,69,29,145,31,200,31,13,31,13,30,13,29,188,31,188,30,237,31,237,30,233,31,28,31,28,30,222,31,24,31,79,31,71,31,71,30,71,29,25,31,132,31,71,31,96,31,185,31,203,31,192,31,133,31,67,31,37,31,183,31,147,31,147,30,83,31,83,30,170,31,51,31,51,30,108,31,211,31,237,31,145,31,145,30,79,31,79,30,88,31,94,31,54,31,160,31,120,31,191,31,254,31,68,31,78,31,169,31,169,30,203,31,203,30,125,31,222,31,222,30,152,31,162,31,162,30,234,31,9,31,9,31,9,30,9,29,9,28,9,27,11,31,5,31,194,31,186,31,156,31,55,31,226,31,226,30,244,31,244,30,34,31,34,30,19,31,95,31,95,30,109,31,96,31,153,31,197,31,197,30,246,31,221,31,29,31,104,31,217,31,232,31,250,31,112,31,71,31,71,30,163,31,68,31,164,31,117,31,25,31,241,31,180,31,168,31,195,31,195,30,4,31,130,31,209,31,141,31,185,31,45,31,163,31,163,30,228,31,228,30,12,31,12,30,106,31,106,30,233,31,226,31,150,31,60,31,89,31,233,31,182,31,113,31,201,31,191,31,9,31,163,31,109,31,195,31,122,31,145,31,236,31,56,31,43,31,43,30,60,31,147,31,147,30,14,31,145,31,137,31,137,30,151,31,151,30,152,31,18,31,21,31,138,31,231,31,65,31,85,31,85,30,137,31,137,30,107,31,69,31,227,31,177,31,195,31,249,31,202,31,183,31,166,31,20,31,22,31,243,31,164,31,159,31,199,31,199,30,199,29,223,31,66,31,98,31,38,31,11,31,27,31,62,31,161,31,84,31,245,31,143,31,50,31,63,31,130,31,155,31,155,30,204,31,138,31,166,31,179,31,119,31,119,30,150,31,3,31,10,31,106,31,139,31,54,31,54,30,121,31,117,31,117,30,78,31,112,31,92,31,132,31,201,31,147,31,233,31,233,31,121,31,22,31,65,31,232,31,109,31,109,30,109,29,231,31,120,31,193,31,45,31,197,31,81,31,160,31,160,30,160,29,88,31,229,31,163,31,78,31,78,30,86,31,11,31,218,31,79,31,79,30,79,29,239,31,43,31,43,30,126,31,73,31,251,31,149,31,122,31,230,31,108,31,127,31,7,31,124,31,233,31,233,30,233,29,27,31,179,31,64,31,251,31,251,30,194,31,194,30,24,31,155,31,230,31,28,31,28,30,24,31,205,31,205,30,241,31,71,31,249,31,157,31,4,31,225,31,53,31,217,31,145,31,133,31,133,30,236,31,163,31,249,31,249,30,174,31,246,31,115,31,2,31,2,31,122,31,182,31,182,30,182,29,183,31,158,31,158,30,23,31,101,31,144,31,71,31,13,31,206,31,45,31,45,30,159,31,24,31,140,31,30,31,47,31,137,31,62,31,245,31,132,31,194,31,134,31,220,31,13,31,147,31,147,30,125,31,224,31,226,31,161,31,161,30,119,31,119,30,223,31,22,31,152,31,152,30,67,31,250,31,250,30,250,29,250,28,101,31,89,31,89,30,89,29,35,31,247,31,233,31,233,30,233,29,15,31,48,31,65,31,249,31,190,31,99,31,209,31,50,31,102,31,50,31,112,31,120,31,120,30,47,31,50,31,85,31,85,30,240,31,240,30,200,31,13,31,202,31,209,31,209,30,196,31,203,31,203,30,112,31,156,31,156,30,223,31,223,30,238,31,201,31,241,31,105,31,47,31,47,30,54,31,181,31,84,31,158,31,158,30,71,31,102,31,121,31,184,31,26,31,26,30,60,31,60,30,98,31,98,30,144,31,152,31,124,31,29,31,126,31,64,31,221,31,61,31,239,31,131,31,131,30,191,31,94,31,228,31,10,31,51,31,51,30,51,29,120,31,120,30,3,31,15,31,15,30,32,31,175,31,40,31,40,30,247,31,33,31,14,31,255,31,67,31,100,31,92,31,128,31,128,30,159,31,16,31,150,31,70,31,43,31,108,31,108,30,237,31,232,31,232,30,109,31,134,31,196,31,196,30,196,29,58,31,58,30,80,31,208,31,92,31,92,30,229,31,229,30,98,31,44,31,44,30,44,29,44,28,104,31,150,31,149,31,232,31,183,31,90,31,29,31,155,31,156,31,47,31,36,31,214,31,197,31,37,31,158,31,15,31,43,31,43,30,105,31,90,31,157,31,160,31,234,31,234,30,207,31,105,31,105,30,104,31,159,31,159,30,143,31,253,31,157,31,82,31,185,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
