-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_31 is
end project_tb_31;

architecture project_tb_arch_31 of project_tb_31 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 355;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (56,0,0,0,33,0,33,0,38,0,45,0,165,0,229,0,83,0,47,0,138,0,0,0,218,0,152,0,90,0,117,0,29,0,0,0,187,0,208,0,252,0,193,0,253,0,244,0,35,0,32,0,57,0,0,0,0,0,0,0,0,0,7,0,24,0,0,0,166,0,0,0,72,0,0,0,134,0,80,0,0,0,205,0,0,0,243,0,0,0,225,0,65,0,253,0,147,0,213,0,0,0,0,0,199,0,0,0,30,0,221,0,28,0,0,0,51,0,68,0,13,0,0,0,173,0,57,0,148,0,118,0,161,0,0,0,47,0,139,0,0,0,167,0,95,0,96,0,0,0,221,0,0,0,254,0,194,0,125,0,8,0,15,0,211,0,161,0,21,0,127,0,211,0,16,0,118,0,0,0,42,0,172,0,140,0,64,0,127,0,227,0,1,0,10,0,64,0,39,0,87,0,149,0,31,0,233,0,105,0,60,0,0,0,187,0,169,0,0,0,129,0,216,0,183,0,0,0,141,0,128,0,161,0,0,0,205,0,0,0,179,0,83,0,15,0,13,0,0,0,245,0,0,0,199,0,0,0,14,0,21,0,52,0,48,0,120,0,69,0,130,0,235,0,91,0,43,0,99,0,168,0,97,0,139,0,179,0,53,0,121,0,0,0,0,0,72,0,0,0,154,0,0,0,226,0,0,0,0,0,0,0,255,0,247,0,72,0,205,0,0,0,103,0,139,0,186,0,240,0,204,0,140,0,0,0,86,0,0,0,46,0,157,0,47,0,42,0,0,0,0,0,157,0,0,0,223,0,194,0,69,0,236,0,175,0,124,0,124,0,170,0,155,0,201,0,240,0,193,0,142,0,158,0,117,0,0,0,177,0,82,0,0,0,36,0,44,0,165,0,31,0,43,0,0,0,170,0,116,0,98,0,172,0,0,0,168,0,58,0,44,0,213,0,155,0,0,0,0,0,133,0,187,0,156,0,0,0,215,0,241,0,226,0,209,0,150,0,254,0,0,0,96,0,123,0,143,0,30,0,169,0,153,0,0,0,217,0,250,0,174,0,228,0,61,0,220,0,65,0,230,0,222,0,12,0,0,0,205,0,0,0,27,0,224,0,254,0,83,0,140,0,93,0,138,0,0,0,97,0,226,0,192,0,1,0,226,0,23,0,0,0,216,0,141,0,204,0,135,0,145,0,169,0,53,0,26,0,206,0,21,0,65,0,0,0,7,0,243,0,225,0,191,0,0,0,0,0,143,0,99,0,79,0,179,0,0,0,0,0,190,0,250,0,131,0,135,0,114,0,197,0,102,0,231,0,0,0,224,0,50,0,0,0,0,0,0,0,0,0,0,0,99,0,0,0,90,0,84,0,190,0,182,0,111,0,41,0,43,0,0,0,24,0,34,0,151,0,0,0,0,0,0,0,17,0,140,0,0,0,64,0,78,0,20,0,197,0,118,0,205,0,0,0,0,0,202,0,52,0,131,0,143,0,0,0,65,0,36,0,152,0,0,0,218,0,151,0,0,0,212,0,0,0,171,0,0,0,181,0,218,0,41,0,171,0,251,0,109,0,0,0,14,0,1,0,0,0,12,0);
signal scenario_full  : scenario_type := (56,31,56,30,33,31,33,31,38,31,45,31,165,31,229,31,83,31,47,31,138,31,138,30,218,31,152,31,90,31,117,31,29,31,29,30,187,31,208,31,252,31,193,31,253,31,244,31,35,31,32,31,57,31,57,30,57,29,57,28,57,27,7,31,24,31,24,30,166,31,166,30,72,31,72,30,134,31,80,31,80,30,205,31,205,30,243,31,243,30,225,31,65,31,253,31,147,31,213,31,213,30,213,29,199,31,199,30,30,31,221,31,28,31,28,30,51,31,68,31,13,31,13,30,173,31,57,31,148,31,118,31,161,31,161,30,47,31,139,31,139,30,167,31,95,31,96,31,96,30,221,31,221,30,254,31,194,31,125,31,8,31,15,31,211,31,161,31,21,31,127,31,211,31,16,31,118,31,118,30,42,31,172,31,140,31,64,31,127,31,227,31,1,31,10,31,64,31,39,31,87,31,149,31,31,31,233,31,105,31,60,31,60,30,187,31,169,31,169,30,129,31,216,31,183,31,183,30,141,31,128,31,161,31,161,30,205,31,205,30,179,31,83,31,15,31,13,31,13,30,245,31,245,30,199,31,199,30,14,31,21,31,52,31,48,31,120,31,69,31,130,31,235,31,91,31,43,31,99,31,168,31,97,31,139,31,179,31,53,31,121,31,121,30,121,29,72,31,72,30,154,31,154,30,226,31,226,30,226,29,226,28,255,31,247,31,72,31,205,31,205,30,103,31,139,31,186,31,240,31,204,31,140,31,140,30,86,31,86,30,46,31,157,31,47,31,42,31,42,30,42,29,157,31,157,30,223,31,194,31,69,31,236,31,175,31,124,31,124,31,170,31,155,31,201,31,240,31,193,31,142,31,158,31,117,31,117,30,177,31,82,31,82,30,36,31,44,31,165,31,31,31,43,31,43,30,170,31,116,31,98,31,172,31,172,30,168,31,58,31,44,31,213,31,155,31,155,30,155,29,133,31,187,31,156,31,156,30,215,31,241,31,226,31,209,31,150,31,254,31,254,30,96,31,123,31,143,31,30,31,169,31,153,31,153,30,217,31,250,31,174,31,228,31,61,31,220,31,65,31,230,31,222,31,12,31,12,30,205,31,205,30,27,31,224,31,254,31,83,31,140,31,93,31,138,31,138,30,97,31,226,31,192,31,1,31,226,31,23,31,23,30,216,31,141,31,204,31,135,31,145,31,169,31,53,31,26,31,206,31,21,31,65,31,65,30,7,31,243,31,225,31,191,31,191,30,191,29,143,31,99,31,79,31,179,31,179,30,179,29,190,31,250,31,131,31,135,31,114,31,197,31,102,31,231,31,231,30,224,31,50,31,50,30,50,29,50,28,50,27,50,26,99,31,99,30,90,31,84,31,190,31,182,31,111,31,41,31,43,31,43,30,24,31,34,31,151,31,151,30,151,29,151,28,17,31,140,31,140,30,64,31,78,31,20,31,197,31,118,31,205,31,205,30,205,29,202,31,52,31,131,31,143,31,143,30,65,31,36,31,152,31,152,30,218,31,151,31,151,30,212,31,212,30,171,31,171,30,181,31,218,31,41,31,171,31,251,31,109,31,109,30,14,31,1,31,1,30,12,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
