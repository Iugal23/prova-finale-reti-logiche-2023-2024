-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_454 is
end project_tb_454;

architecture project_tb_arch_454 of project_tb_454 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 833;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (64,0,123,0,122,0,188,0,0,0,106,0,193,0,0,0,214,0,209,0,170,0,0,0,235,0,57,0,0,0,35,0,29,0,64,0,59,0,254,0,244,0,136,0,209,0,224,0,247,0,0,0,0,0,112,0,0,0,0,0,155,0,0,0,10,0,200,0,242,0,210,0,231,0,0,0,78,0,221,0,221,0,118,0,24,0,33,0,123,0,38,0,136,0,136,0,217,0,0,0,125,0,0,0,233,0,54,0,176,0,116,0,192,0,190,0,9,0,127,0,89,0,186,0,0,0,0,0,0,0,138,0,246,0,208,0,240,0,149,0,0,0,101,0,0,0,150,0,0,0,15,0,164,0,198,0,0,0,166,0,129,0,231,0,79,0,34,0,198,0,205,0,230,0,147,0,252,0,0,0,125,0,148,0,184,0,0,0,193,0,15,0,3,0,28,0,175,0,0,0,117,0,187,0,210,0,83,0,30,0,0,0,209,0,171,0,62,0,60,0,239,0,220,0,66,0,93,0,163,0,30,0,19,0,101,0,0,0,238,0,145,0,149,0,0,0,134,0,10,0,176,0,124,0,162,0,0,0,219,0,85,0,30,0,127,0,0,0,73,0,0,0,62,0,157,0,0,0,228,0,224,0,0,0,181,0,65,0,75,0,192,0,84,0,185,0,222,0,37,0,74,0,198,0,69,0,241,0,232,0,83,0,0,0,191,0,220,0,230,0,103,0,168,0,41,0,0,0,184,0,222,0,0,0,0,0,187,0,234,0,181,0,91,0,13,0,198,0,114,0,0,0,166,0,161,0,240,0,226,0,221,0,191,0,159,0,20,0,214,0,0,0,234,0,154,0,84,0,45,0,124,0,69,0,20,0,61,0,35,0,126,0,0,0,182,0,7,0,254,0,66,0,162,0,32,0,182,0,183,0,51,0,170,0,0,0,111,0,0,0,0,0,44,0,139,0,243,0,186,0,22,0,0,0,243,0,34,0,45,0,166,0,100,0,134,0,173,0,0,0,0,0,228,0,240,0,203,0,73,0,176,0,58,0,220,0,60,0,181,0,178,0,224,0,0,0,0,0,87,0,169,0,93,0,0,0,206,0,0,0,30,0,38,0,138,0,229,0,223,0,0,0,240,0,46,0,252,0,207,0,219,0,0,0,0,0,190,0,0,0,194,0,134,0,227,0,0,0,0,0,38,0,150,0,39,0,219,0,208,0,0,0,0,0,140,0,0,0,114,0,236,0,179,0,4,0,18,0,0,0,169,0,194,0,79,0,246,0,99,0,83,0,33,0,17,0,76,0,54,0,17,0,28,0,0,0,192,0,166,0,133,0,0,0,153,0,61,0,0,0,122,0,33,0,35,0,129,0,113,0,0,0,163,0,53,0,187,0,0,0,0,0,171,0,81,0,201,0,118,0,254,0,0,0,235,0,56,0,0,0,12,0,102,0,53,0,27,0,70,0,138,0,16,0,0,0,0,0,87,0,248,0,134,0,147,0,234,0,30,0,0,0,156,0,23,0,163,0,24,0,6,0,79,0,171,0,42,0,156,0,159,0,202,0,74,0,0,0,159,0,120,0,168,0,87,0,127,0,0,0,9,0,0,0,143,0,0,0,88,0,169,0,246,0,133,0,243,0,215,0,74,0,90,0,71,0,81,0,0,0,112,0,0,0,0,0,249,0,75,0,175,0,59,0,121,0,0,0,243,0,0,0,172,0,172,0,44,0,187,0,235,0,0,0,44,0,225,0,85,0,159,0,252,0,20,0,0,0,94,0,0,0,61,0,84,0,228,0,89,0,0,0,0,0,92,0,113,0,24,0,107,0,56,0,79,0,6,0,68,0,0,0,104,0,190,0,0,0,59,0,153,0,73,0,97,0,0,0,233,0,53,0,241,0,0,0,18,0,42,0,7,0,218,0,8,0,0,0,84,0,142,0,158,0,0,0,211,0,84,0,54,0,254,0,70,0,93,0,169,0,58,0,107,0,44,0,132,0,71,0,0,0,167,0,241,0,135,0,156,0,253,0,51,0,140,0,200,0,205,0,217,0,82,0,216,0,227,0,54,0,94,0,120,0,22,0,82,0,185,0,102,0,117,0,0,0,99,0,6,0,111,0,22,0,174,0,142,0,101,0,131,0,70,0,65,0,59,0,245,0,236,0,154,0,126,0,164,0,81,0,42,0,0,0,244,0,136,0,22,0,68,0,19,0,0,0,57,0,0,0,41,0,0,0,47,0,7,0,0,0,116,0,0,0,106,0,145,0,210,0,153,0,101,0,60,0,240,0,80,0,124,0,163,0,162,0,189,0,0,0,70,0,95,0,155,0,0,0,167,0,30,0,63,0,203,0,82,0,200,0,1,0,205,0,96,0,0,0,231,0,185,0,136,0,193,0,0,0,34,0,0,0,74,0,229,0,154,0,0,0,0,0,0,0,0,0,66,0,46,0,0,0,12,0,0,0,0,0,3,0,93,0,179,0,48,0,0,0,148,0,106,0,145,0,17,0,0,0,133,0,68,0,0,0,24,0,162,0,195,0,169,0,193,0,9,0,47,0,56,0,203,0,84,0,134,0,51,0,216,0,44,0,158,0,242,0,208,0,82,0,58,0,41,0,180,0,205,0,247,0,175,0,0,0,159,0,235,0,149,0,0,0,118,0,199,0,191,0,220,0,96,0,135,0,56,0,4,0,139,0,26,0,19,0,73,0,115,0,226,0,152,0,122,0,243,0,21,0,118,0,181,0,203,0,0,0,148,0,212,0,201,0,71,0,67,0,5,0,201,0,0,0,0,0,196,0,180,0,176,0,228,0,198,0,76,0,235,0,45,0,24,0,0,0,96,0,249,0,204,0,192,0,102,0,0,0,99,0,0,0,1,0,0,0,219,0,168,0,232,0,133,0,138,0,0,0,217,0,238,0,236,0,118,0,12,0,89,0,155,0,92,0,155,0,80,0,0,0,216,0,223,0,0,0,0,0,152,0,226,0,236,0,159,0,176,0,0,0,194,0,210,0,180,0,71,0,115,0,0,0,102,0,81,0,63,0,165,0,55,0,144,0,25,0,0,0,0,0,76,0,42,0,138,0,234,0,204,0,0,0,0,0,178,0,27,0,14,0,83,0,41,0,156,0,170,0,230,0,235,0,82,0,250,0,68,0,170,0,0,0,177,0,0,0,254,0,16,0,98,0,168,0,8,0,115,0,107,0,57,0,82,0,214,0,0,0,224,0,0,0,167,0,154,0,92,0,0,0,205,0,34,0,216,0,153,0,54,0,19,0,132,0,154,0,0,0,65,0,23,0,231,0,249,0,171,0,180,0,144,0,54,0,95,0,104,0,211,0,0,0,0,0,0,0,35,0,165,0,153,0,194,0,123,0,102,0,19,0,118,0,114,0,162,0,0,0,81,0,49,0,190,0,200,0,140,0,46,0,20,0,54,0,0,0,22,0,220,0,11,0,205,0,250,0,100,0,125,0,0,0,29,0,0,0,204,0,128,0,23,0,138,0,0,0,0,0,229,0,0,0,215,0,61,0,180,0,36,0,206,0,68,0,152,0,0,0,0,0,0,0,0,0,36,0,0,0,0,0,0,0,182,0,0,0,124,0,73,0,71,0,172,0,174,0,74,0,0,0,0,0,0,0,147,0,0,0,249,0,219,0,107,0,143,0,123,0,169,0,76,0,220,0,12,0,177,0,60,0,23,0,50,0,177,0,0,0,43,0,0,0,0,0,17,0,0,0);
signal scenario_full  : scenario_type := (64,31,123,31,122,31,188,31,188,30,106,31,193,31,193,30,214,31,209,31,170,31,170,30,235,31,57,31,57,30,35,31,29,31,64,31,59,31,254,31,244,31,136,31,209,31,224,31,247,31,247,30,247,29,112,31,112,30,112,29,155,31,155,30,10,31,200,31,242,31,210,31,231,31,231,30,78,31,221,31,221,31,118,31,24,31,33,31,123,31,38,31,136,31,136,31,217,31,217,30,125,31,125,30,233,31,54,31,176,31,116,31,192,31,190,31,9,31,127,31,89,31,186,31,186,30,186,29,186,28,138,31,246,31,208,31,240,31,149,31,149,30,101,31,101,30,150,31,150,30,15,31,164,31,198,31,198,30,166,31,129,31,231,31,79,31,34,31,198,31,205,31,230,31,147,31,252,31,252,30,125,31,148,31,184,31,184,30,193,31,15,31,3,31,28,31,175,31,175,30,117,31,187,31,210,31,83,31,30,31,30,30,209,31,171,31,62,31,60,31,239,31,220,31,66,31,93,31,163,31,30,31,19,31,101,31,101,30,238,31,145,31,149,31,149,30,134,31,10,31,176,31,124,31,162,31,162,30,219,31,85,31,30,31,127,31,127,30,73,31,73,30,62,31,157,31,157,30,228,31,224,31,224,30,181,31,65,31,75,31,192,31,84,31,185,31,222,31,37,31,74,31,198,31,69,31,241,31,232,31,83,31,83,30,191,31,220,31,230,31,103,31,168,31,41,31,41,30,184,31,222,31,222,30,222,29,187,31,234,31,181,31,91,31,13,31,198,31,114,31,114,30,166,31,161,31,240,31,226,31,221,31,191,31,159,31,20,31,214,31,214,30,234,31,154,31,84,31,45,31,124,31,69,31,20,31,61,31,35,31,126,31,126,30,182,31,7,31,254,31,66,31,162,31,32,31,182,31,183,31,51,31,170,31,170,30,111,31,111,30,111,29,44,31,139,31,243,31,186,31,22,31,22,30,243,31,34,31,45,31,166,31,100,31,134,31,173,31,173,30,173,29,228,31,240,31,203,31,73,31,176,31,58,31,220,31,60,31,181,31,178,31,224,31,224,30,224,29,87,31,169,31,93,31,93,30,206,31,206,30,30,31,38,31,138,31,229,31,223,31,223,30,240,31,46,31,252,31,207,31,219,31,219,30,219,29,190,31,190,30,194,31,134,31,227,31,227,30,227,29,38,31,150,31,39,31,219,31,208,31,208,30,208,29,140,31,140,30,114,31,236,31,179,31,4,31,18,31,18,30,169,31,194,31,79,31,246,31,99,31,83,31,33,31,17,31,76,31,54,31,17,31,28,31,28,30,192,31,166,31,133,31,133,30,153,31,61,31,61,30,122,31,33,31,35,31,129,31,113,31,113,30,163,31,53,31,187,31,187,30,187,29,171,31,81,31,201,31,118,31,254,31,254,30,235,31,56,31,56,30,12,31,102,31,53,31,27,31,70,31,138,31,16,31,16,30,16,29,87,31,248,31,134,31,147,31,234,31,30,31,30,30,156,31,23,31,163,31,24,31,6,31,79,31,171,31,42,31,156,31,159,31,202,31,74,31,74,30,159,31,120,31,168,31,87,31,127,31,127,30,9,31,9,30,143,31,143,30,88,31,169,31,246,31,133,31,243,31,215,31,74,31,90,31,71,31,81,31,81,30,112,31,112,30,112,29,249,31,75,31,175,31,59,31,121,31,121,30,243,31,243,30,172,31,172,31,44,31,187,31,235,31,235,30,44,31,225,31,85,31,159,31,252,31,20,31,20,30,94,31,94,30,61,31,84,31,228,31,89,31,89,30,89,29,92,31,113,31,24,31,107,31,56,31,79,31,6,31,68,31,68,30,104,31,190,31,190,30,59,31,153,31,73,31,97,31,97,30,233,31,53,31,241,31,241,30,18,31,42,31,7,31,218,31,8,31,8,30,84,31,142,31,158,31,158,30,211,31,84,31,54,31,254,31,70,31,93,31,169,31,58,31,107,31,44,31,132,31,71,31,71,30,167,31,241,31,135,31,156,31,253,31,51,31,140,31,200,31,205,31,217,31,82,31,216,31,227,31,54,31,94,31,120,31,22,31,82,31,185,31,102,31,117,31,117,30,99,31,6,31,111,31,22,31,174,31,142,31,101,31,131,31,70,31,65,31,59,31,245,31,236,31,154,31,126,31,164,31,81,31,42,31,42,30,244,31,136,31,22,31,68,31,19,31,19,30,57,31,57,30,41,31,41,30,47,31,7,31,7,30,116,31,116,30,106,31,145,31,210,31,153,31,101,31,60,31,240,31,80,31,124,31,163,31,162,31,189,31,189,30,70,31,95,31,155,31,155,30,167,31,30,31,63,31,203,31,82,31,200,31,1,31,205,31,96,31,96,30,231,31,185,31,136,31,193,31,193,30,34,31,34,30,74,31,229,31,154,31,154,30,154,29,154,28,154,27,66,31,46,31,46,30,12,31,12,30,12,29,3,31,93,31,179,31,48,31,48,30,148,31,106,31,145,31,17,31,17,30,133,31,68,31,68,30,24,31,162,31,195,31,169,31,193,31,9,31,47,31,56,31,203,31,84,31,134,31,51,31,216,31,44,31,158,31,242,31,208,31,82,31,58,31,41,31,180,31,205,31,247,31,175,31,175,30,159,31,235,31,149,31,149,30,118,31,199,31,191,31,220,31,96,31,135,31,56,31,4,31,139,31,26,31,19,31,73,31,115,31,226,31,152,31,122,31,243,31,21,31,118,31,181,31,203,31,203,30,148,31,212,31,201,31,71,31,67,31,5,31,201,31,201,30,201,29,196,31,180,31,176,31,228,31,198,31,76,31,235,31,45,31,24,31,24,30,96,31,249,31,204,31,192,31,102,31,102,30,99,31,99,30,1,31,1,30,219,31,168,31,232,31,133,31,138,31,138,30,217,31,238,31,236,31,118,31,12,31,89,31,155,31,92,31,155,31,80,31,80,30,216,31,223,31,223,30,223,29,152,31,226,31,236,31,159,31,176,31,176,30,194,31,210,31,180,31,71,31,115,31,115,30,102,31,81,31,63,31,165,31,55,31,144,31,25,31,25,30,25,29,76,31,42,31,138,31,234,31,204,31,204,30,204,29,178,31,27,31,14,31,83,31,41,31,156,31,170,31,230,31,235,31,82,31,250,31,68,31,170,31,170,30,177,31,177,30,254,31,16,31,98,31,168,31,8,31,115,31,107,31,57,31,82,31,214,31,214,30,224,31,224,30,167,31,154,31,92,31,92,30,205,31,34,31,216,31,153,31,54,31,19,31,132,31,154,31,154,30,65,31,23,31,231,31,249,31,171,31,180,31,144,31,54,31,95,31,104,31,211,31,211,30,211,29,211,28,35,31,165,31,153,31,194,31,123,31,102,31,19,31,118,31,114,31,162,31,162,30,81,31,49,31,190,31,200,31,140,31,46,31,20,31,54,31,54,30,22,31,220,31,11,31,205,31,250,31,100,31,125,31,125,30,29,31,29,30,204,31,128,31,23,31,138,31,138,30,138,29,229,31,229,30,215,31,61,31,180,31,36,31,206,31,68,31,152,31,152,30,152,29,152,28,152,27,36,31,36,30,36,29,36,28,182,31,182,30,124,31,73,31,71,31,172,31,174,31,74,31,74,30,74,29,74,28,147,31,147,30,249,31,219,31,107,31,143,31,123,31,169,31,76,31,220,31,12,31,177,31,60,31,23,31,50,31,177,31,177,30,43,31,43,30,43,29,17,31,17,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
