-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_317 is
end project_tb_317;

architecture project_tb_arch_317 of project_tb_317 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 291;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (158,0,189,0,43,0,47,0,135,0,3,0,249,0,0,0,181,0,43,0,83,0,52,0,28,0,206,0,0,0,253,0,0,0,0,0,253,0,146,0,150,0,0,0,163,0,76,0,151,0,42,0,255,0,0,0,242,0,54,0,0,0,244,0,168,0,234,0,0,0,125,0,0,0,184,0,118,0,0,0,239,0,0,0,138,0,210,0,0,0,175,0,134,0,23,0,155,0,0,0,165,0,0,0,0,0,120,0,65,0,198,0,84,0,0,0,68,0,0,0,12,0,22,0,162,0,45,0,189,0,0,0,1,0,0,0,0,0,184,0,202,0,60,0,162,0,0,0,65,0,34,0,229,0,0,0,0,0,0,0,125,0,1,0,28,0,25,0,141,0,122,0,19,0,89,0,8,0,110,0,174,0,234,0,19,0,0,0,0,0,221,0,84,0,32,0,9,0,13,0,124,0,6,0,153,0,103,0,0,0,214,0,209,0,17,0,240,0,114,0,223,0,223,0,98,0,103,0,117,0,0,0,178,0,0,0,251,0,140,0,0,0,210,0,88,0,0,0,18,0,0,0,21,0,195,0,0,0,214,0,220,0,136,0,249,0,198,0,234,0,171,0,152,0,65,0,28,0,157,0,0,0,81,0,236,0,231,0,234,0,0,0,100,0,95,0,0,0,169,0,106,0,63,0,43,0,8,0,79,0,178,0,0,0,244,0,0,0,0,0,0,0,4,0,0,0,141,0,20,0,77,0,0,0,120,0,200,0,78,0,131,0,163,0,37,0,191,0,59,0,153,0,216,0,200,0,173,0,0,0,142,0,97,0,94,0,116,0,189,0,153,0,0,0,0,0,154,0,185,0,57,0,158,0,231,0,137,0,25,0,136,0,72,0,22,0,36,0,37,0,57,0,0,0,53,0,16,0,95,0,190,0,227,0,250,0,0,0,117,0,254,0,143,0,29,0,121,0,173,0,175,0,0,0,171,0,131,0,192,0,101,0,243,0,26,0,129,0,0,0,2,0,149,0,87,0,0,0,185,0,24,0,126,0,37,0,206,0,250,0,202,0,162,0,217,0,77,0,254,0,71,0,0,0,253,0,147,0,69,0,144,0,0,0,0,0,0,0,119,0,0,0,0,0,77,0,33,0,75,0,0,0,106,0,107,0,23,0,208,0,83,0,95,0,145,0,0,0,0,0,50,0,0,0,126,0,110,0,0,0,23,0,108,0,188,0,0,0,0,0,48,0,0,0,187,0,0,0,97,0,227,0,113,0,0,0,206,0,0,0,0,0,117,0,0,0,0,0,114,0,0,0);
signal scenario_full  : scenario_type := (158,31,189,31,43,31,47,31,135,31,3,31,249,31,249,30,181,31,43,31,83,31,52,31,28,31,206,31,206,30,253,31,253,30,253,29,253,31,146,31,150,31,150,30,163,31,76,31,151,31,42,31,255,31,255,30,242,31,54,31,54,30,244,31,168,31,234,31,234,30,125,31,125,30,184,31,118,31,118,30,239,31,239,30,138,31,210,31,210,30,175,31,134,31,23,31,155,31,155,30,165,31,165,30,165,29,120,31,65,31,198,31,84,31,84,30,68,31,68,30,12,31,22,31,162,31,45,31,189,31,189,30,1,31,1,30,1,29,184,31,202,31,60,31,162,31,162,30,65,31,34,31,229,31,229,30,229,29,229,28,125,31,1,31,28,31,25,31,141,31,122,31,19,31,89,31,8,31,110,31,174,31,234,31,19,31,19,30,19,29,221,31,84,31,32,31,9,31,13,31,124,31,6,31,153,31,103,31,103,30,214,31,209,31,17,31,240,31,114,31,223,31,223,31,98,31,103,31,117,31,117,30,178,31,178,30,251,31,140,31,140,30,210,31,88,31,88,30,18,31,18,30,21,31,195,31,195,30,214,31,220,31,136,31,249,31,198,31,234,31,171,31,152,31,65,31,28,31,157,31,157,30,81,31,236,31,231,31,234,31,234,30,100,31,95,31,95,30,169,31,106,31,63,31,43,31,8,31,79,31,178,31,178,30,244,31,244,30,244,29,244,28,4,31,4,30,141,31,20,31,77,31,77,30,120,31,200,31,78,31,131,31,163,31,37,31,191,31,59,31,153,31,216,31,200,31,173,31,173,30,142,31,97,31,94,31,116,31,189,31,153,31,153,30,153,29,154,31,185,31,57,31,158,31,231,31,137,31,25,31,136,31,72,31,22,31,36,31,37,31,57,31,57,30,53,31,16,31,95,31,190,31,227,31,250,31,250,30,117,31,254,31,143,31,29,31,121,31,173,31,175,31,175,30,171,31,131,31,192,31,101,31,243,31,26,31,129,31,129,30,2,31,149,31,87,31,87,30,185,31,24,31,126,31,37,31,206,31,250,31,202,31,162,31,217,31,77,31,254,31,71,31,71,30,253,31,147,31,69,31,144,31,144,30,144,29,144,28,119,31,119,30,119,29,77,31,33,31,75,31,75,30,106,31,107,31,23,31,208,31,83,31,95,31,145,31,145,30,145,29,50,31,50,30,126,31,110,31,110,30,23,31,108,31,188,31,188,30,188,29,48,31,48,30,187,31,187,30,97,31,227,31,113,31,113,30,206,31,206,30,206,29,117,31,117,30,117,29,114,31,114,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
