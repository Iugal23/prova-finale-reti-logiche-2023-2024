-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_35 is
end project_tb_35;

architecture project_tb_arch_35 of project_tb_35 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 791;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (234,0,137,0,226,0,61,0,143,0,0,0,202,0,106,0,50,0,0,0,79,0,0,0,229,0,128,0,0,0,0,0,135,0,0,0,0,0,191,0,96,0,196,0,9,0,239,0,205,0,26,0,164,0,159,0,115,0,83,0,0,0,108,0,51,0,0,0,118,0,221,0,119,0,227,0,88,0,0,0,37,0,226,0,27,0,79,0,61,0,135,0,72,0,0,0,159,0,0,0,213,0,0,0,20,0,0,0,199,0,37,0,95,0,237,0,37,0,244,0,157,0,21,0,30,0,20,0,24,0,81,0,0,0,4,0,230,0,246,0,108,0,66,0,137,0,237,0,84,0,45,0,38,0,0,0,119,0,5,0,1,0,0,0,0,0,211,0,55,0,0,0,136,0,113,0,0,0,158,0,1,0,168,0,199,0,133,0,0,0,74,0,142,0,177,0,140,0,246,0,163,0,82,0,169,0,224,0,222,0,0,0,95,0,0,0,77,0,189,0,0,0,60,0,192,0,20,0,0,0,35,0,79,0,161,0,235,0,0,0,250,0,61,0,156,0,38,0,49,0,149,0,150,0,241,0,0,0,0,0,197,0,212,0,186,0,183,0,169,0,104,0,17,0,109,0,0,0,134,0,170,0,44,0,152,0,180,0,0,0,201,0,128,0,96,0,166,0,152,0,224,0,71,0,193,0,101,0,0,0,165,0,235,0,179,0,120,0,183,0,61,0,64,0,233,0,23,0,27,0,47,0,35,0,19,0,21,0,117,0,89,0,124,0,181,0,176,0,12,0,0,0,0,0,0,0,48,0,59,0,37,0,242,0,0,0,101,0,37,0,33,0,214,0,0,0,167,0,0,0,168,0,49,0,255,0,0,0,222,0,42,0,116,0,136,0,0,0,230,0,176,0,229,0,89,0,231,0,97,0,0,0,0,0,0,0,241,0,0,0,214,0,79,0,205,0,136,0,209,0,173,0,0,0,213,0,0,0,1,0,254,0,170,0,0,0,182,0,163,0,190,0,72,0,240,0,220,0,79,0,0,0,0,0,141,0,0,0,226,0,158,0,13,0,28,0,72,0,189,0,182,0,219,0,191,0,76,0,103,0,121,0,215,0,101,0,222,0,0,0,149,0,59,0,41,0,244,0,0,0,34,0,24,0,178,0,112,0,204,0,163,0,198,0,112,0,44,0,131,0,136,0,255,0,146,0,210,0,242,0,193,0,63,0,0,0,91,0,27,0,15,0,0,0,189,0,147,0,2,0,104,0,0,0,45,0,193,0,119,0,179,0,172,0,111,0,240,0,132,0,234,0,247,0,0,0,136,0,73,0,0,0,0,0,0,0,195,0,124,0,87,0,27,0,212,0,72,0,254,0,26,0,137,0,250,0,216,0,218,0,0,0,32,0,214,0,248,0,115,0,0,0,221,0,104,0,0,0,21,0,140,0,240,0,113,0,0,0,0,0,117,0,0,0,192,0,0,0,79,0,67,0,0,0,163,0,170,0,31,0,226,0,232,0,236,0,0,0,78,0,8,0,8,0,0,0,234,0,36,0,231,0,153,0,0,0,0,0,51,0,88,0,84,0,31,0,0,0,245,0,249,0,63,0,224,0,203,0,218,0,63,0,0,0,85,0,170,0,196,0,123,0,0,0,103,0,0,0,41,0,0,0,0,0,0,0,124,0,113,0,0,0,69,0,112,0,226,0,0,0,125,0,0,0,224,0,139,0,0,0,241,0,243,0,79,0,205,0,0,0,0,0,196,0,189,0,0,0,61,0,132,0,13,0,0,0,0,0,82,0,241,0,195,0,110,0,122,0,113,0,134,0,208,0,43,0,94,0,123,0,222,0,138,0,117,0,44,0,228,0,209,0,83,0,0,0,0,0,57,0,48,0,0,0,232,0,96,0,32,0,103,0,22,0,196,0,244,0,239,0,246,0,0,0,164,0,179,0,0,0,44,0,184,0,137,0,131,0,74,0,61,0,0,0,37,0,0,0,0,0,34,0,0,0,200,0,240,0,151,0,23,0,108,0,229,0,68,0,173,0,53,0,3,0,65,0,0,0,0,0,0,0,96,0,154,0,243,0,138,0,29,0,36,0,157,0,85,0,220,0,85,0,90,0,114,0,111,0,245,0,151,0,0,0,247,0,9,0,90,0,78,0,84,0,71,0,73,0,7,0,0,0,165,0,33,0,72,0,0,0,166,0,25,0,239,0,83,0,0,0,174,0,0,0,90,0,216,0,75,0,0,0,0,0,0,0,148,0,72,0,240,0,15,0,0,0,156,0,130,0,16,0,14,0,198,0,137,0,0,0,212,0,122,0,60,0,198,0,176,0,127,0,0,0,0,0,233,0,190,0,81,0,181,0,131,0,244,0,58,0,167,0,0,0,0,0,216,0,25,0,220,0,0,0,0,0,23,0,169,0,202,0,164,0,83,0,0,0,125,0,0,0,116,0,229,0,0,0,155,0,189,0,8,0,0,0,103,0,172,0,211,0,186,0,13,0,62,0,234,0,114,0,193,0,178,0,132,0,0,0,97,0,201,0,180,0,121,0,194,0,219,0,20,0,141,0,0,0,56,0,221,0,38,0,38,0,0,0,196,0,0,0,181,0,0,0,0,0,49,0,2,0,120,0,0,0,225,0,106,0,217,0,45,0,210,0,156,0,162,0,176,0,213,0,35,0,96,0,155,0,172,0,0,0,0,0,156,0,193,0,43,0,102,0,0,0,0,0,64,0,0,0,118,0,0,0,237,0,126,0,195,0,57,0,98,0,0,0,122,0,0,0,222,0,179,0,148,0,94,0,0,0,113,0,148,0,0,0,151,0,232,0,239,0,212,0,102,0,207,0,116,0,221,0,67,0,147,0,176,0,248,0,0,0,207,0,224,0,24,0,105,0,0,0,8,0,174,0,67,0,249,0,0,0,217,0,251,0,0,0,115,0,51,0,140,0,161,0,136,0,105,0,125,0,155,0,174,0,18,0,114,0,0,0,246,0,0,0,18,0,206,0,251,0,237,0,0,0,165,0,95,0,86,0,0,0,103,0,176,0,0,0,1,0,207,0,122,0,112,0,102,0,0,0,242,0,199,0,91,0,0,0,146,0,67,0,252,0,222,0,144,0,0,0,100,0,176,0,224,0,212,0,50,0,240,0,216,0,0,0,214,0,103,0,166,0,246,0,0,0,67,0,62,0,17,0,0,0,121,0,172,0,141,0,0,0,201,0,117,0,254,0,13,0,213,0,152,0,124,0,147,0,73,0,189,0,50,0,167,0,193,0,13,0,211,0,0,0,0,0,85,0,0,0,113,0,27,0,120,0,0,0,36,0,0,0,166,0,251,0,217,0,241,0,111,0,125,0,0,0,0,0,47,0,114,0,49,0,126,0,188,0,100,0,115,0,242,0,15,0,0,0,0,0,144,0,0,0,23,0,0,0,0,0,169,0,33,0,143,0,138,0,0,0,237,0,0,0,0,0,217,0,20,0,44,0,225,0,65,0,47,0,124,0,181,0,0,0,0,0,55,0,0,0,1,0,35,0,161,0,46,0);
signal scenario_full  : scenario_type := (234,31,137,31,226,31,61,31,143,31,143,30,202,31,106,31,50,31,50,30,79,31,79,30,229,31,128,31,128,30,128,29,135,31,135,30,135,29,191,31,96,31,196,31,9,31,239,31,205,31,26,31,164,31,159,31,115,31,83,31,83,30,108,31,51,31,51,30,118,31,221,31,119,31,227,31,88,31,88,30,37,31,226,31,27,31,79,31,61,31,135,31,72,31,72,30,159,31,159,30,213,31,213,30,20,31,20,30,199,31,37,31,95,31,237,31,37,31,244,31,157,31,21,31,30,31,20,31,24,31,81,31,81,30,4,31,230,31,246,31,108,31,66,31,137,31,237,31,84,31,45,31,38,31,38,30,119,31,5,31,1,31,1,30,1,29,211,31,55,31,55,30,136,31,113,31,113,30,158,31,1,31,168,31,199,31,133,31,133,30,74,31,142,31,177,31,140,31,246,31,163,31,82,31,169,31,224,31,222,31,222,30,95,31,95,30,77,31,189,31,189,30,60,31,192,31,20,31,20,30,35,31,79,31,161,31,235,31,235,30,250,31,61,31,156,31,38,31,49,31,149,31,150,31,241,31,241,30,241,29,197,31,212,31,186,31,183,31,169,31,104,31,17,31,109,31,109,30,134,31,170,31,44,31,152,31,180,31,180,30,201,31,128,31,96,31,166,31,152,31,224,31,71,31,193,31,101,31,101,30,165,31,235,31,179,31,120,31,183,31,61,31,64,31,233,31,23,31,27,31,47,31,35,31,19,31,21,31,117,31,89,31,124,31,181,31,176,31,12,31,12,30,12,29,12,28,48,31,59,31,37,31,242,31,242,30,101,31,37,31,33,31,214,31,214,30,167,31,167,30,168,31,49,31,255,31,255,30,222,31,42,31,116,31,136,31,136,30,230,31,176,31,229,31,89,31,231,31,97,31,97,30,97,29,97,28,241,31,241,30,214,31,79,31,205,31,136,31,209,31,173,31,173,30,213,31,213,30,1,31,254,31,170,31,170,30,182,31,163,31,190,31,72,31,240,31,220,31,79,31,79,30,79,29,141,31,141,30,226,31,158,31,13,31,28,31,72,31,189,31,182,31,219,31,191,31,76,31,103,31,121,31,215,31,101,31,222,31,222,30,149,31,59,31,41,31,244,31,244,30,34,31,24,31,178,31,112,31,204,31,163,31,198,31,112,31,44,31,131,31,136,31,255,31,146,31,210,31,242,31,193,31,63,31,63,30,91,31,27,31,15,31,15,30,189,31,147,31,2,31,104,31,104,30,45,31,193,31,119,31,179,31,172,31,111,31,240,31,132,31,234,31,247,31,247,30,136,31,73,31,73,30,73,29,73,28,195,31,124,31,87,31,27,31,212,31,72,31,254,31,26,31,137,31,250,31,216,31,218,31,218,30,32,31,214,31,248,31,115,31,115,30,221,31,104,31,104,30,21,31,140,31,240,31,113,31,113,30,113,29,117,31,117,30,192,31,192,30,79,31,67,31,67,30,163,31,170,31,31,31,226,31,232,31,236,31,236,30,78,31,8,31,8,31,8,30,234,31,36,31,231,31,153,31,153,30,153,29,51,31,88,31,84,31,31,31,31,30,245,31,249,31,63,31,224,31,203,31,218,31,63,31,63,30,85,31,170,31,196,31,123,31,123,30,103,31,103,30,41,31,41,30,41,29,41,28,124,31,113,31,113,30,69,31,112,31,226,31,226,30,125,31,125,30,224,31,139,31,139,30,241,31,243,31,79,31,205,31,205,30,205,29,196,31,189,31,189,30,61,31,132,31,13,31,13,30,13,29,82,31,241,31,195,31,110,31,122,31,113,31,134,31,208,31,43,31,94,31,123,31,222,31,138,31,117,31,44,31,228,31,209,31,83,31,83,30,83,29,57,31,48,31,48,30,232,31,96,31,32,31,103,31,22,31,196,31,244,31,239,31,246,31,246,30,164,31,179,31,179,30,44,31,184,31,137,31,131,31,74,31,61,31,61,30,37,31,37,30,37,29,34,31,34,30,200,31,240,31,151,31,23,31,108,31,229,31,68,31,173,31,53,31,3,31,65,31,65,30,65,29,65,28,96,31,154,31,243,31,138,31,29,31,36,31,157,31,85,31,220,31,85,31,90,31,114,31,111,31,245,31,151,31,151,30,247,31,9,31,90,31,78,31,84,31,71,31,73,31,7,31,7,30,165,31,33,31,72,31,72,30,166,31,25,31,239,31,83,31,83,30,174,31,174,30,90,31,216,31,75,31,75,30,75,29,75,28,148,31,72,31,240,31,15,31,15,30,156,31,130,31,16,31,14,31,198,31,137,31,137,30,212,31,122,31,60,31,198,31,176,31,127,31,127,30,127,29,233,31,190,31,81,31,181,31,131,31,244,31,58,31,167,31,167,30,167,29,216,31,25,31,220,31,220,30,220,29,23,31,169,31,202,31,164,31,83,31,83,30,125,31,125,30,116,31,229,31,229,30,155,31,189,31,8,31,8,30,103,31,172,31,211,31,186,31,13,31,62,31,234,31,114,31,193,31,178,31,132,31,132,30,97,31,201,31,180,31,121,31,194,31,219,31,20,31,141,31,141,30,56,31,221,31,38,31,38,31,38,30,196,31,196,30,181,31,181,30,181,29,49,31,2,31,120,31,120,30,225,31,106,31,217,31,45,31,210,31,156,31,162,31,176,31,213,31,35,31,96,31,155,31,172,31,172,30,172,29,156,31,193,31,43,31,102,31,102,30,102,29,64,31,64,30,118,31,118,30,237,31,126,31,195,31,57,31,98,31,98,30,122,31,122,30,222,31,179,31,148,31,94,31,94,30,113,31,148,31,148,30,151,31,232,31,239,31,212,31,102,31,207,31,116,31,221,31,67,31,147,31,176,31,248,31,248,30,207,31,224,31,24,31,105,31,105,30,8,31,174,31,67,31,249,31,249,30,217,31,251,31,251,30,115,31,51,31,140,31,161,31,136,31,105,31,125,31,155,31,174,31,18,31,114,31,114,30,246,31,246,30,18,31,206,31,251,31,237,31,237,30,165,31,95,31,86,31,86,30,103,31,176,31,176,30,1,31,207,31,122,31,112,31,102,31,102,30,242,31,199,31,91,31,91,30,146,31,67,31,252,31,222,31,144,31,144,30,100,31,176,31,224,31,212,31,50,31,240,31,216,31,216,30,214,31,103,31,166,31,246,31,246,30,67,31,62,31,17,31,17,30,121,31,172,31,141,31,141,30,201,31,117,31,254,31,13,31,213,31,152,31,124,31,147,31,73,31,189,31,50,31,167,31,193,31,13,31,211,31,211,30,211,29,85,31,85,30,113,31,27,31,120,31,120,30,36,31,36,30,166,31,251,31,217,31,241,31,111,31,125,31,125,30,125,29,47,31,114,31,49,31,126,31,188,31,100,31,115,31,242,31,15,31,15,30,15,29,144,31,144,30,23,31,23,30,23,29,169,31,33,31,143,31,138,31,138,30,237,31,237,30,237,29,217,31,20,31,44,31,225,31,65,31,47,31,124,31,181,31,181,30,181,29,55,31,55,30,1,31,35,31,161,31,46,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
