-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 189;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (84,0,98,0,245,0,148,0,189,0,21,0,121,0,108,0,132,0,112,0,23,0,34,0,0,0,248,0,0,0,0,0,234,0,160,0,225,0,120,0,93,0,8,0,126,0,0,0,203,0,230,0,161,0,71,0,52,0,0,0,0,0,0,0,0,0,63,0,228,0,224,0,211,0,35,0,200,0,10,0,86,0,0,0,26,0,0,0,247,0,235,0,0,0,0,0,195,0,235,0,50,0,41,0,181,0,189,0,70,0,134,0,70,0,0,0,155,0,115,0,38,0,0,0,222,0,205,0,36,0,0,0,51,0,0,0,0,0,56,0,247,0,157,0,192,0,192,0,209,0,212,0,90,0,27,0,0,0,183,0,0,0,173,0,210,0,0,0,135,0,229,0,131,0,218,0,138,0,43,0,26,0,231,0,222,0,75,0,0,0,248,0,66,0,0,0,72,0,244,0,0,0,30,0,77,0,0,0,235,0,238,0,84,0,104,0,139,0,0,0,55,0,125,0,5,0,104,0,40,0,183,0,228,0,177,0,94,0,141,0,76,0,227,0,0,0,64,0,169,0,231,0,231,0,39,0,0,0,36,0,0,0,7,0,199,0,0,0,49,0,4,0,0,0,35,0,223,0,243,0,81,0,0,0,88,0,147,0,180,0,150,0,233,0,142,0,111,0,171,0,53,0,239,0,130,0,16,0,103,0,210,0,141,0,172,0,193,0,1,0,122,0,116,0,47,0,0,0,0,0,115,0,91,0,108,0,79,0,103,0,19,0,22,0,0,0,110,0,15,0,54,0,44,0,0,0,245,0,129,0,210,0,123,0,110,0,0,0,9,0,0,0,0,0,103,0,0,0);
signal scenario_full  : scenario_type := (84,31,98,31,245,31,148,31,189,31,21,31,121,31,108,31,132,31,112,31,23,31,34,31,34,30,248,31,248,30,248,29,234,31,160,31,225,31,120,31,93,31,8,31,126,31,126,30,203,31,230,31,161,31,71,31,52,31,52,30,52,29,52,28,52,27,63,31,228,31,224,31,211,31,35,31,200,31,10,31,86,31,86,30,26,31,26,30,247,31,235,31,235,30,235,29,195,31,235,31,50,31,41,31,181,31,189,31,70,31,134,31,70,31,70,30,155,31,115,31,38,31,38,30,222,31,205,31,36,31,36,30,51,31,51,30,51,29,56,31,247,31,157,31,192,31,192,31,209,31,212,31,90,31,27,31,27,30,183,31,183,30,173,31,210,31,210,30,135,31,229,31,131,31,218,31,138,31,43,31,26,31,231,31,222,31,75,31,75,30,248,31,66,31,66,30,72,31,244,31,244,30,30,31,77,31,77,30,235,31,238,31,84,31,104,31,139,31,139,30,55,31,125,31,5,31,104,31,40,31,183,31,228,31,177,31,94,31,141,31,76,31,227,31,227,30,64,31,169,31,231,31,231,31,39,31,39,30,36,31,36,30,7,31,199,31,199,30,49,31,4,31,4,30,35,31,223,31,243,31,81,31,81,30,88,31,147,31,180,31,150,31,233,31,142,31,111,31,171,31,53,31,239,31,130,31,16,31,103,31,210,31,141,31,172,31,193,31,1,31,122,31,116,31,47,31,47,30,47,29,115,31,91,31,108,31,79,31,103,31,19,31,22,31,22,30,110,31,15,31,54,31,44,31,44,30,245,31,129,31,210,31,123,31,110,31,110,30,9,31,9,30,9,29,103,31,103,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
