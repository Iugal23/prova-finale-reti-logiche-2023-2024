-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_832 is
end project_tb_832;

architecture project_tb_arch_832 of project_tb_832 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 876;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (10,0,192,0,254,0,0,0,157,0,208,0,107,0,188,0,242,0,42,0,0,0,50,0,20,0,18,0,109,0,223,0,0,0,99,0,75,0,71,0,249,0,131,0,127,0,0,0,127,0,195,0,32,0,35,0,32,0,215,0,178,0,144,0,250,0,187,0,232,0,178,0,30,0,96,0,182,0,0,0,0,0,0,0,218,0,62,0,174,0,249,0,88,0,73,0,204,0,40,0,28,0,149,0,0,0,12,0,131,0,243,0,0,0,217,0,14,0,240,0,249,0,156,0,81,0,0,0,170,0,14,0,0,0,75,0,0,0,20,0,237,0,115,0,6,0,46,0,22,0,3,0,65,0,0,0,230,0,0,0,0,0,64,0,131,0,0,0,0,0,77,0,0,0,46,0,250,0,38,0,251,0,25,0,243,0,0,0,32,0,190,0,86,0,97,0,128,0,0,0,144,0,230,0,169,0,231,0,0,0,229,0,33,0,238,0,164,0,140,0,117,0,175,0,50,0,129,0,170,0,63,0,192,0,207,0,14,0,136,0,137,0,51,0,81,0,171,0,68,0,43,0,0,0,35,0,145,0,89,0,130,0,215,0,204,0,0,0,48,0,0,0,116,0,72,0,82,0,110,0,107,0,0,0,146,0,75,0,126,0,236,0,8,0,129,0,253,0,133,0,0,0,200,0,0,0,29,0,191,0,0,0,0,0,110,0,247,0,0,0,235,0,74,0,183,0,143,0,0,0,0,0,59,0,48,0,50,0,0,0,250,0,80,0,72,0,90,0,0,0,128,0,84,0,214,0,215,0,189,0,211,0,2,0,63,0,220,0,98,0,89,0,182,0,83,0,133,0,156,0,166,0,201,0,70,0,0,0,0,0,45,0,184,0,146,0,17,0,189,0,154,0,175,0,137,0,25,0,29,0,94,0,85,0,103,0,189,0,139,0,0,0,85,0,172,0,195,0,57,0,11,0,209,0,0,0,100,0,52,0,25,0,5,0,219,0,163,0,0,0,60,0,0,0,193,0,93,0,129,0,10,0,5,0,0,0,88,0,46,0,0,0,0,0,106,0,0,0,113,0,0,0,97,0,0,0,85,0,16,0,51,0,107,0,6,0,230,0,159,0,245,0,97,0,120,0,208,0,209,0,204,0,0,0,0,0,89,0,72,0,173,0,11,0,47,0,62,0,20,0,254,0,22,0,70,0,0,0,0,0,102,0,248,0,0,0,51,0,14,0,79,0,8,0,162,0,188,0,38,0,228,0,194,0,0,0,216,0,122,0,204,0,232,0,0,0,228,0,0,0,226,0,231,0,0,0,134,0,127,0,0,0,226,0,0,0,95,0,107,0,0,0,137,0,86,0,201,0,200,0,180,0,168,0,90,0,0,0,81,0,0,0,83,0,137,0,72,0,163,0,0,0,0,0,0,0,0,0,22,0,74,0,101,0,62,0,39,0,0,0,0,0,211,0,0,0,0,0,0,0,105,0,91,0,36,0,0,0,252,0,0,0,0,0,100,0,233,0,211,0,4,0,0,0,0,0,131,0,136,0,151,0,184,0,214,0,82,0,134,0,64,0,61,0,24,0,201,0,150,0,160,0,215,0,184,0,80,0,157,0,98,0,0,0,206,0,177,0,166,0,146,0,80,0,5,0,67,0,25,0,246,0,0,0,129,0,162,0,43,0,247,0,170,0,194,0,56,0,90,0,117,0,109,0,201,0,0,0,127,0,191,0,201,0,32,0,156,0,209,0,246,0,170,0,0,0,52,0,37,0,42,0,20,0,82,0,62,0,22,0,25,0,243,0,145,0,57,0,11,0,0,0,77,0,226,0,0,0,24,0,229,0,202,0,108,0,124,0,0,0,157,0,218,0,254,0,53,0,106,0,161,0,186,0,0,0,163,0,136,0,0,0,105,0,122,0,124,0,12,0,70,0,212,0,152,0,0,0,117,0,250,0,109,0,66,0,63,0,109,0,0,0,212,0,216,0,113,0,151,0,146,0,16,0,255,0,69,0,0,0,15,0,58,0,169,0,13,0,160,0,245,0,167,0,209,0,0,0,98,0,21,0,155,0,48,0,244,0,8,0,142,0,18,0,230,0,0,0,97,0,0,0,133,0,0,0,71,0,29,0,29,0,92,0,0,0,0,0,0,0,45,0,32,0,42,0,241,0,192,0,59,0,67,0,46,0,24,0,135,0,210,0,122,0,140,0,0,0,195,0,245,0,0,0,0,0,166,0,248,0,0,0,0,0,166,0,143,0,11,0,228,0,220,0,249,0,0,0,0,0,28,0,0,0,212,0,30,0,137,0,36,0,0,0,56,0,138,0,50,0,40,0,28,0,0,0,238,0,66,0,88,0,235,0,200,0,0,0,170,0,98,0,81,0,191,0,61,0,218,0,10,0,148,0,0,0,112,0,0,0,0,0,176,0,126,0,0,0,45,0,234,0,0,0,0,0,193,0,6,0,192,0,19,0,105,0,200,0,12,0,57,0,31,0,135,0,29,0,22,0,0,0,0,0,0,0,0,0,148,0,97,0,192,0,10,0,218,0,0,0,43,0,61,0,207,0,165,0,75,0,188,0,162,0,2,0,0,0,50,0,58,0,39,0,237,0,251,0,112,0,150,0,34,0,0,0,0,0,241,0,210,0,184,0,0,0,188,0,151,0,229,0,133,0,0,0,94,0,0,0,56,0,115,0,0,0,0,0,0,0,149,0,213,0,71,0,216,0,105,0,0,0,0,0,106,0,69,0,135,0,6,0,227,0,211,0,0,0,231,0,213,0,218,0,125,0,253,0,103,0,25,0,158,0,216,0,0,0,39,0,117,0,0,0,64,0,22,0,0,0,64,0,167,0,134,0,230,0,4,0,210,0,171,0,68,0,0,0,179,0,209,0,208,0,231,0,125,0,46,0,255,0,0,0,122,0,160,0,31,0,173,0,44,0,69,0,130,0,201,0,67,0,134,0,247,0,0,0,180,0,6,0,7,0,0,0,145,0,6,0,32,0,0,0,95,0,149,0,109,0,77,0,0,0,58,0,208,0,50,0,0,0,0,0,197,0,214,0,0,0,0,0,0,0,92,0,176,0,0,0,113,0,0,0,0,0,242,0,173,0,0,0,240,0,126,0,85,0,0,0,172,0,0,0,170,0,239,0,55,0,225,0,0,0,200,0,249,0,0,0,231,0,168,0,213,0,189,0,245,0,0,0,86,0,226,0,161,0,165,0,219,0,0,0,38,0,0,0,41,0,147,0,172,0,0,0,182,0,175,0,152,0,126,0,120,0,0,0,100,0,143,0,77,0,56,0,74,0,234,0,0,0,69,0,0,0,119,0,132,0,133,0,0,0,160,0,234,0,138,0,151,0,236,0,0,0,219,0,219,0,83,0,60,0,0,0,27,0,184,0,201,0,87,0,27,0,220,0,173,0,230,0,155,0,13,0,64,0,79,0,210,0,100,0,0,0,25,0,0,0,253,0,152,0,0,0,214,0,97,0,123,0,0,0,120,0,0,0,12,0,0,0,0,0,227,0,218,0,79,0,0,0,83,0,78,0,104,0,0,0,104,0,137,0,222,0,95,0,0,0,0,0,118,0,98,0,110,0,150,0,147,0,71,0,0,0,75,0,115,0,190,0,122,0,212,0,198,0,46,0,199,0,112,0,182,0,227,0,131,0,99,0,234,0,0,0,24,0,0,0,192,0,93,0,241,0,93,0,122,0,0,0,89,0,188,0,61,0,20,0,32,0,162,0,120,0,142,0,229,0,86,0,0,0,237,0,231,0,0,0,199,0,185,0,0,0,10,0,210,0,242,0,231,0,0,0,142,0,141,0,79,0,200,0,0,0,236,0,249,0,0,0,0,0,166,0,0,0,44,0,208,0,95,0,18,0,0,0,65,0,58,0,65,0,54,0,220,0,149,0,27,0);
signal scenario_full  : scenario_type := (10,31,192,31,254,31,254,30,157,31,208,31,107,31,188,31,242,31,42,31,42,30,50,31,20,31,18,31,109,31,223,31,223,30,99,31,75,31,71,31,249,31,131,31,127,31,127,30,127,31,195,31,32,31,35,31,32,31,215,31,178,31,144,31,250,31,187,31,232,31,178,31,30,31,96,31,182,31,182,30,182,29,182,28,218,31,62,31,174,31,249,31,88,31,73,31,204,31,40,31,28,31,149,31,149,30,12,31,131,31,243,31,243,30,217,31,14,31,240,31,249,31,156,31,81,31,81,30,170,31,14,31,14,30,75,31,75,30,20,31,237,31,115,31,6,31,46,31,22,31,3,31,65,31,65,30,230,31,230,30,230,29,64,31,131,31,131,30,131,29,77,31,77,30,46,31,250,31,38,31,251,31,25,31,243,31,243,30,32,31,190,31,86,31,97,31,128,31,128,30,144,31,230,31,169,31,231,31,231,30,229,31,33,31,238,31,164,31,140,31,117,31,175,31,50,31,129,31,170,31,63,31,192,31,207,31,14,31,136,31,137,31,51,31,81,31,171,31,68,31,43,31,43,30,35,31,145,31,89,31,130,31,215,31,204,31,204,30,48,31,48,30,116,31,72,31,82,31,110,31,107,31,107,30,146,31,75,31,126,31,236,31,8,31,129,31,253,31,133,31,133,30,200,31,200,30,29,31,191,31,191,30,191,29,110,31,247,31,247,30,235,31,74,31,183,31,143,31,143,30,143,29,59,31,48,31,50,31,50,30,250,31,80,31,72,31,90,31,90,30,128,31,84,31,214,31,215,31,189,31,211,31,2,31,63,31,220,31,98,31,89,31,182,31,83,31,133,31,156,31,166,31,201,31,70,31,70,30,70,29,45,31,184,31,146,31,17,31,189,31,154,31,175,31,137,31,25,31,29,31,94,31,85,31,103,31,189,31,139,31,139,30,85,31,172,31,195,31,57,31,11,31,209,31,209,30,100,31,52,31,25,31,5,31,219,31,163,31,163,30,60,31,60,30,193,31,93,31,129,31,10,31,5,31,5,30,88,31,46,31,46,30,46,29,106,31,106,30,113,31,113,30,97,31,97,30,85,31,16,31,51,31,107,31,6,31,230,31,159,31,245,31,97,31,120,31,208,31,209,31,204,31,204,30,204,29,89,31,72,31,173,31,11,31,47,31,62,31,20,31,254,31,22,31,70,31,70,30,70,29,102,31,248,31,248,30,51,31,14,31,79,31,8,31,162,31,188,31,38,31,228,31,194,31,194,30,216,31,122,31,204,31,232,31,232,30,228,31,228,30,226,31,231,31,231,30,134,31,127,31,127,30,226,31,226,30,95,31,107,31,107,30,137,31,86,31,201,31,200,31,180,31,168,31,90,31,90,30,81,31,81,30,83,31,137,31,72,31,163,31,163,30,163,29,163,28,163,27,22,31,74,31,101,31,62,31,39,31,39,30,39,29,211,31,211,30,211,29,211,28,105,31,91,31,36,31,36,30,252,31,252,30,252,29,100,31,233,31,211,31,4,31,4,30,4,29,131,31,136,31,151,31,184,31,214,31,82,31,134,31,64,31,61,31,24,31,201,31,150,31,160,31,215,31,184,31,80,31,157,31,98,31,98,30,206,31,177,31,166,31,146,31,80,31,5,31,67,31,25,31,246,31,246,30,129,31,162,31,43,31,247,31,170,31,194,31,56,31,90,31,117,31,109,31,201,31,201,30,127,31,191,31,201,31,32,31,156,31,209,31,246,31,170,31,170,30,52,31,37,31,42,31,20,31,82,31,62,31,22,31,25,31,243,31,145,31,57,31,11,31,11,30,77,31,226,31,226,30,24,31,229,31,202,31,108,31,124,31,124,30,157,31,218,31,254,31,53,31,106,31,161,31,186,31,186,30,163,31,136,31,136,30,105,31,122,31,124,31,12,31,70,31,212,31,152,31,152,30,117,31,250,31,109,31,66,31,63,31,109,31,109,30,212,31,216,31,113,31,151,31,146,31,16,31,255,31,69,31,69,30,15,31,58,31,169,31,13,31,160,31,245,31,167,31,209,31,209,30,98,31,21,31,155,31,48,31,244,31,8,31,142,31,18,31,230,31,230,30,97,31,97,30,133,31,133,30,71,31,29,31,29,31,92,31,92,30,92,29,92,28,45,31,32,31,42,31,241,31,192,31,59,31,67,31,46,31,24,31,135,31,210,31,122,31,140,31,140,30,195,31,245,31,245,30,245,29,166,31,248,31,248,30,248,29,166,31,143,31,11,31,228,31,220,31,249,31,249,30,249,29,28,31,28,30,212,31,30,31,137,31,36,31,36,30,56,31,138,31,50,31,40,31,28,31,28,30,238,31,66,31,88,31,235,31,200,31,200,30,170,31,98,31,81,31,191,31,61,31,218,31,10,31,148,31,148,30,112,31,112,30,112,29,176,31,126,31,126,30,45,31,234,31,234,30,234,29,193,31,6,31,192,31,19,31,105,31,200,31,12,31,57,31,31,31,135,31,29,31,22,31,22,30,22,29,22,28,22,27,148,31,97,31,192,31,10,31,218,31,218,30,43,31,61,31,207,31,165,31,75,31,188,31,162,31,2,31,2,30,50,31,58,31,39,31,237,31,251,31,112,31,150,31,34,31,34,30,34,29,241,31,210,31,184,31,184,30,188,31,151,31,229,31,133,31,133,30,94,31,94,30,56,31,115,31,115,30,115,29,115,28,149,31,213,31,71,31,216,31,105,31,105,30,105,29,106,31,69,31,135,31,6,31,227,31,211,31,211,30,231,31,213,31,218,31,125,31,253,31,103,31,25,31,158,31,216,31,216,30,39,31,117,31,117,30,64,31,22,31,22,30,64,31,167,31,134,31,230,31,4,31,210,31,171,31,68,31,68,30,179,31,209,31,208,31,231,31,125,31,46,31,255,31,255,30,122,31,160,31,31,31,173,31,44,31,69,31,130,31,201,31,67,31,134,31,247,31,247,30,180,31,6,31,7,31,7,30,145,31,6,31,32,31,32,30,95,31,149,31,109,31,77,31,77,30,58,31,208,31,50,31,50,30,50,29,197,31,214,31,214,30,214,29,214,28,92,31,176,31,176,30,113,31,113,30,113,29,242,31,173,31,173,30,240,31,126,31,85,31,85,30,172,31,172,30,170,31,239,31,55,31,225,31,225,30,200,31,249,31,249,30,231,31,168,31,213,31,189,31,245,31,245,30,86,31,226,31,161,31,165,31,219,31,219,30,38,31,38,30,41,31,147,31,172,31,172,30,182,31,175,31,152,31,126,31,120,31,120,30,100,31,143,31,77,31,56,31,74,31,234,31,234,30,69,31,69,30,119,31,132,31,133,31,133,30,160,31,234,31,138,31,151,31,236,31,236,30,219,31,219,31,83,31,60,31,60,30,27,31,184,31,201,31,87,31,27,31,220,31,173,31,230,31,155,31,13,31,64,31,79,31,210,31,100,31,100,30,25,31,25,30,253,31,152,31,152,30,214,31,97,31,123,31,123,30,120,31,120,30,12,31,12,30,12,29,227,31,218,31,79,31,79,30,83,31,78,31,104,31,104,30,104,31,137,31,222,31,95,31,95,30,95,29,118,31,98,31,110,31,150,31,147,31,71,31,71,30,75,31,115,31,190,31,122,31,212,31,198,31,46,31,199,31,112,31,182,31,227,31,131,31,99,31,234,31,234,30,24,31,24,30,192,31,93,31,241,31,93,31,122,31,122,30,89,31,188,31,61,31,20,31,32,31,162,31,120,31,142,31,229,31,86,31,86,30,237,31,231,31,231,30,199,31,185,31,185,30,10,31,210,31,242,31,231,31,231,30,142,31,141,31,79,31,200,31,200,30,236,31,249,31,249,30,249,29,166,31,166,30,44,31,208,31,95,31,18,31,18,30,65,31,58,31,65,31,54,31,220,31,149,31,27,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
