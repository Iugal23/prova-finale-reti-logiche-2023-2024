-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 967;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (146,0,230,0,0,0,224,0,0,0,195,0,0,0,38,0,0,0,0,0,103,0,99,0,178,0,164,0,10,0,234,0,137,0,115,0,74,0,153,0,87,0,69,0,25,0,160,0,144,0,214,0,171,0,60,0,63,0,237,0,252,0,51,0,0,0,142,0,43,0,68,0,232,0,197,0,193,0,33,0,95,0,0,0,0,0,242,0,0,0,189,0,111,0,81,0,223,0,174,0,2,0,104,0,247,0,103,0,46,0,248,0,20,0,204,0,0,0,215,0,141,0,26,0,42,0,118,0,98,0,74,0,0,0,227,0,95,0,185,0,137,0,74,0,43,0,0,0,0,0,154,0,0,0,229,0,10,0,71,0,226,0,165,0,41,0,0,0,206,0,232,0,229,0,150,0,91,0,0,0,70,0,131,0,164,0,170,0,0,0,169,0,208,0,23,0,117,0,92,0,50,0,0,0,51,0,48,0,38,0,191,0,216,0,100,0,0,0,110,0,37,0,177,0,129,0,162,0,200,0,189,0,240,0,138,0,169,0,83,0,6,0,0,0,99,0,44,0,221,0,247,0,224,0,116,0,0,0,231,0,0,0,0,0,14,0,25,0,63,0,0,0,238,0,129,0,101,0,157,0,0,0,178,0,157,0,174,0,61,0,254,0,96,0,0,0,185,0,121,0,0,0,12,0,145,0,147,0,0,0,244,0,55,0,180,0,159,0,87,0,75,0,43,0,80,0,234,0,0,0,0,0,146,0,179,0,113,0,111,0,58,0,38,0,156,0,0,0,97,0,132,0,23,0,27,0,235,0,229,0,189,0,0,0,0,0,0,0,103,0,8,0,0,0,2,0,192,0,0,0,107,0,0,0,212,0,189,0,248,0,137,0,0,0,66,0,183,0,251,0,133,0,14,0,0,0,55,0,0,0,187,0,93,0,0,0,166,0,161,0,79,0,164,0,195,0,78,0,0,0,220,0,58,0,22,0,73,0,213,0,161,0,0,0,0,0,0,0,79,0,88,0,25,0,0,0,170,0,7,0,166,0,0,0,54,0,128,0,217,0,91,0,155,0,83,0,0,0,169,0,246,0,238,0,71,0,0,0,131,0,55,0,91,0,176,0,232,0,0,0,147,0,228,0,214,0,54,0,90,0,121,0,44,0,166,0,206,0,217,0,216,0,198,0,84,0,0,0,155,0,107,0,20,0,55,0,20,0,115,0,38,0,236,0,112,0,219,0,218,0,168,0,198,0,0,0,73,0,61,0,11,0,64,0,198,0,113,0,59,0,239,0,34,0,183,0,24,0,44,0,184,0,40,0,252,0,137,0,44,0,229,0,92,0,0,0,50,0,119,0,107,0,0,0,146,0,129,0,71,0,83,0,55,0,0,0,88,0,130,0,156,0,101,0,188,0,112,0,116,0,0,0,0,0,148,0,53,0,88,0,172,0,170,0,128,0,188,0,0,0,0,0,0,0,210,0,36,0,134,0,81,0,34,0,146,0,170,0,144,0,143,0,230,0,189,0,135,0,0,0,127,0,129,0,130,0,101,0,43,0,128,0,218,0,168,0,142,0,166,0,244,0,185,0,209,0,176,0,219,0,206,0,0,0,137,0,207,0,134,0,76,0,47,0,107,0,182,0,215,0,151,0,23,0,68,0,208,0,160,0,224,0,212,0,186,0,0,0,95,0,0,0,254,0,74,0,180,0,0,0,3,0,192,0,115,0,0,0,243,0,64,0,134,0,0,0,102,0,164,0,118,0,0,0,129,0,39,0,43,0,0,0,118,0,0,0,9,0,192,0,0,0,0,0,130,0,16,0,46,0,187,0,4,0,151,0,233,0,237,0,74,0,208,0,219,0,26,0,149,0,5,0,111,0,30,0,0,0,131,0,248,0,0,0,219,0,3,0,25,0,0,0,56,0,249,0,145,0,120,0,149,0,156,0,0,0,0,0,104,0,0,0,41,0,13,0,248,0,133,0,211,0,7,0,119,0,13,0,89,0,0,0,89,0,0,0,75,0,250,0,172,0,114,0,104,0,84,0,251,0,194,0,0,0,191,0,88,0,8,0,0,0,18,0,82,0,34,0,221,0,199,0,235,0,183,0,0,0,209,0,0,0,0,0,163,0,203,0,0,0,164,0,0,0,32,0,174,0,204,0,63,0,0,0,113,0,158,0,214,0,16,0,35,0,159,0,219,0,152,0,1,0,223,0,0,0,91,0,0,0,0,0,66,0,0,0,31,0,28,0,91,0,220,0,56,0,21,0,189,0,160,0,127,0,160,0,235,0,134,0,227,0,226,0,0,0,198,0,9,0,84,0,95,0,155,0,49,0,59,0,0,0,154,0,165,0,187,0,173,0,216,0,100,0,97,0,252,0,68,0,0,0,189,0,201,0,240,0,163,0,249,0,0,0,104,0,5,0,0,0,4,0,61,0,119,0,24,0,43,0,24,0,250,0,0,0,160,0,185,0,244,0,0,0,37,0,121,0,44,0,0,0,179,0,85,0,82,0,0,0,0,0,224,0,82,0,0,0,105,0,168,0,8,0,151,0,0,0,161,0,0,0,201,0,95,0,85,0,156,0,0,0,141,0,14,0,155,0,207,0,0,0,159,0,4,0,0,0,184,0,0,0,0,0,0,0,0,0,121,0,213,0,123,0,0,0,0,0,64,0,0,0,92,0,106,0,81,0,12,0,64,0,185,0,125,0,140,0,0,0,82,0,154,0,81,0,230,0,107,0,146,0,77,0,222,0,52,0,80,0,106,0,76,0,162,0,39,0,0,0,0,0,130,0,104,0,119,0,209,0,0,0,38,0,150,0,48,0,54,0,122,0,0,0,253,0,224,0,91,0,109,0,183,0,160,0,196,0,0,0,39,0,222,0,99,0,149,0,127,0,0,0,191,0,86,0,246,0,0,0,75,0,145,0,4,0,68,0,205,0,223,0,24,0,0,0,204,0,24,0,65,0,248,0,17,0,0,0,72,0,24,0,51,0,99,0,68,0,51,0,225,0,134,0,153,0,46,0,214,0,148,0,115,0,0,0,132,0,0,0,88,0,0,0,96,0,57,0,126,0,12,0,214,0,208,0,110,0,83,0,29,0,224,0,155,0,58,0,147,0,0,0,160,0,61,0,145,0,31,0,140,0,7,0,107,0,1,0,11,0,0,0,236,0,17,0,0,0,164,0,145,0,28,0,77,0,158,0,83,0,36,0,85,0,78,0,0,0,65,0,171,0,168,0,0,0,0,0,134,0,117,0,234,0,0,0,18,0,179,0,197,0,0,0,51,0,246,0,250,0,142,0,43,0,0,0,43,0,124,0,0,0,254,0,6,0,0,0,6,0,0,0,132,0,0,0,9,0,161,0,93,0,188,0,224,0,79,0,121,0,97,0,0,0,61,0,6,0,225,0,0,0,5,0,120,0,12,0,217,0,183,0,31,0,134,0,201,0,213,0,130,0,252,0,138,0,78,0,0,0,37,0,145,0,0,0,196,0,78,0,148,0,37,0,225,0,36,0,200,0,0,0,121,0,28,0,215,0,41,0,0,0,0,0,58,0,57,0,106,0,77,0,4,0,197,0,182,0,222,0,97,0,233,0,6,0,0,0,123,0,24,0,0,0,0,0,136,0,102,0,182,0,116,0,154,0,182,0,0,0,0,0,63,0,175,0,195,0,95,0,136,0,82,0,61,0,178,0,15,0,97,0,189,0,187,0,107,0,0,0,243,0,188,0,0,0,0,0,107,0,211,0,31,0,90,0,161,0,0,0,126,0,54,0,254,0,0,0,0,0,64,0,161,0,134,0,230,0,188,0,173,0,0,0,196,0,57,0,0,0,81,0,67,0,154,0,220,0,16,0,0,0,107,0,147,0,111,0,0,0,129,0,222,0,80,0,141,0,42,0,0,0,0,0,67,0,134,0,107,0,232,0,70,0,0,0,120,0,238,0,236,0,208,0,159,0,0,0,178,0,59,0,20,0,17,0,207,0,56,0,0,0,184,0,0,0,0,0,21,0,26,0,233,0,175,0,26,0,0,0,7,0,92,0,52,0,225,0,0,0,0,0,11,0,163,0,0,0,0,0,2,0,0,0,177,0,175,0,188,0,197,0,0,0,135,0,230,0,176,0,3,0,143,0,48,0,15,0,220,0,253,0,123,0,180,0,249,0,162,0,28,0,254,0,245,0,0,0,227,0,0,0,0,0,16,0,218,0,136,0,107,0,92,0,119,0,99,0,5,0,248,0,105,0,235,0,46,0,82,0,35,0,90,0,209,0,126,0,3,0,192,0,238,0,0,0,22,0,25,0,197,0,221,0,213,0,189,0,221,0,16,0,25,0);
signal scenario_full  : scenario_type := (146,31,230,31,230,30,224,31,224,30,195,31,195,30,38,31,38,30,38,29,103,31,99,31,178,31,164,31,10,31,234,31,137,31,115,31,74,31,153,31,87,31,69,31,25,31,160,31,144,31,214,31,171,31,60,31,63,31,237,31,252,31,51,31,51,30,142,31,43,31,68,31,232,31,197,31,193,31,33,31,95,31,95,30,95,29,242,31,242,30,189,31,111,31,81,31,223,31,174,31,2,31,104,31,247,31,103,31,46,31,248,31,20,31,204,31,204,30,215,31,141,31,26,31,42,31,118,31,98,31,74,31,74,30,227,31,95,31,185,31,137,31,74,31,43,31,43,30,43,29,154,31,154,30,229,31,10,31,71,31,226,31,165,31,41,31,41,30,206,31,232,31,229,31,150,31,91,31,91,30,70,31,131,31,164,31,170,31,170,30,169,31,208,31,23,31,117,31,92,31,50,31,50,30,51,31,48,31,38,31,191,31,216,31,100,31,100,30,110,31,37,31,177,31,129,31,162,31,200,31,189,31,240,31,138,31,169,31,83,31,6,31,6,30,99,31,44,31,221,31,247,31,224,31,116,31,116,30,231,31,231,30,231,29,14,31,25,31,63,31,63,30,238,31,129,31,101,31,157,31,157,30,178,31,157,31,174,31,61,31,254,31,96,31,96,30,185,31,121,31,121,30,12,31,145,31,147,31,147,30,244,31,55,31,180,31,159,31,87,31,75,31,43,31,80,31,234,31,234,30,234,29,146,31,179,31,113,31,111,31,58,31,38,31,156,31,156,30,97,31,132,31,23,31,27,31,235,31,229,31,189,31,189,30,189,29,189,28,103,31,8,31,8,30,2,31,192,31,192,30,107,31,107,30,212,31,189,31,248,31,137,31,137,30,66,31,183,31,251,31,133,31,14,31,14,30,55,31,55,30,187,31,93,31,93,30,166,31,161,31,79,31,164,31,195,31,78,31,78,30,220,31,58,31,22,31,73,31,213,31,161,31,161,30,161,29,161,28,79,31,88,31,25,31,25,30,170,31,7,31,166,31,166,30,54,31,128,31,217,31,91,31,155,31,83,31,83,30,169,31,246,31,238,31,71,31,71,30,131,31,55,31,91,31,176,31,232,31,232,30,147,31,228,31,214,31,54,31,90,31,121,31,44,31,166,31,206,31,217,31,216,31,198,31,84,31,84,30,155,31,107,31,20,31,55,31,20,31,115,31,38,31,236,31,112,31,219,31,218,31,168,31,198,31,198,30,73,31,61,31,11,31,64,31,198,31,113,31,59,31,239,31,34,31,183,31,24,31,44,31,184,31,40,31,252,31,137,31,44,31,229,31,92,31,92,30,50,31,119,31,107,31,107,30,146,31,129,31,71,31,83,31,55,31,55,30,88,31,130,31,156,31,101,31,188,31,112,31,116,31,116,30,116,29,148,31,53,31,88,31,172,31,170,31,128,31,188,31,188,30,188,29,188,28,210,31,36,31,134,31,81,31,34,31,146,31,170,31,144,31,143,31,230,31,189,31,135,31,135,30,127,31,129,31,130,31,101,31,43,31,128,31,218,31,168,31,142,31,166,31,244,31,185,31,209,31,176,31,219,31,206,31,206,30,137,31,207,31,134,31,76,31,47,31,107,31,182,31,215,31,151,31,23,31,68,31,208,31,160,31,224,31,212,31,186,31,186,30,95,31,95,30,254,31,74,31,180,31,180,30,3,31,192,31,115,31,115,30,243,31,64,31,134,31,134,30,102,31,164,31,118,31,118,30,129,31,39,31,43,31,43,30,118,31,118,30,9,31,192,31,192,30,192,29,130,31,16,31,46,31,187,31,4,31,151,31,233,31,237,31,74,31,208,31,219,31,26,31,149,31,5,31,111,31,30,31,30,30,131,31,248,31,248,30,219,31,3,31,25,31,25,30,56,31,249,31,145,31,120,31,149,31,156,31,156,30,156,29,104,31,104,30,41,31,13,31,248,31,133,31,211,31,7,31,119,31,13,31,89,31,89,30,89,31,89,30,75,31,250,31,172,31,114,31,104,31,84,31,251,31,194,31,194,30,191,31,88,31,8,31,8,30,18,31,82,31,34,31,221,31,199,31,235,31,183,31,183,30,209,31,209,30,209,29,163,31,203,31,203,30,164,31,164,30,32,31,174,31,204,31,63,31,63,30,113,31,158,31,214,31,16,31,35,31,159,31,219,31,152,31,1,31,223,31,223,30,91,31,91,30,91,29,66,31,66,30,31,31,28,31,91,31,220,31,56,31,21,31,189,31,160,31,127,31,160,31,235,31,134,31,227,31,226,31,226,30,198,31,9,31,84,31,95,31,155,31,49,31,59,31,59,30,154,31,165,31,187,31,173,31,216,31,100,31,97,31,252,31,68,31,68,30,189,31,201,31,240,31,163,31,249,31,249,30,104,31,5,31,5,30,4,31,61,31,119,31,24,31,43,31,24,31,250,31,250,30,160,31,185,31,244,31,244,30,37,31,121,31,44,31,44,30,179,31,85,31,82,31,82,30,82,29,224,31,82,31,82,30,105,31,168,31,8,31,151,31,151,30,161,31,161,30,201,31,95,31,85,31,156,31,156,30,141,31,14,31,155,31,207,31,207,30,159,31,4,31,4,30,184,31,184,30,184,29,184,28,184,27,121,31,213,31,123,31,123,30,123,29,64,31,64,30,92,31,106,31,81,31,12,31,64,31,185,31,125,31,140,31,140,30,82,31,154,31,81,31,230,31,107,31,146,31,77,31,222,31,52,31,80,31,106,31,76,31,162,31,39,31,39,30,39,29,130,31,104,31,119,31,209,31,209,30,38,31,150,31,48,31,54,31,122,31,122,30,253,31,224,31,91,31,109,31,183,31,160,31,196,31,196,30,39,31,222,31,99,31,149,31,127,31,127,30,191,31,86,31,246,31,246,30,75,31,145,31,4,31,68,31,205,31,223,31,24,31,24,30,204,31,24,31,65,31,248,31,17,31,17,30,72,31,24,31,51,31,99,31,68,31,51,31,225,31,134,31,153,31,46,31,214,31,148,31,115,31,115,30,132,31,132,30,88,31,88,30,96,31,57,31,126,31,12,31,214,31,208,31,110,31,83,31,29,31,224,31,155,31,58,31,147,31,147,30,160,31,61,31,145,31,31,31,140,31,7,31,107,31,1,31,11,31,11,30,236,31,17,31,17,30,164,31,145,31,28,31,77,31,158,31,83,31,36,31,85,31,78,31,78,30,65,31,171,31,168,31,168,30,168,29,134,31,117,31,234,31,234,30,18,31,179,31,197,31,197,30,51,31,246,31,250,31,142,31,43,31,43,30,43,31,124,31,124,30,254,31,6,31,6,30,6,31,6,30,132,31,132,30,9,31,161,31,93,31,188,31,224,31,79,31,121,31,97,31,97,30,61,31,6,31,225,31,225,30,5,31,120,31,12,31,217,31,183,31,31,31,134,31,201,31,213,31,130,31,252,31,138,31,78,31,78,30,37,31,145,31,145,30,196,31,78,31,148,31,37,31,225,31,36,31,200,31,200,30,121,31,28,31,215,31,41,31,41,30,41,29,58,31,57,31,106,31,77,31,4,31,197,31,182,31,222,31,97,31,233,31,6,31,6,30,123,31,24,31,24,30,24,29,136,31,102,31,182,31,116,31,154,31,182,31,182,30,182,29,63,31,175,31,195,31,95,31,136,31,82,31,61,31,178,31,15,31,97,31,189,31,187,31,107,31,107,30,243,31,188,31,188,30,188,29,107,31,211,31,31,31,90,31,161,31,161,30,126,31,54,31,254,31,254,30,254,29,64,31,161,31,134,31,230,31,188,31,173,31,173,30,196,31,57,31,57,30,81,31,67,31,154,31,220,31,16,31,16,30,107,31,147,31,111,31,111,30,129,31,222,31,80,31,141,31,42,31,42,30,42,29,67,31,134,31,107,31,232,31,70,31,70,30,120,31,238,31,236,31,208,31,159,31,159,30,178,31,59,31,20,31,17,31,207,31,56,31,56,30,184,31,184,30,184,29,21,31,26,31,233,31,175,31,26,31,26,30,7,31,92,31,52,31,225,31,225,30,225,29,11,31,163,31,163,30,163,29,2,31,2,30,177,31,175,31,188,31,197,31,197,30,135,31,230,31,176,31,3,31,143,31,48,31,15,31,220,31,253,31,123,31,180,31,249,31,162,31,28,31,254,31,245,31,245,30,227,31,227,30,227,29,16,31,218,31,136,31,107,31,92,31,119,31,99,31,5,31,248,31,105,31,235,31,46,31,82,31,35,31,90,31,209,31,126,31,3,31,192,31,238,31,238,30,22,31,25,31,197,31,221,31,213,31,189,31,221,31,16,31,25,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
