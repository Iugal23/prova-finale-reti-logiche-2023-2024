-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 863;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,118,0,108,0,202,0,151,0,49,0,249,0,118,0,0,0,28,0,92,0,186,0,0,0,156,0,83,0,100,0,224,0,0,0,254,0,223,0,94,0,62,0,111,0,49,0,178,0,180,0,83,0,251,0,225,0,15,0,0,0,0,0,207,0,0,0,0,0,0,0,254,0,111,0,242,0,0,0,145,0,60,0,140,0,32,0,0,0,40,0,248,0,240,0,0,0,71,0,0,0,180,0,18,0,0,0,3,0,198,0,183,0,0,0,209,0,0,0,240,0,128,0,27,0,132,0,250,0,116,0,0,0,70,0,205,0,217,0,35,0,0,0,0,0,229,0,121,0,129,0,197,0,0,0,160,0,105,0,104,0,65,0,97,0,35,0,0,0,0,0,210,0,73,0,0,0,38,0,0,0,235,0,0,0,0,0,0,0,187,0,248,0,41,0,79,0,37,0,156,0,122,0,67,0,181,0,200,0,86,0,55,0,187,0,201,0,104,0,0,0,42,0,1,0,59,0,58,0,47,0,0,0,0,0,65,0,242,0,2,0,185,0,249,0,0,0,49,0,16,0,117,0,0,0,188,0,132,0,239,0,199,0,124,0,248,0,0,0,51,0,54,0,110,0,95,0,121,0,0,0,0,0,75,0,0,0,3,0,161,0,130,0,0,0,213,0,252,0,0,0,247,0,172,0,154,0,71,0,3,0,14,0,171,0,136,0,231,0,188,0,209,0,80,0,131,0,248,0,31,0,20,0,0,0,67,0,31,0,205,0,16,0,74,0,0,0,152,0,161,0,196,0,219,0,57,0,171,0,218,0,88,0,198,0,139,0,123,0,86,0,151,0,119,0,107,0,0,0,106,0,60,0,55,0,231,0,57,0,3,0,119,0,224,0,66,0,0,0,32,0,150,0,36,0,155,0,0,0,195,0,82,0,0,0,7,0,245,0,112,0,145,0,129,0,154,0,33,0,13,0,237,0,0,0,117,0,97,0,7,0,100,0,160,0,95,0,236,0,49,0,225,0,152,0,234,0,27,0,25,0,163,0,206,0,0,0,110,0,120,0,225,0,151,0,0,0,0,0,240,0,203,0,149,0,25,0,173,0,96,0,55,0,254,0,245,0,137,0,2,0,108,0,217,0,33,0,251,0,0,0,191,0,151,0,0,0,77,0,83,0,217,0,208,0,229,0,114,0,142,0,133,0,69,0,160,0,1,0,106,0,132,0,182,0,0,0,0,0,208,0,46,0,55,0,0,0,0,0,218,0,23,0,88,0,87,0,181,0,0,0,162,0,184,0,16,0,88,0,214,0,228,0,153,0,0,0,255,0,52,0,249,0,110,0,198,0,161,0,191,0,154,0,0,0,26,0,196,0,150,0,57,0,19,0,189,0,113,0,0,0,81,0,105,0,57,0,32,0,38,0,191,0,58,0,85,0,234,0,25,0,120,0,0,0,0,0,231,0,37,0,93,0,255,0,126,0,0,0,0,0,69,0,145,0,0,0,6,0,250,0,195,0,57,0,35,0,109,0,14,0,43,0,0,0,0,0,138,0,198,0,18,0,138,0,155,0,0,0,0,0,189,0,183,0,52,0,0,0,58,0,15,0,0,0,0,0,58,0,239,0,0,0,222,0,0,0,25,0,44,0,168,0,14,0,0,0,78,0,248,0,0,0,198,0,172,0,75,0,142,0,99,0,155,0,41,0,0,0,43,0,173,0,141,0,113,0,246,0,0,0,120,0,217,0,223,0,92,0,84,0,241,0,219,0,0,0,209,0,152,0,144,0,0,0,80,0,0,0,248,0,5,0,201,0,0,0,95,0,19,0,249,0,225,0,36,0,106,0,186,0,208,0,179,0,140,0,200,0,45,0,241,0,159,0,190,0,133,0,167,0,59,0,116,0,174,0,0,0,37,0,0,0,215,0,0,0,82,0,63,0,146,0,95,0,207,0,0,0,149,0,97,0,29,0,68,0,77,0,160,0,40,0,230,0,90,0,167,0,88,0,200,0,145,0,245,0,127,0,110,0,78,0,198,0,17,0,0,0,0,0,90,0,57,0,0,0,142,0,130,0,42,0,113,0,28,0,0,0,173,0,142,0,145,0,0,0,148,0,144,0,0,0,0,0,168,0,41,0,0,0,4,0,0,0,247,0,77,0,37,0,213,0,98,0,148,0,68,0,193,0,0,0,244,0,0,0,149,0,0,0,214,0,0,0,144,0,135,0,183,0,0,0,211,0,125,0,135,0,69,0,159,0,49,0,0,0,156,0,96,0,80,0,168,0,64,0,51,0,0,0,199,0,144,0,43,0,212,0,165,0,53,0,230,0,132,0,240,0,138,0,135,0,28,0,67,0,58,0,247,0,93,0,0,0,0,0,54,0,150,0,230,0,149,0,222,0,160,0,8,0,0,0,54,0,0,0,52,0,0,0,70,0,0,0,176,0,197,0,34,0,138,0,58,0,87,0,170,0,195,0,196,0,129,0,236,0,157,0,199,0,128,0,0,0,0,0,63,0,178,0,168,0,233,0,204,0,248,0,29,0,164,0,0,0,237,0,119,0,182,0,212,0,85,0,26,0,65,0,0,0,92,0,254,0,0,0,0,0,48,0,182,0,152,0,27,0,96,0,0,0,7,0,55,0,58,0,243,0,10,0,24,0,0,0,0,0,211,0,0,0,234,0,54,0,175,0,152,0,248,0,147,0,218,0,65,0,81,0,27,0,98,0,0,0,66,0,15,0,83,0,179,0,244,0,0,0,191,0,0,0,25,0,213,0,18,0,128,0,0,0,223,0,184,0,18,0,73,0,132,0,120,0,0,0,0,0,0,0,185,0,8,0,176,0,0,0,0,0,185,0,29,0,130,0,97,0,155,0,111,0,57,0,142,0,124,0,67,0,95,0,108,0,247,0,0,0,89,0,0,0,239,0,0,0,241,0,84,0,233,0,8,0,0,0,40,0,227,0,53,0,171,0,5,0,193,0,119,0,202,0,11,0,30,0,37,0,254,0,16,0,0,0,187,0,14,0,14,0,231,0,88,0,173,0,125,0,190,0,0,0,0,0,0,0,80,0,90,0,239,0,68,0,79,0,42,0,0,0,103,0,135,0,207,0,204,0,242,0,99,0,188,0,33,0,92,0,22,0,160,0,137,0,33,0,0,0,0,0,134,0,231,0,53,0,0,0,105,0,187,0,213,0,0,0,213,0,0,0,128,0,59,0,231,0,199,0,92,0,140,0,0,0,10,0,0,0,56,0,163,0,61,0,203,0,194,0,12,0,0,0,109,0,106,0,39,0,222,0,11,0,55,0,182,0,148,0,78,0,128,0,144,0,0,0,21,0,126,0,179,0,37,0,89,0,194,0,0,0,207,0,157,0,121,0,0,0,121,0,152,0,36,0,158,0,105,0,0,0,128,0,66,0,244,0,55,0,9,0,119,0,166,0,255,0,26,0,119,0,138,0,0,0,95,0,9,0,66,0,244,0,148,0,0,0,191,0,154,0,180,0,6,0,146,0,25,0,36,0,0,0,109,0,56,0,47,0,0,0,11,0,27,0,131,0,164,0,0,0,0,0,0,0,0,0,248,0,49,0,3,0,143,0,216,0,227,0,53,0,37,0,41,0,215,0,124,0,201,0,197,0,0,0,157,0,42,0,62,0,196,0,56,0,55,0,16,0,112,0,88,0,75,0,160,0,118,0,201,0,88,0,147,0,246,0,219,0,0,0,226,0,154,0,0,0,241,0,0,0,141,0,176,0,175,0,0,0,125,0,0,0,130,0,207,0,76,0,235,0,83,0,0,0,5,0,165,0,84,0,210,0,74,0,250,0,46,0,0,0,93,0,137,0,0,0,246,0,9,0,73,0,44,0,164,0);
signal scenario_full  : scenario_type := (0,0,118,31,108,31,202,31,151,31,49,31,249,31,118,31,118,30,28,31,92,31,186,31,186,30,156,31,83,31,100,31,224,31,224,30,254,31,223,31,94,31,62,31,111,31,49,31,178,31,180,31,83,31,251,31,225,31,15,31,15,30,15,29,207,31,207,30,207,29,207,28,254,31,111,31,242,31,242,30,145,31,60,31,140,31,32,31,32,30,40,31,248,31,240,31,240,30,71,31,71,30,180,31,18,31,18,30,3,31,198,31,183,31,183,30,209,31,209,30,240,31,128,31,27,31,132,31,250,31,116,31,116,30,70,31,205,31,217,31,35,31,35,30,35,29,229,31,121,31,129,31,197,31,197,30,160,31,105,31,104,31,65,31,97,31,35,31,35,30,35,29,210,31,73,31,73,30,38,31,38,30,235,31,235,30,235,29,235,28,187,31,248,31,41,31,79,31,37,31,156,31,122,31,67,31,181,31,200,31,86,31,55,31,187,31,201,31,104,31,104,30,42,31,1,31,59,31,58,31,47,31,47,30,47,29,65,31,242,31,2,31,185,31,249,31,249,30,49,31,16,31,117,31,117,30,188,31,132,31,239,31,199,31,124,31,248,31,248,30,51,31,54,31,110,31,95,31,121,31,121,30,121,29,75,31,75,30,3,31,161,31,130,31,130,30,213,31,252,31,252,30,247,31,172,31,154,31,71,31,3,31,14,31,171,31,136,31,231,31,188,31,209,31,80,31,131,31,248,31,31,31,20,31,20,30,67,31,31,31,205,31,16,31,74,31,74,30,152,31,161,31,196,31,219,31,57,31,171,31,218,31,88,31,198,31,139,31,123,31,86,31,151,31,119,31,107,31,107,30,106,31,60,31,55,31,231,31,57,31,3,31,119,31,224,31,66,31,66,30,32,31,150,31,36,31,155,31,155,30,195,31,82,31,82,30,7,31,245,31,112,31,145,31,129,31,154,31,33,31,13,31,237,31,237,30,117,31,97,31,7,31,100,31,160,31,95,31,236,31,49,31,225,31,152,31,234,31,27,31,25,31,163,31,206,31,206,30,110,31,120,31,225,31,151,31,151,30,151,29,240,31,203,31,149,31,25,31,173,31,96,31,55,31,254,31,245,31,137,31,2,31,108,31,217,31,33,31,251,31,251,30,191,31,151,31,151,30,77,31,83,31,217,31,208,31,229,31,114,31,142,31,133,31,69,31,160,31,1,31,106,31,132,31,182,31,182,30,182,29,208,31,46,31,55,31,55,30,55,29,218,31,23,31,88,31,87,31,181,31,181,30,162,31,184,31,16,31,88,31,214,31,228,31,153,31,153,30,255,31,52,31,249,31,110,31,198,31,161,31,191,31,154,31,154,30,26,31,196,31,150,31,57,31,19,31,189,31,113,31,113,30,81,31,105,31,57,31,32,31,38,31,191,31,58,31,85,31,234,31,25,31,120,31,120,30,120,29,231,31,37,31,93,31,255,31,126,31,126,30,126,29,69,31,145,31,145,30,6,31,250,31,195,31,57,31,35,31,109,31,14,31,43,31,43,30,43,29,138,31,198,31,18,31,138,31,155,31,155,30,155,29,189,31,183,31,52,31,52,30,58,31,15,31,15,30,15,29,58,31,239,31,239,30,222,31,222,30,25,31,44,31,168,31,14,31,14,30,78,31,248,31,248,30,198,31,172,31,75,31,142,31,99,31,155,31,41,31,41,30,43,31,173,31,141,31,113,31,246,31,246,30,120,31,217,31,223,31,92,31,84,31,241,31,219,31,219,30,209,31,152,31,144,31,144,30,80,31,80,30,248,31,5,31,201,31,201,30,95,31,19,31,249,31,225,31,36,31,106,31,186,31,208,31,179,31,140,31,200,31,45,31,241,31,159,31,190,31,133,31,167,31,59,31,116,31,174,31,174,30,37,31,37,30,215,31,215,30,82,31,63,31,146,31,95,31,207,31,207,30,149,31,97,31,29,31,68,31,77,31,160,31,40,31,230,31,90,31,167,31,88,31,200,31,145,31,245,31,127,31,110,31,78,31,198,31,17,31,17,30,17,29,90,31,57,31,57,30,142,31,130,31,42,31,113,31,28,31,28,30,173,31,142,31,145,31,145,30,148,31,144,31,144,30,144,29,168,31,41,31,41,30,4,31,4,30,247,31,77,31,37,31,213,31,98,31,148,31,68,31,193,31,193,30,244,31,244,30,149,31,149,30,214,31,214,30,144,31,135,31,183,31,183,30,211,31,125,31,135,31,69,31,159,31,49,31,49,30,156,31,96,31,80,31,168,31,64,31,51,31,51,30,199,31,144,31,43,31,212,31,165,31,53,31,230,31,132,31,240,31,138,31,135,31,28,31,67,31,58,31,247,31,93,31,93,30,93,29,54,31,150,31,230,31,149,31,222,31,160,31,8,31,8,30,54,31,54,30,52,31,52,30,70,31,70,30,176,31,197,31,34,31,138,31,58,31,87,31,170,31,195,31,196,31,129,31,236,31,157,31,199,31,128,31,128,30,128,29,63,31,178,31,168,31,233,31,204,31,248,31,29,31,164,31,164,30,237,31,119,31,182,31,212,31,85,31,26,31,65,31,65,30,92,31,254,31,254,30,254,29,48,31,182,31,152,31,27,31,96,31,96,30,7,31,55,31,58,31,243,31,10,31,24,31,24,30,24,29,211,31,211,30,234,31,54,31,175,31,152,31,248,31,147,31,218,31,65,31,81,31,27,31,98,31,98,30,66,31,15,31,83,31,179,31,244,31,244,30,191,31,191,30,25,31,213,31,18,31,128,31,128,30,223,31,184,31,18,31,73,31,132,31,120,31,120,30,120,29,120,28,185,31,8,31,176,31,176,30,176,29,185,31,29,31,130,31,97,31,155,31,111,31,57,31,142,31,124,31,67,31,95,31,108,31,247,31,247,30,89,31,89,30,239,31,239,30,241,31,84,31,233,31,8,31,8,30,40,31,227,31,53,31,171,31,5,31,193,31,119,31,202,31,11,31,30,31,37,31,254,31,16,31,16,30,187,31,14,31,14,31,231,31,88,31,173,31,125,31,190,31,190,30,190,29,190,28,80,31,90,31,239,31,68,31,79,31,42,31,42,30,103,31,135,31,207,31,204,31,242,31,99,31,188,31,33,31,92,31,22,31,160,31,137,31,33,31,33,30,33,29,134,31,231,31,53,31,53,30,105,31,187,31,213,31,213,30,213,31,213,30,128,31,59,31,231,31,199,31,92,31,140,31,140,30,10,31,10,30,56,31,163,31,61,31,203,31,194,31,12,31,12,30,109,31,106,31,39,31,222,31,11,31,55,31,182,31,148,31,78,31,128,31,144,31,144,30,21,31,126,31,179,31,37,31,89,31,194,31,194,30,207,31,157,31,121,31,121,30,121,31,152,31,36,31,158,31,105,31,105,30,128,31,66,31,244,31,55,31,9,31,119,31,166,31,255,31,26,31,119,31,138,31,138,30,95,31,9,31,66,31,244,31,148,31,148,30,191,31,154,31,180,31,6,31,146,31,25,31,36,31,36,30,109,31,56,31,47,31,47,30,11,31,27,31,131,31,164,31,164,30,164,29,164,28,164,27,248,31,49,31,3,31,143,31,216,31,227,31,53,31,37,31,41,31,215,31,124,31,201,31,197,31,197,30,157,31,42,31,62,31,196,31,56,31,55,31,16,31,112,31,88,31,75,31,160,31,118,31,201,31,88,31,147,31,246,31,219,31,219,30,226,31,154,31,154,30,241,31,241,30,141,31,176,31,175,31,175,30,125,31,125,30,130,31,207,31,76,31,235,31,83,31,83,30,5,31,165,31,84,31,210,31,74,31,250,31,46,31,46,30,93,31,137,31,137,30,246,31,9,31,73,31,44,31,164,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
