-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_446 is
end project_tb_446;

architecture project_tb_arch_446 of project_tb_446 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 859;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (189,0,102,0,133,0,207,0,78,0,56,0,0,0,119,0,235,0,74,0,0,0,0,0,216,0,0,0,99,0,72,0,56,0,143,0,95,0,154,0,173,0,0,0,0,0,176,0,90,0,21,0,0,0,0,0,0,0,207,0,60,0,106,0,234,0,98,0,245,0,0,0,0,0,145,0,131,0,206,0,201,0,247,0,118,0,70,0,246,0,141,0,0,0,0,0,0,0,151,0,94,0,0,0,0,0,92,0,33,0,126,0,9,0,164,0,90,0,56,0,65,0,172,0,75,0,87,0,180,0,40,0,58,0,137,0,119,0,223,0,244,0,72,0,57,0,0,0,134,0,0,0,66,0,195,0,0,0,223,0,123,0,232,0,77,0,140,0,156,0,73,0,0,0,190,0,58,0,0,0,0,0,170,0,141,0,167,0,131,0,222,0,18,0,46,0,80,0,166,0,176,0,35,0,105,0,96,0,132,0,109,0,0,0,30,0,60,0,47,0,69,0,0,0,11,0,177,0,214,0,161,0,0,0,181,0,193,0,227,0,232,0,98,0,0,0,185,0,103,0,125,0,109,0,0,0,5,0,136,0,29,0,0,0,170,0,27,0,126,0,0,0,189,0,58,0,145,0,55,0,209,0,60,0,15,0,0,0,147,0,0,0,0,0,159,0,127,0,8,0,0,0,132,0,17,0,207,0,0,0,203,0,204,0,228,0,23,0,57,0,253,0,0,0,249,0,254,0,148,0,146,0,0,0,0,0,163,0,181,0,27,0,111,0,9,0,158,0,0,0,91,0,0,0,90,0,83,0,161,0,47,0,209,0,192,0,166,0,247,0,111,0,0,0,0,0,154,0,183,0,55,0,0,0,160,0,163,0,68,0,0,0,0,0,204,0,140,0,2,0,0,0,7,0,99,0,182,0,124,0,0,0,184,0,38,0,181,0,200,0,206,0,22,0,3,0,112,0,150,0,184,0,126,0,63,0,96,0,0,0,75,0,248,0,0,0,0,0,0,0,57,0,87,0,175,0,116,0,0,0,196,0,118,0,220,0,0,0,95,0,144,0,6,0,93,0,95,0,126,0,0,0,2,0,158,0,66,0,214,0,115,0,181,0,44,0,122,0,219,0,103,0,64,0,186,0,0,0,57,0,74,0,71,0,59,0,89,0,0,0,0,0,231,0,65,0,226,0,110,0,0,0,231,0,153,0,166,0,78,0,56,0,19,0,233,0,197,0,130,0,89,0,187,0,220,0,1,0,221,0,160,0,101,0,39,0,38,0,217,0,94,0,202,0,94,0,233,0,97,0,55,0,246,0,133,0,51,0,156,0,255,0,202,0,104,0,91,0,213,0,186,0,111,0,125,0,22,0,0,0,46,0,177,0,0,0,221,0,143,0,250,0,255,0,253,0,235,0,244,0,97,0,133,0,206,0,193,0,229,0,0,0,0,0,179,0,138,0,93,0,127,0,59,0,52,0,21,0,0,0,0,0,0,0,18,0,0,0,144,0,138,0,161,0,113,0,146,0,150,0,247,0,0,0,228,0,0,0,127,0,0,0,0,0,123,0,0,0,188,0,187,0,107,0,231,0,0,0,0,0,122,0,27,0,143,0,211,0,67,0,39,0,197,0,45,0,35,0,103,0,30,0,80,0,86,0,0,0,0,0,12,0,115,0,67,0,246,0,0,0,18,0,51,0,6,0,0,0,113,0,11,0,140,0,14,0,202,0,90,0,0,0,49,0,0,0,194,0,0,0,55,0,107,0,0,0,87,0,129,0,130,0,142,0,0,0,220,0,17,0,0,0,83,0,98,0,249,0,101,0,0,0,187,0,78,0,147,0,82,0,0,0,141,0,145,0,236,0,0,0,101,0,126,0,1,0,0,0,28,0,163,0,0,0,77,0,80,0,58,0,77,0,39,0,12,0,0,0,0,0,236,0,0,0,23,0,11,0,159,0,124,0,105,0,3,0,72,0,170,0,239,0,155,0,156,0,182,0,132,0,0,0,170,0,0,0,110,0,140,0,30,0,252,0,0,0,128,0,210,0,131,0,144,0,156,0,237,0,30,0,41,0,101,0,231,0,21,0,40,0,0,0,162,0,84,0,108,0,12,0,9,0,233,0,140,0,0,0,232,0,0,0,0,0,210,0,26,0,83,0,236,0,246,0,57,0,60,0,0,0,108,0,248,0,107,0,56,0,165,0,0,0,255,0,184,0,17,0,39,0,0,0,0,0,111,0,0,0,209,0,71,0,0,0,47,0,242,0,0,0,127,0,0,0,97,0,254,0,247,0,0,0,0,0,192,0,194,0,101,0,37,0,188,0,254,0,99,0,81,0,0,0,137,0,192,0,0,0,0,0,248,0,71,0,104,0,209,0,153,0,10,0,23,0,52,0,184,0,145,0,255,0,33,0,0,0,17,0,197,0,209,0,242,0,0,0,29,0,6,0,19,0,159,0,169,0,76,0,42,0,0,0,139,0,7,0,37,0,187,0,0,0,171,0,0,0,18,0,58,0,0,0,0,0,0,0,198,0,10,0,30,0,89,0,85,0,128,0,209,0,80,0,245,0,59,0,119,0,112,0,117,0,243,0,250,0,0,0,188,0,181,0,71,0,255,0,213,0,162,0,92,0,106,0,0,0,208,0,35,0,252,0,58,0,108,0,137,0,210,0,15,0,132,0,0,0,34,0,62,0,126,0,23,0,0,0,33,0,209,0,70,0,0,0,0,0,153,0,147,0,191,0,155,0,0,0,67,0,217,0,0,0,49,0,0,0,73,0,0,0,140,0,196,0,248,0,45,0,219,0,222,0,153,0,218,0,227,0,57,0,102,0,30,0,203,0,176,0,196,0,17,0,0,0,29,0,105,0,216,0,4,0,70,0,64,0,64,0,160,0,206,0,33,0,88,0,66,0,0,0,0,0,0,0,0,0,95,0,0,0,0,0,242,0,0,0,149,0,33,0,219,0,36,0,39,0,0,0,116,0,0,0,83,0,111,0,172,0,18,0,0,0,170,0,203,0,0,0,192,0,139,0,0,0,96,0,0,0,15,0,0,0,203,0,182,0,187,0,136,0,0,0,0,0,50,0,186,0,7,0,214,0,25,0,160,0,2,0,0,0,147,0,26,0,0,0,112,0,49,0,150,0,0,0,0,0,187,0,47,0,104,0,10,0,50,0,245,0,215,0,104,0,214,0,222,0,21,0,0,0,251,0,35,0,36,0,43,0,124,0,0,0,129,0,0,0,218,0,81,0,90,0,142,0,0,0,141,0,165,0,198,0,0,0,133,0,103,0,0,0,76,0,18,0,37,0,189,0,0,0,199,0,57,0,116,0,133,0,0,0,216,0,53,0,76,0,35,0,186,0,106,0,82,0,174,0,118,0,42,0,166,0,112,0,212,0,13,0,83,0,164,0,126,0,102,0,37,0,238,0,132,0,176,0,195,0,3,0,116,0,28,0,202,0,151,0,206,0,0,0,121,0,31,0,228,0,140,0,56,0,62,0,244,0,83,0,170,0,0,0,122,0,0,0,28,0,204,0,85,0,0,0,39,0,186,0,197,0,176,0,72,0,169,0,237,0,238,0,255,0,176,0,147,0,0,0,229,0,154,0,252,0,7,0,82,0,21,0,24,0,199,0,59,0,40,0,225,0,181,0,78,0,229,0,0,0,206,0,51,0,0,0,32,0,10,0,8,0,195,0,132,0,0,0,5,0,202,0,220,0,71,0,238,0,27,0,17,0,101,0,151,0,17,0,224,0,57,0,247,0,0,0,0,0,28,0,69,0,132,0,0,0,0,0,230,0,145,0,0,0,167,0,167,0,53,0,0,0,0,0,233,0,55,0,28,0,132,0);
signal scenario_full  : scenario_type := (189,31,102,31,133,31,207,31,78,31,56,31,56,30,119,31,235,31,74,31,74,30,74,29,216,31,216,30,99,31,72,31,56,31,143,31,95,31,154,31,173,31,173,30,173,29,176,31,90,31,21,31,21,30,21,29,21,28,207,31,60,31,106,31,234,31,98,31,245,31,245,30,245,29,145,31,131,31,206,31,201,31,247,31,118,31,70,31,246,31,141,31,141,30,141,29,141,28,151,31,94,31,94,30,94,29,92,31,33,31,126,31,9,31,164,31,90,31,56,31,65,31,172,31,75,31,87,31,180,31,40,31,58,31,137,31,119,31,223,31,244,31,72,31,57,31,57,30,134,31,134,30,66,31,195,31,195,30,223,31,123,31,232,31,77,31,140,31,156,31,73,31,73,30,190,31,58,31,58,30,58,29,170,31,141,31,167,31,131,31,222,31,18,31,46,31,80,31,166,31,176,31,35,31,105,31,96,31,132,31,109,31,109,30,30,31,60,31,47,31,69,31,69,30,11,31,177,31,214,31,161,31,161,30,181,31,193,31,227,31,232,31,98,31,98,30,185,31,103,31,125,31,109,31,109,30,5,31,136,31,29,31,29,30,170,31,27,31,126,31,126,30,189,31,58,31,145,31,55,31,209,31,60,31,15,31,15,30,147,31,147,30,147,29,159,31,127,31,8,31,8,30,132,31,17,31,207,31,207,30,203,31,204,31,228,31,23,31,57,31,253,31,253,30,249,31,254,31,148,31,146,31,146,30,146,29,163,31,181,31,27,31,111,31,9,31,158,31,158,30,91,31,91,30,90,31,83,31,161,31,47,31,209,31,192,31,166,31,247,31,111,31,111,30,111,29,154,31,183,31,55,31,55,30,160,31,163,31,68,31,68,30,68,29,204,31,140,31,2,31,2,30,7,31,99,31,182,31,124,31,124,30,184,31,38,31,181,31,200,31,206,31,22,31,3,31,112,31,150,31,184,31,126,31,63,31,96,31,96,30,75,31,248,31,248,30,248,29,248,28,57,31,87,31,175,31,116,31,116,30,196,31,118,31,220,31,220,30,95,31,144,31,6,31,93,31,95,31,126,31,126,30,2,31,158,31,66,31,214,31,115,31,181,31,44,31,122,31,219,31,103,31,64,31,186,31,186,30,57,31,74,31,71,31,59,31,89,31,89,30,89,29,231,31,65,31,226,31,110,31,110,30,231,31,153,31,166,31,78,31,56,31,19,31,233,31,197,31,130,31,89,31,187,31,220,31,1,31,221,31,160,31,101,31,39,31,38,31,217,31,94,31,202,31,94,31,233,31,97,31,55,31,246,31,133,31,51,31,156,31,255,31,202,31,104,31,91,31,213,31,186,31,111,31,125,31,22,31,22,30,46,31,177,31,177,30,221,31,143,31,250,31,255,31,253,31,235,31,244,31,97,31,133,31,206,31,193,31,229,31,229,30,229,29,179,31,138,31,93,31,127,31,59,31,52,31,21,31,21,30,21,29,21,28,18,31,18,30,144,31,138,31,161,31,113,31,146,31,150,31,247,31,247,30,228,31,228,30,127,31,127,30,127,29,123,31,123,30,188,31,187,31,107,31,231,31,231,30,231,29,122,31,27,31,143,31,211,31,67,31,39,31,197,31,45,31,35,31,103,31,30,31,80,31,86,31,86,30,86,29,12,31,115,31,67,31,246,31,246,30,18,31,51,31,6,31,6,30,113,31,11,31,140,31,14,31,202,31,90,31,90,30,49,31,49,30,194,31,194,30,55,31,107,31,107,30,87,31,129,31,130,31,142,31,142,30,220,31,17,31,17,30,83,31,98,31,249,31,101,31,101,30,187,31,78,31,147,31,82,31,82,30,141,31,145,31,236,31,236,30,101,31,126,31,1,31,1,30,28,31,163,31,163,30,77,31,80,31,58,31,77,31,39,31,12,31,12,30,12,29,236,31,236,30,23,31,11,31,159,31,124,31,105,31,3,31,72,31,170,31,239,31,155,31,156,31,182,31,132,31,132,30,170,31,170,30,110,31,140,31,30,31,252,31,252,30,128,31,210,31,131,31,144,31,156,31,237,31,30,31,41,31,101,31,231,31,21,31,40,31,40,30,162,31,84,31,108,31,12,31,9,31,233,31,140,31,140,30,232,31,232,30,232,29,210,31,26,31,83,31,236,31,246,31,57,31,60,31,60,30,108,31,248,31,107,31,56,31,165,31,165,30,255,31,184,31,17,31,39,31,39,30,39,29,111,31,111,30,209,31,71,31,71,30,47,31,242,31,242,30,127,31,127,30,97,31,254,31,247,31,247,30,247,29,192,31,194,31,101,31,37,31,188,31,254,31,99,31,81,31,81,30,137,31,192,31,192,30,192,29,248,31,71,31,104,31,209,31,153,31,10,31,23,31,52,31,184,31,145,31,255,31,33,31,33,30,17,31,197,31,209,31,242,31,242,30,29,31,6,31,19,31,159,31,169,31,76,31,42,31,42,30,139,31,7,31,37,31,187,31,187,30,171,31,171,30,18,31,58,31,58,30,58,29,58,28,198,31,10,31,30,31,89,31,85,31,128,31,209,31,80,31,245,31,59,31,119,31,112,31,117,31,243,31,250,31,250,30,188,31,181,31,71,31,255,31,213,31,162,31,92,31,106,31,106,30,208,31,35,31,252,31,58,31,108,31,137,31,210,31,15,31,132,31,132,30,34,31,62,31,126,31,23,31,23,30,33,31,209,31,70,31,70,30,70,29,153,31,147,31,191,31,155,31,155,30,67,31,217,31,217,30,49,31,49,30,73,31,73,30,140,31,196,31,248,31,45,31,219,31,222,31,153,31,218,31,227,31,57,31,102,31,30,31,203,31,176,31,196,31,17,31,17,30,29,31,105,31,216,31,4,31,70,31,64,31,64,31,160,31,206,31,33,31,88,31,66,31,66,30,66,29,66,28,66,27,95,31,95,30,95,29,242,31,242,30,149,31,33,31,219,31,36,31,39,31,39,30,116,31,116,30,83,31,111,31,172,31,18,31,18,30,170,31,203,31,203,30,192,31,139,31,139,30,96,31,96,30,15,31,15,30,203,31,182,31,187,31,136,31,136,30,136,29,50,31,186,31,7,31,214,31,25,31,160,31,2,31,2,30,147,31,26,31,26,30,112,31,49,31,150,31,150,30,150,29,187,31,47,31,104,31,10,31,50,31,245,31,215,31,104,31,214,31,222,31,21,31,21,30,251,31,35,31,36,31,43,31,124,31,124,30,129,31,129,30,218,31,81,31,90,31,142,31,142,30,141,31,165,31,198,31,198,30,133,31,103,31,103,30,76,31,18,31,37,31,189,31,189,30,199,31,57,31,116,31,133,31,133,30,216,31,53,31,76,31,35,31,186,31,106,31,82,31,174,31,118,31,42,31,166,31,112,31,212,31,13,31,83,31,164,31,126,31,102,31,37,31,238,31,132,31,176,31,195,31,3,31,116,31,28,31,202,31,151,31,206,31,206,30,121,31,31,31,228,31,140,31,56,31,62,31,244,31,83,31,170,31,170,30,122,31,122,30,28,31,204,31,85,31,85,30,39,31,186,31,197,31,176,31,72,31,169,31,237,31,238,31,255,31,176,31,147,31,147,30,229,31,154,31,252,31,7,31,82,31,21,31,24,31,199,31,59,31,40,31,225,31,181,31,78,31,229,31,229,30,206,31,51,31,51,30,32,31,10,31,8,31,195,31,132,31,132,30,5,31,202,31,220,31,71,31,238,31,27,31,17,31,101,31,151,31,17,31,224,31,57,31,247,31,247,30,247,29,28,31,69,31,132,31,132,30,132,29,230,31,145,31,145,30,167,31,167,31,53,31,53,30,53,29,233,31,55,31,28,31,132,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
