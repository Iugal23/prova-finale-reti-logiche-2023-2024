-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_769 is
end project_tb_769;

architecture project_tb_arch_769 of project_tb_769 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 872;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,125,0,34,0,29,0,69,0,158,0,167,0,55,0,159,0,223,0,251,0,146,0,189,0,9,0,90,0,0,0,65,0,41,0,217,0,200,0,13,0,220,0,156,0,0,0,4,0,188,0,236,0,0,0,77,0,0,0,254,0,61,0,0,0,204,0,153,0,109,0,161,0,97,0,0,0,0,0,0,0,2,0,92,0,111,0,43,0,73,0,17,0,89,0,158,0,67,0,231,0,170,0,65,0,84,0,255,0,112,0,214,0,235,0,0,0,0,0,146,0,0,0,165,0,86,0,68,0,70,0,214,0,97,0,124,0,237,0,0,0,193,0,0,0,0,0,0,0,0,0,164,0,231,0,31,0,179,0,0,0,0,0,0,0,232,0,0,0,0,0,97,0,47,0,0,0,37,0,213,0,147,0,103,0,46,0,46,0,253,0,163,0,0,0,31,0,64,0,184,0,158,0,29,0,0,0,119,0,181,0,111,0,134,0,57,0,165,0,36,0,162,0,124,0,183,0,0,0,175,0,212,0,15,0,167,0,42,0,100,0,148,0,14,0,231,0,81,0,51,0,24,0,96,0,61,0,70,0,157,0,254,0,236,0,213,0,48,0,0,0,245,0,0,0,34,0,80,0,49,0,67,0,0,0,195,0,127,0,0,0,55,0,236,0,254,0,112,0,117,0,121,0,2,0,198,0,175,0,53,0,148,0,172,0,92,0,16,0,169,0,0,0,90,0,214,0,235,0,175,0,168,0,18,0,0,0,248,0,132,0,0,0,86,0,4,0,59,0,20,0,71,0,218,0,0,0,171,0,0,0,0,0,0,0,52,0,0,0,117,0,0,0,113,0,15,0,26,0,131,0,64,0,61,0,252,0,149,0,139,0,0,0,143,0,0,0,141,0,154,0,42,0,0,0,102,0,0,0,123,0,0,0,114,0,91,0,63,0,227,0,74,0,202,0,40,0,0,0,125,0,65,0,215,0,11,0,195,0,65,0,250,0,53,0,43,0,0,0,206,0,106,0,0,0,181,0,0,0,195,0,5,0,0,0,0,0,212,0,125,0,98,0,0,0,200,0,0,0,129,0,137,0,0,0,0,0,203,0,217,0,164,0,172,0,0,0,0,0,74,0,214,0,229,0,58,0,0,0,128,0,0,0,217,0,195,0,57,0,224,0,60,0,231,0,52,0,30,0,228,0,141,0,71,0,0,0,126,0,158,0,73,0,255,0,133,0,196,0,0,0,72,0,62,0,77,0,239,0,27,0,13,0,238,0,185,0,21,0,88,0,40,0,162,0,183,0,246,0,0,0,0,0,0,0,157,0,0,0,16,0,232,0,194,0,20,0,244,0,0,0,28,0,39,0,30,0,225,0,141,0,170,0,30,0,214,0,69,0,171,0,0,0,49,0,148,0,162,0,201,0,0,0,111,0,171,0,213,0,20,0,60,0,110,0,245,0,17,0,0,0,50,0,58,0,58,0,82,0,69,0,168,0,142,0,0,0,30,0,34,0,0,0,33,0,0,0,242,0,51,0,123,0,180,0,251,0,0,0,94,0,0,0,71,0,59,0,199,0,117,0,35,0,50,0,115,0,120,0,0,0,0,0,0,0,55,0,0,0,15,0,0,0,0,0,133,0,148,0,231,0,0,0,0,0,50,0,0,0,62,0,46,0,13,0,209,0,46,0,182,0,137,0,153,0,51,0,118,0,110,0,214,0,36,0,234,0,0,0,0,0,148,0,25,0,236,0,120,0,213,0,140,0,107,0,0,0,0,0,54,0,216,0,144,0,94,0,250,0,174,0,91,0,134,0,190,0,0,0,196,0,1,0,0,0,0,0,0,0,150,0,74,0,167,0,0,0,56,0,0,0,105,0,43,0,84,0,250,0,36,0,108,0,31,0,139,0,244,0,201,0,195,0,55,0,0,0,26,0,15,0,182,0,29,0,10,0,45,0,191,0,209,0,0,0,71,0,0,0,44,0,190,0,34,0,97,0,153,0,51,0,147,0,0,0,0,0,110,0,224,0,28,0,0,0,15,0,221,0,86,0,98,0,166,0,255,0,0,0,18,0,137,0,164,0,2,0,31,0,120,0,97,0,134,0,0,0,123,0,0,0,74,0,0,0,66,0,187,0,99,0,248,0,114,0,118,0,0,0,214,0,74,0,52,0,0,0,204,0,169,0,90,0,46,0,0,0,36,0,46,0,212,0,2,0,0,0,0,0,159,0,146,0,230,0,0,0,248,0,200,0,253,0,20,0,103,0,57,0,82,0,230,0,0,0,169,0,0,0,225,0,250,0,189,0,92,0,28,0,138,0,109,0,250,0,86,0,0,0,95,0,67,0,79,0,51,0,55,0,188,0,229,0,173,0,0,0,218,0,179,0,0,0,241,0,0,0,160,0,41,0,100,0,55,0,143,0,118,0,189,0,84,0,178,0,215,0,210,0,79,0,112,0,114,0,20,0,0,0,230,0,0,0,23,0,80,0,220,0,202,0,66,0,119,0,0,0,189,0,244,0,136,0,38,0,255,0,5,0,0,0,138,0,8,0,122,0,101,0,0,0,154,0,141,0,0,0,37,0,45,0,237,0,25,0,113,0,0,0,0,0,138,0,123,0,205,0,55,0,154,0,166,0,126,0,33,0,23,0,54,0,21,0,0,0,0,0,121,0,73,0,156,0,127,0,0,0,152,0,195,0,35,0,0,0,223,0,14,0,77,0,162,0,62,0,0,0,193,0,35,0,215,0,0,0,65,0,204,0,178,0,0,0,0,0,0,0,29,0,0,0,53,0,75,0,204,0,168,0,0,0,253,0,14,0,61,0,87,0,160,0,35,0,254,0,0,0,10,0,0,0,195,0,153,0,203,0,175,0,181,0,0,0,214,0,0,0,233,0,69,0,69,0,243,0,120,0,172,0,175,0,18,0,228,0,72,0,11,0,106,0,0,0,0,0,202,0,21,0,238,0,156,0,111,0,59,0,0,0,17,0,158,0,100,0,49,0,0,0,0,0,169,0,0,0,190,0,0,0,0,0,119,0,210,0,109,0,0,0,73,0,42,0,1,0,254,0,208,0,0,0,72,0,97,0,234,0,108,0,77,0,92,0,79,0,154,0,0,0,58,0,0,0,75,0,232,0,0,0,120,0,169,0,228,0,144,0,9,0,125,0,32,0,0,0,138,0,0,0,10,0,149,0,20,0,9,0,0,0,174,0,48,0,178,0,206,0,0,0,238,0,0,0,117,0,182,0,121,0,177,0,174,0,157,0,231,0,95,0,54,0,6,0,144,0,101,0,241,0,0,0,0,0,195,0,0,0,0,0,0,0,74,0,26,0,0,0,0,0,76,0,235,0,230,0,250,0,171,0,49,0,254,0,193,0,170,0,167,0,0,0,187,0,148,0,223,0,35,0,203,0,112,0,82,0,44,0,228,0,0,0,117,0,24,0,35,0,0,0,215,0,201,0,99,0,48,0,0,0,0,0,18,0,191,0,74,0,26,0,42,0,127,0,0,0,31,0,227,0,126,0,71,0,49,0,0,0,125,0,23,0,163,0,70,0,27,0,67,0,120,0,25,0,92,0,0,0,0,0,187,0,0,0,83,0,0,0,178,0,61,0,0,0,214,0,0,0,111,0,85,0,184,0,107,0,225,0,147,0,235,0,27,0,87,0,145,0,162,0,140,0,231,0,3,0,129,0,93,0,187,0,144,0,0,0,173,0,79,0,120,0,94,0,198,0,104,0,131,0,79,0,0,0,0,0,26,0,192,0,191,0,88,0,103,0,240,0,168,0,251,0,162,0,185,0,245,0,222,0,0,0,87,0,13,0,81,0,0,0,0,0,0,0,0,0,135,0,221,0,234,0,0,0,241,0,228,0,167,0,0,0,36,0,215,0,36,0,0,0,88,0,254,0);
signal scenario_full  : scenario_type := (0,0,125,31,34,31,29,31,69,31,158,31,167,31,55,31,159,31,223,31,251,31,146,31,189,31,9,31,90,31,90,30,65,31,41,31,217,31,200,31,13,31,220,31,156,31,156,30,4,31,188,31,236,31,236,30,77,31,77,30,254,31,61,31,61,30,204,31,153,31,109,31,161,31,97,31,97,30,97,29,97,28,2,31,92,31,111,31,43,31,73,31,17,31,89,31,158,31,67,31,231,31,170,31,65,31,84,31,255,31,112,31,214,31,235,31,235,30,235,29,146,31,146,30,165,31,86,31,68,31,70,31,214,31,97,31,124,31,237,31,237,30,193,31,193,30,193,29,193,28,193,27,164,31,231,31,31,31,179,31,179,30,179,29,179,28,232,31,232,30,232,29,97,31,47,31,47,30,37,31,213,31,147,31,103,31,46,31,46,31,253,31,163,31,163,30,31,31,64,31,184,31,158,31,29,31,29,30,119,31,181,31,111,31,134,31,57,31,165,31,36,31,162,31,124,31,183,31,183,30,175,31,212,31,15,31,167,31,42,31,100,31,148,31,14,31,231,31,81,31,51,31,24,31,96,31,61,31,70,31,157,31,254,31,236,31,213,31,48,31,48,30,245,31,245,30,34,31,80,31,49,31,67,31,67,30,195,31,127,31,127,30,55,31,236,31,254,31,112,31,117,31,121,31,2,31,198,31,175,31,53,31,148,31,172,31,92,31,16,31,169,31,169,30,90,31,214,31,235,31,175,31,168,31,18,31,18,30,248,31,132,31,132,30,86,31,4,31,59,31,20,31,71,31,218,31,218,30,171,31,171,30,171,29,171,28,52,31,52,30,117,31,117,30,113,31,15,31,26,31,131,31,64,31,61,31,252,31,149,31,139,31,139,30,143,31,143,30,141,31,154,31,42,31,42,30,102,31,102,30,123,31,123,30,114,31,91,31,63,31,227,31,74,31,202,31,40,31,40,30,125,31,65,31,215,31,11,31,195,31,65,31,250,31,53,31,43,31,43,30,206,31,106,31,106,30,181,31,181,30,195,31,5,31,5,30,5,29,212,31,125,31,98,31,98,30,200,31,200,30,129,31,137,31,137,30,137,29,203,31,217,31,164,31,172,31,172,30,172,29,74,31,214,31,229,31,58,31,58,30,128,31,128,30,217,31,195,31,57,31,224,31,60,31,231,31,52,31,30,31,228,31,141,31,71,31,71,30,126,31,158,31,73,31,255,31,133,31,196,31,196,30,72,31,62,31,77,31,239,31,27,31,13,31,238,31,185,31,21,31,88,31,40,31,162,31,183,31,246,31,246,30,246,29,246,28,157,31,157,30,16,31,232,31,194,31,20,31,244,31,244,30,28,31,39,31,30,31,225,31,141,31,170,31,30,31,214,31,69,31,171,31,171,30,49,31,148,31,162,31,201,31,201,30,111,31,171,31,213,31,20,31,60,31,110,31,245,31,17,31,17,30,50,31,58,31,58,31,82,31,69,31,168,31,142,31,142,30,30,31,34,31,34,30,33,31,33,30,242,31,51,31,123,31,180,31,251,31,251,30,94,31,94,30,71,31,59,31,199,31,117,31,35,31,50,31,115,31,120,31,120,30,120,29,120,28,55,31,55,30,15,31,15,30,15,29,133,31,148,31,231,31,231,30,231,29,50,31,50,30,62,31,46,31,13,31,209,31,46,31,182,31,137,31,153,31,51,31,118,31,110,31,214,31,36,31,234,31,234,30,234,29,148,31,25,31,236,31,120,31,213,31,140,31,107,31,107,30,107,29,54,31,216,31,144,31,94,31,250,31,174,31,91,31,134,31,190,31,190,30,196,31,1,31,1,30,1,29,1,28,150,31,74,31,167,31,167,30,56,31,56,30,105,31,43,31,84,31,250,31,36,31,108,31,31,31,139,31,244,31,201,31,195,31,55,31,55,30,26,31,15,31,182,31,29,31,10,31,45,31,191,31,209,31,209,30,71,31,71,30,44,31,190,31,34,31,97,31,153,31,51,31,147,31,147,30,147,29,110,31,224,31,28,31,28,30,15,31,221,31,86,31,98,31,166,31,255,31,255,30,18,31,137,31,164,31,2,31,31,31,120,31,97,31,134,31,134,30,123,31,123,30,74,31,74,30,66,31,187,31,99,31,248,31,114,31,118,31,118,30,214,31,74,31,52,31,52,30,204,31,169,31,90,31,46,31,46,30,36,31,46,31,212,31,2,31,2,30,2,29,159,31,146,31,230,31,230,30,248,31,200,31,253,31,20,31,103,31,57,31,82,31,230,31,230,30,169,31,169,30,225,31,250,31,189,31,92,31,28,31,138,31,109,31,250,31,86,31,86,30,95,31,67,31,79,31,51,31,55,31,188,31,229,31,173,31,173,30,218,31,179,31,179,30,241,31,241,30,160,31,41,31,100,31,55,31,143,31,118,31,189,31,84,31,178,31,215,31,210,31,79,31,112,31,114,31,20,31,20,30,230,31,230,30,23,31,80,31,220,31,202,31,66,31,119,31,119,30,189,31,244,31,136,31,38,31,255,31,5,31,5,30,138,31,8,31,122,31,101,31,101,30,154,31,141,31,141,30,37,31,45,31,237,31,25,31,113,31,113,30,113,29,138,31,123,31,205,31,55,31,154,31,166,31,126,31,33,31,23,31,54,31,21,31,21,30,21,29,121,31,73,31,156,31,127,31,127,30,152,31,195,31,35,31,35,30,223,31,14,31,77,31,162,31,62,31,62,30,193,31,35,31,215,31,215,30,65,31,204,31,178,31,178,30,178,29,178,28,29,31,29,30,53,31,75,31,204,31,168,31,168,30,253,31,14,31,61,31,87,31,160,31,35,31,254,31,254,30,10,31,10,30,195,31,153,31,203,31,175,31,181,31,181,30,214,31,214,30,233,31,69,31,69,31,243,31,120,31,172,31,175,31,18,31,228,31,72,31,11,31,106,31,106,30,106,29,202,31,21,31,238,31,156,31,111,31,59,31,59,30,17,31,158,31,100,31,49,31,49,30,49,29,169,31,169,30,190,31,190,30,190,29,119,31,210,31,109,31,109,30,73,31,42,31,1,31,254,31,208,31,208,30,72,31,97,31,234,31,108,31,77,31,92,31,79,31,154,31,154,30,58,31,58,30,75,31,232,31,232,30,120,31,169,31,228,31,144,31,9,31,125,31,32,31,32,30,138,31,138,30,10,31,149,31,20,31,9,31,9,30,174,31,48,31,178,31,206,31,206,30,238,31,238,30,117,31,182,31,121,31,177,31,174,31,157,31,231,31,95,31,54,31,6,31,144,31,101,31,241,31,241,30,241,29,195,31,195,30,195,29,195,28,74,31,26,31,26,30,26,29,76,31,235,31,230,31,250,31,171,31,49,31,254,31,193,31,170,31,167,31,167,30,187,31,148,31,223,31,35,31,203,31,112,31,82,31,44,31,228,31,228,30,117,31,24,31,35,31,35,30,215,31,201,31,99,31,48,31,48,30,48,29,18,31,191,31,74,31,26,31,42,31,127,31,127,30,31,31,227,31,126,31,71,31,49,31,49,30,125,31,23,31,163,31,70,31,27,31,67,31,120,31,25,31,92,31,92,30,92,29,187,31,187,30,83,31,83,30,178,31,61,31,61,30,214,31,214,30,111,31,85,31,184,31,107,31,225,31,147,31,235,31,27,31,87,31,145,31,162,31,140,31,231,31,3,31,129,31,93,31,187,31,144,31,144,30,173,31,79,31,120,31,94,31,198,31,104,31,131,31,79,31,79,30,79,29,26,31,192,31,191,31,88,31,103,31,240,31,168,31,251,31,162,31,185,31,245,31,222,31,222,30,87,31,13,31,81,31,81,30,81,29,81,28,81,27,135,31,221,31,234,31,234,30,241,31,228,31,167,31,167,30,36,31,215,31,36,31,36,30,88,31,254,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
