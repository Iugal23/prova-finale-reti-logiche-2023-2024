-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_337 is
end project_tb_337;

architecture project_tb_arch_337 of project_tb_337 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 843;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (186,0,124,0,0,0,201,0,0,0,63,0,154,0,78,0,0,0,28,0,61,0,186,0,255,0,0,0,252,0,14,0,134,0,56,0,115,0,112,0,22,0,31,0,107,0,224,0,167,0,102,0,215,0,53,0,118,0,233,0,176,0,0,0,110,0,137,0,57,0,29,0,0,0,102,0,164,0,0,0,86,0,64,0,42,0,244,0,54,0,117,0,0,0,3,0,36,0,191,0,70,0,253,0,232,0,30,0,157,0,9,0,174,0,0,0,43,0,118,0,111,0,32,0,152,0,61,0,122,0,35,0,61,0,224,0,107,0,65,0,199,0,0,0,13,0,15,0,153,0,254,0,0,0,31,0,225,0,13,0,232,0,203,0,204,0,133,0,129,0,0,0,112,0,134,0,221,0,196,0,65,0,107,0,166,0,66,0,151,0,141,0,233,0,178,0,55,0,48,0,39,0,0,0,14,0,115,0,47,0,0,0,218,0,18,0,0,0,96,0,160,0,0,0,145,0,76,0,21,0,74,0,170,0,97,0,159,0,142,0,72,0,163,0,0,0,198,0,0,0,48,0,125,0,0,0,10,0,0,0,0,0,231,0,35,0,52,0,129,0,178,0,97,0,115,0,0,0,196,0,0,0,139,0,253,0,31,0,101,0,26,0,0,0,23,0,74,0,144,0,62,0,34,0,49,0,221,0,47,0,102,0,25,0,149,0,247,0,112,0,164,0,74,0,23,0,113,0,124,0,58,0,32,0,0,0,169,0,136,0,133,0,33,0,76,0,167,0,38,0,80,0,0,0,69,0,118,0,195,0,179,0,35,0,45,0,64,0,188,0,187,0,192,0,0,0,200,0,186,0,226,0,0,0,0,0,174,0,151,0,87,0,210,0,176,0,137,0,241,0,213,0,73,0,249,0,0,0,0,0,42,0,205,0,8,0,75,0,112,0,3,0,0,0,54,0,204,0,0,0,0,0,252,0,222,0,201,0,0,0,7,0,203,0,0,0,239,0,118,0,11,0,0,0,120,0,195,0,144,0,214,0,148,0,242,0,22,0,71,0,147,0,102,0,127,0,85,0,73,0,0,0,80,0,89,0,67,0,209,0,0,0,204,0,172,0,196,0,83,0,169,0,146,0,108,0,70,0,186,0,215,0,39,0,0,0,171,0,111,0,186,0,0,0,117,0,0,0,5,0,120,0,58,0,208,0,0,0,236,0,0,0,82,0,142,0,194,0,63,0,0,0,51,0,143,0,0,0,33,0,48,0,207,0,0,0,87,0,113,0,104,0,255,0,0,0,211,0,76,0,73,0,0,0,207,0,87,0,14,0,61,0,195,0,109,0,121,0,113,0,108,0,39,0,126,0,19,0,21,0,250,0,0,0,0,0,13,0,111,0,0,0,124,0,152,0,195,0,60,0,106,0,97,0,208,0,0,0,20,0,0,0,194,0,206,0,165,0,208,0,130,0,210,0,248,0,235,0,0,0,166,0,179,0,0,0,110,0,120,0,9,0,0,0,120,0,189,0,151,0,0,0,197,0,112,0,12,0,142,0,13,0,200,0,116,0,249,0,232,0,23,0,0,0,50,0,253,0,220,0,240,0,247,0,197,0,28,0,98,0,221,0,51,0,236,0,68,0,45,0,77,0,114,0,121,0,29,0,0,0,0,0,173,0,130,0,217,0,154,0,0,0,197,0,190,0,220,0,161,0,156,0,241,0,136,0,193,0,191,0,126,0,183,0,201,0,169,0,113,0,39,0,0,0,253,0,34,0,78,0,65,0,0,0,188,0,0,0,160,0,116,0,109,0,0,0,212,0,36,0,160,0,91,0,64,0,211,0,193,0,156,0,178,0,153,0,186,0,164,0,144,0,30,0,237,0,0,0,138,0,167,0,77,0,116,0,63,0,0,0,92,0,231,0,38,0,0,0,25,0,0,0,0,0,130,0,25,0,0,0,167,0,53,0,125,0,0,0,0,0,58,0,0,0,51,0,107,0,0,0,231,0,64,0,244,0,93,0,7,0,208,0,163,0,123,0,216,0,15,0,182,0,60,0,217,0,117,0,35,0,33,0,169,0,221,0,91,0,188,0,189,0,9,0,232,0,245,0,0,0,196,0,0,0,0,0,242,0,193,0,134,0,72,0,247,0,121,0,47,0,0,0,92,0,0,0,242,0,228,0,58,0,143,0,210,0,0,0,0,0,234,0,252,0,218,0,36,0,25,0,143,0,241,0,226,0,52,0,207,0,187,0,229,0,111,0,8,0,0,0,0,0,77,0,194,0,0,0,116,0,197,0,0,0,228,0,59,0,0,0,199,0,0,0,0,0,22,0,135,0,0,0,0,0,72,0,107,0,0,0,0,0,247,0,250,0,139,0,189,0,96,0,75,0,7,0,225,0,57,0,0,0,185,0,158,0,0,0,124,0,81,0,51,0,119,0,0,0,153,0,50,0,0,0,69,0,0,0,27,0,126,0,0,0,112,0,120,0,0,0,62,0,10,0,166,0,0,0,129,0,228,0,7,0,101,0,154,0,46,0,233,0,36,0,153,0,190,0,48,0,124,0,144,0,138,0,0,0,127,0,2,0,212,0,0,0,25,0,157,0,236,0,30,0,14,0,3,0,88,0,158,0,179,0,10,0,27,0,0,0,129,0,112,0,0,0,180,0,0,0,37,0,84,0,0,0,0,0,0,0,110,0,0,0,0,0,106,0,192,0,85,0,124,0,139,0,235,0,123,0,0,0,90,0,139,0,242,0,26,0,7,0,158,0,83,0,0,0,0,0,0,0,252,0,0,0,0,0,179,0,84,0,23,0,0,0,105,0,198,0,11,0,161,0,72,0,158,0,124,0,125,0,212,0,184,0,52,0,174,0,201,0,88,0,253,0,188,0,0,0,246,0,241,0,0,0,84,0,168,0,0,0,123,0,171,0,66,0,117,0,0,0,130,0,106,0,77,0,50,0,134,0,0,0,0,0,0,0,39,0,86,0,0,0,104,0,235,0,180,0,160,0,0,0,127,0,92,0,227,0,0,0,169,0,44,0,23,0,109,0,0,0,227,0,0,0,94,0,209,0,234,0,54,0,139,0,245,0,245,0,0,0,35,0,18,0,0,0,234,0,146,0,60,0,162,0,0,0,124,0,100,0,232,0,0,0,0,0,93,0,179,0,58,0,55,0,0,0,153,0,107,0,101,0,0,0,0,0,211,0,190,0,186,0,0,0,29,0,0,0,153,0,150,0,36,0,124,0,237,0,16,0,241,0,196,0,247,0,91,0,213,0,194,0,215,0,188,0,0,0,21,0,155,0,0,0,125,0,200,0,190,0,113,0,120,0,90,0,0,0,0,0,226,0,124,0,189,0,96,0,96,0,0,0,60,0,236,0,0,0,217,0,221,0,0,0,0,0,127,0,184,0,17,0,137,0,45,0,44,0,66,0,53,0,109,0,52,0,0,0,77,0,0,0,141,0,223,0,1,0,178,0,223,0,97,0,121,0,210,0,24,0,193,0,183,0,84,0,115,0,141,0,0,0,221,0,0,0,29,0,236,0,226,0,155,0,166,0,0,0,149,0,227,0,69,0,54,0,80,0,0,0,54,0,184,0,4,0,139,0,101,0,127,0,49,0,43,0,142,0,0,0,238,0,132,0,210,0,251,0,73,0,52,0,179,0,85,0,68,0,132,0,34,0,204,0,76,0,0,0,161,0,9,0,88,0,126,0,255,0,0,0,0,0,31,0,0,0,182,0,21,0,113,0,121,0,147,0,1,0,34,0,122,0,107,0);
signal scenario_full  : scenario_type := (186,31,124,31,124,30,201,31,201,30,63,31,154,31,78,31,78,30,28,31,61,31,186,31,255,31,255,30,252,31,14,31,134,31,56,31,115,31,112,31,22,31,31,31,107,31,224,31,167,31,102,31,215,31,53,31,118,31,233,31,176,31,176,30,110,31,137,31,57,31,29,31,29,30,102,31,164,31,164,30,86,31,64,31,42,31,244,31,54,31,117,31,117,30,3,31,36,31,191,31,70,31,253,31,232,31,30,31,157,31,9,31,174,31,174,30,43,31,118,31,111,31,32,31,152,31,61,31,122,31,35,31,61,31,224,31,107,31,65,31,199,31,199,30,13,31,15,31,153,31,254,31,254,30,31,31,225,31,13,31,232,31,203,31,204,31,133,31,129,31,129,30,112,31,134,31,221,31,196,31,65,31,107,31,166,31,66,31,151,31,141,31,233,31,178,31,55,31,48,31,39,31,39,30,14,31,115,31,47,31,47,30,218,31,18,31,18,30,96,31,160,31,160,30,145,31,76,31,21,31,74,31,170,31,97,31,159,31,142,31,72,31,163,31,163,30,198,31,198,30,48,31,125,31,125,30,10,31,10,30,10,29,231,31,35,31,52,31,129,31,178,31,97,31,115,31,115,30,196,31,196,30,139,31,253,31,31,31,101,31,26,31,26,30,23,31,74,31,144,31,62,31,34,31,49,31,221,31,47,31,102,31,25,31,149,31,247,31,112,31,164,31,74,31,23,31,113,31,124,31,58,31,32,31,32,30,169,31,136,31,133,31,33,31,76,31,167,31,38,31,80,31,80,30,69,31,118,31,195,31,179,31,35,31,45,31,64,31,188,31,187,31,192,31,192,30,200,31,186,31,226,31,226,30,226,29,174,31,151,31,87,31,210,31,176,31,137,31,241,31,213,31,73,31,249,31,249,30,249,29,42,31,205,31,8,31,75,31,112,31,3,31,3,30,54,31,204,31,204,30,204,29,252,31,222,31,201,31,201,30,7,31,203,31,203,30,239,31,118,31,11,31,11,30,120,31,195,31,144,31,214,31,148,31,242,31,22,31,71,31,147,31,102,31,127,31,85,31,73,31,73,30,80,31,89,31,67,31,209,31,209,30,204,31,172,31,196,31,83,31,169,31,146,31,108,31,70,31,186,31,215,31,39,31,39,30,171,31,111,31,186,31,186,30,117,31,117,30,5,31,120,31,58,31,208,31,208,30,236,31,236,30,82,31,142,31,194,31,63,31,63,30,51,31,143,31,143,30,33,31,48,31,207,31,207,30,87,31,113,31,104,31,255,31,255,30,211,31,76,31,73,31,73,30,207,31,87,31,14,31,61,31,195,31,109,31,121,31,113,31,108,31,39,31,126,31,19,31,21,31,250,31,250,30,250,29,13,31,111,31,111,30,124,31,152,31,195,31,60,31,106,31,97,31,208,31,208,30,20,31,20,30,194,31,206,31,165,31,208,31,130,31,210,31,248,31,235,31,235,30,166,31,179,31,179,30,110,31,120,31,9,31,9,30,120,31,189,31,151,31,151,30,197,31,112,31,12,31,142,31,13,31,200,31,116,31,249,31,232,31,23,31,23,30,50,31,253,31,220,31,240,31,247,31,197,31,28,31,98,31,221,31,51,31,236,31,68,31,45,31,77,31,114,31,121,31,29,31,29,30,29,29,173,31,130,31,217,31,154,31,154,30,197,31,190,31,220,31,161,31,156,31,241,31,136,31,193,31,191,31,126,31,183,31,201,31,169,31,113,31,39,31,39,30,253,31,34,31,78,31,65,31,65,30,188,31,188,30,160,31,116,31,109,31,109,30,212,31,36,31,160,31,91,31,64,31,211,31,193,31,156,31,178,31,153,31,186,31,164,31,144,31,30,31,237,31,237,30,138,31,167,31,77,31,116,31,63,31,63,30,92,31,231,31,38,31,38,30,25,31,25,30,25,29,130,31,25,31,25,30,167,31,53,31,125,31,125,30,125,29,58,31,58,30,51,31,107,31,107,30,231,31,64,31,244,31,93,31,7,31,208,31,163,31,123,31,216,31,15,31,182,31,60,31,217,31,117,31,35,31,33,31,169,31,221,31,91,31,188,31,189,31,9,31,232,31,245,31,245,30,196,31,196,30,196,29,242,31,193,31,134,31,72,31,247,31,121,31,47,31,47,30,92,31,92,30,242,31,228,31,58,31,143,31,210,31,210,30,210,29,234,31,252,31,218,31,36,31,25,31,143,31,241,31,226,31,52,31,207,31,187,31,229,31,111,31,8,31,8,30,8,29,77,31,194,31,194,30,116,31,197,31,197,30,228,31,59,31,59,30,199,31,199,30,199,29,22,31,135,31,135,30,135,29,72,31,107,31,107,30,107,29,247,31,250,31,139,31,189,31,96,31,75,31,7,31,225,31,57,31,57,30,185,31,158,31,158,30,124,31,81,31,51,31,119,31,119,30,153,31,50,31,50,30,69,31,69,30,27,31,126,31,126,30,112,31,120,31,120,30,62,31,10,31,166,31,166,30,129,31,228,31,7,31,101,31,154,31,46,31,233,31,36,31,153,31,190,31,48,31,124,31,144,31,138,31,138,30,127,31,2,31,212,31,212,30,25,31,157,31,236,31,30,31,14,31,3,31,88,31,158,31,179,31,10,31,27,31,27,30,129,31,112,31,112,30,180,31,180,30,37,31,84,31,84,30,84,29,84,28,110,31,110,30,110,29,106,31,192,31,85,31,124,31,139,31,235,31,123,31,123,30,90,31,139,31,242,31,26,31,7,31,158,31,83,31,83,30,83,29,83,28,252,31,252,30,252,29,179,31,84,31,23,31,23,30,105,31,198,31,11,31,161,31,72,31,158,31,124,31,125,31,212,31,184,31,52,31,174,31,201,31,88,31,253,31,188,31,188,30,246,31,241,31,241,30,84,31,168,31,168,30,123,31,171,31,66,31,117,31,117,30,130,31,106,31,77,31,50,31,134,31,134,30,134,29,134,28,39,31,86,31,86,30,104,31,235,31,180,31,160,31,160,30,127,31,92,31,227,31,227,30,169,31,44,31,23,31,109,31,109,30,227,31,227,30,94,31,209,31,234,31,54,31,139,31,245,31,245,31,245,30,35,31,18,31,18,30,234,31,146,31,60,31,162,31,162,30,124,31,100,31,232,31,232,30,232,29,93,31,179,31,58,31,55,31,55,30,153,31,107,31,101,31,101,30,101,29,211,31,190,31,186,31,186,30,29,31,29,30,153,31,150,31,36,31,124,31,237,31,16,31,241,31,196,31,247,31,91,31,213,31,194,31,215,31,188,31,188,30,21,31,155,31,155,30,125,31,200,31,190,31,113,31,120,31,90,31,90,30,90,29,226,31,124,31,189,31,96,31,96,31,96,30,60,31,236,31,236,30,217,31,221,31,221,30,221,29,127,31,184,31,17,31,137,31,45,31,44,31,66,31,53,31,109,31,52,31,52,30,77,31,77,30,141,31,223,31,1,31,178,31,223,31,97,31,121,31,210,31,24,31,193,31,183,31,84,31,115,31,141,31,141,30,221,31,221,30,29,31,236,31,226,31,155,31,166,31,166,30,149,31,227,31,69,31,54,31,80,31,80,30,54,31,184,31,4,31,139,31,101,31,127,31,49,31,43,31,142,31,142,30,238,31,132,31,210,31,251,31,73,31,52,31,179,31,85,31,68,31,132,31,34,31,204,31,76,31,76,30,161,31,9,31,88,31,126,31,255,31,255,30,255,29,31,31,31,30,182,31,21,31,113,31,121,31,147,31,1,31,34,31,122,31,107,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
