-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_565 is
end project_tb_565;

architecture project_tb_arch_565 of project_tb_565 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 981;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (0,0,0,0,36,0,12,0,190,0,155,0,47,0,0,0,76,0,137,0,7,0,120,0,0,0,14,0,0,0,0,0,192,0,223,0,68,0,120,0,28,0,236,0,0,0,156,0,0,0,39,0,21,0,29,0,234,0,168,0,150,0,47,0,221,0,27,0,233,0,0,0,8,0,204,0,176,0,0,0,48,0,109,0,220,0,96,0,126,0,62,0,0,0,201,0,50,0,141,0,203,0,94,0,206,0,2,0,164,0,0,0,112,0,28,0,174,0,254,0,42,0,84,0,224,0,137,0,0,0,243,0,160,0,0,0,116,0,251,0,0,0,208,0,216,0,204,0,181,0,147,0,40,0,250,0,99,0,211,0,5,0,241,0,41,0,223,0,228,0,232,0,0,0,222,0,240,0,4,0,169,0,0,0,224,0,44,0,0,0,0,0,179,0,186,0,138,0,140,0,68,0,120,0,65,0,179,0,250,0,227,0,0,0,244,0,2,0,239,0,121,0,129,0,163,0,140,0,218,0,0,0,144,0,61,0,163,0,0,0,5,0,32,0,0,0,13,0,0,0,196,0,0,0,120,0,106,0,240,0,36,0,124,0,0,0,11,0,20,0,0,0,39,0,125,0,220,0,50,0,22,0,0,0,118,0,232,0,114,0,200,0,252,0,103,0,88,0,0,0,210,0,71,0,250,0,0,0,0,0,0,0,185,0,245,0,145,0,6,0,0,0,33,0,0,0,229,0,0,0,250,0,250,0,142,0,95,0,199,0,22,0,24,0,194,0,150,0,59,0,36,0,173,0,108,0,96,0,29,0,11,0,29,0,207,0,102,0,30,0,219,0,7,0,0,0,163,0,0,0,78,0,70,0,29,0,0,0,108,0,69,0,21,0,0,0,79,0,203,0,56,0,122,0,0,0,202,0,204,0,177,0,0,0,109,0,31,0,196,0,233,0,103,0,186,0,80,0,47,0,93,0,230,0,196,0,15,0,216,0,129,0,32,0,0,0,0,0,77,0,243,0,65,0,37,0,171,0,202,0,82,0,10,0,191,0,107,0,186,0,54,0,150,0,240,0,176,0,195,0,211,0,0,0,216,0,105,0,153,0,0,0,95,0,144,0,113,0,48,0,95,0,49,0,201,0,200,0,187,0,98,0,163,0,181,0,113,0,6,0,107,0,26,0,20,0,29,0,156,0,0,0,113,0,97,0,80,0,0,0,248,0,37,0,0,0,0,0,190,0,19,0,54,0,182,0,0,0,6,0,152,0,226,0,182,0,30,0,0,0,5,0,197,0,22,0,151,0,105,0,0,0,233,0,253,0,0,0,0,0,0,0,133,0,65,0,0,0,108,0,183,0,232,0,177,0,5,0,12,0,55,0,0,0,0,0,0,0,0,0,164,0,66,0,205,0,23,0,55,0,0,0,202,0,0,0,93,0,51,0,220,0,168,0,63,0,45,0,33,0,252,0,0,0,165,0,186,0,243,0,0,0,105,0,33,0,19,0,125,0,0,0,30,0,0,0,193,0,0,0,22,0,0,0,215,0,211,0,201,0,97,0,127,0,14,0,101,0,0,0,86,0,201,0,71,0,119,0,0,0,84,0,7,0,112,0,14,0,228,0,0,0,0,0,210,0,51,0,143,0,57,0,0,0,49,0,179,0,167,0,77,0,0,0,0,0,72,0,11,0,247,0,24,0,8,0,174,0,216,0,204,0,187,0,177,0,0,0,0,0,106,0,198,0,42,0,0,0,124,0,151,0,199,0,99,0,132,0,0,0,230,0,239,0,0,0,109,0,15,0,97,0,80,0,65,0,47,0,0,0,60,0,223,0,0,0,158,0,161,0,80,0,213,0,237,0,0,0,237,0,163,0,33,0,0,0,0,0,189,0,17,0,131,0,68,0,0,0,0,0,94,0,0,0,8,0,166,0,84,0,178,0,0,0,115,0,0,0,243,0,118,0,94,0,222,0,23,0,0,0,0,0,71,0,0,0,246,0,168,0,91,0,214,0,176,0,11,0,173,0,190,0,148,0,0,0,0,0,254,0,111,0,124,0,37,0,189,0,111,0,158,0,107,0,0,0,54,0,225,0,164,0,250,0,84,0,0,0,47,0,223,0,11,0,200,0,102,0,162,0,0,0,221,0,18,0,212,0,130,0,231,0,0,0,128,0,237,0,0,0,143,0,0,0,65,0,253,0,185,0,125,0,0,0,0,0,138,0,38,0,0,0,86,0,166,0,203,0,208,0,67,0,0,0,4,0,205,0,0,0,229,0,59,0,70,0,119,0,89,0,74,0,0,0,213,0,127,0,73,0,126,0,0,0,0,0,119,0,36,0,145,0,7,0,1,0,76,0,88,0,136,0,190,0,100,0,209,0,124,0,83,0,52,0,97,0,218,0,184,0,35,0,196,0,130,0,5,0,0,0,23,0,15,0,0,0,180,0,8,0,0,0,0,0,64,0,0,0,0,0,33,0,31,0,139,0,253,0,8,0,166,0,248,0,4,0,113,0,33,0,150,0,233,0,169,0,46,0,169,0,191,0,34,0,0,0,0,0,5,0,4,0,195,0,165,0,141,0,149,0,0,0,226,0,0,0,190,0,121,0,0,0,253,0,164,0,0,0,67,0,222,0,235,0,249,0,0,0,1,0,50,0,10,0,140,0,142,0,199,0,160,0,92,0,154,0,0,0,117,0,0,0,108,0,191,0,162,0,232,0,54,0,191,0,165,0,104,0,165,0,211,0,0,0,105,0,189,0,0,0,44,0,160,0,104,0,102,0,225,0,6,0,0,0,190,0,40,0,45,0,211,0,16,0,84,0,94,0,232,0,0,0,71,0,121,0,0,0,215,0,85,0,169,0,0,0,0,0,160,0,71,0,157,0,235,0,157,0,100,0,0,0,250,0,33,0,42,0,94,0,42,0,0,0,212,0,84,0,84,0,33,0,16,0,0,0,230,0,153,0,57,0,245,0,178,0,121,0,165,0,104,0,0,0,22,0,23,0,81,0,243,0,207,0,5,0,170,0,162,0,70,0,0,0,140,0,246,0,54,0,245,0,11,0,255,0,50,0,161,0,163,0,230,0,251,0,0,0,19,0,0,0,106,0,73,0,12,0,68,0,62,0,133,0,57,0,91,0,80,0,26,0,230,0,249,0,43,0,225,0,236,0,0,0,0,0,76,0,178,0,0,0,93,0,215,0,83,0,158,0,142,0,0,0,71,0,78,0,0,0,0,0,95,0,57,0,17,0,46,0,44,0,0,0,68,0,198,0,78,0,247,0,99,0,12,0,205,0,178,0,125,0,107,0,33,0,241,0,61,0,66,0,104,0,173,0,245,0,26,0,134,0,205,0,28,0,160,0,155,0,30,0,0,0,0,0,55,0,0,0,0,0,125,0,208,0,0,0,202,0,107,0,146,0,34,0,0,0,200,0,180,0,74,0,0,0,60,0,68,0,81,0,213,0,0,0,178,0,90,0,223,0,254,0,84,0,166,0,198,0,41,0,136,0,246,0,0,0,121,0,205,0,0,0,244,0,122,0,122,0,103,0,64,0,152,0,68,0,82,0,0,0,0,0,57,0,0,0,242,0,152,0,250,0,230,0,190,0,230,0,29,0,0,0,73,0,5,0,236,0,51,0,0,0,0,0,68,0,199,0,165,0,252,0,37,0,27,0,49,0,0,0,70,0,0,0,0,0,129,0,209,0,197,0,30,0,17,0,142,0,253,0,21,0,72,0,24,0,23,0,255,0,252,0,0,0,46,0,168,0,168,0,6,0,250,0,0,0,27,0,218,0,141,0,247,0,63,0,0,0,72,0,8,0,221,0,19,0,0,0,48,0,0,0,207,0,106,0,66,0,146,0,0,0,54,0,149,0,96,0,67,0,18,0,246,0,64,0,177,0,163,0,221,0,0,0,25,0,0,0,45,0,107,0,0,0,21,0,0,0,93,0,0,0,62,0,166,0,47,0,0,0,40,0,118,0,75,0,5,0,0,0,162,0,212,0,0,0,0,0,82,0,234,0,112,0,108,0,45,0,190,0,210,0,99,0,215,0,234,0,136,0,33,0,239,0,74,0,171,0,0,0,242,0,48,0,0,0,101,0,115,0,72,0,73,0,125,0,0,0,248,0,0,0,0,0,152,0,226,0,155,0,17,0,84,0,199,0,85,0,42,0,0,0,227,0,197,0,252,0,81,0,0,0,176,0,8,0,123,0,103,0,224,0,57,0,94,0,133,0,0,0,0,0,149,0,201,0,16,0,46,0,27,0,217,0,162,0,13,0,29,0,0,0,80,0,161,0,0,0,0,0,37,0,166,0,83,0,201,0,0,0,212,0,52,0,0,0,253,0,0,0,92,0,17,0,28,0,54,0,113,0,36,0,0,0,161,0,34,0,99,0);
signal scenario_full  : scenario_type := (0,0,0,0,36,31,12,31,190,31,155,31,47,31,47,30,76,31,137,31,7,31,120,31,120,30,14,31,14,30,14,29,192,31,223,31,68,31,120,31,28,31,236,31,236,30,156,31,156,30,39,31,21,31,29,31,234,31,168,31,150,31,47,31,221,31,27,31,233,31,233,30,8,31,204,31,176,31,176,30,48,31,109,31,220,31,96,31,126,31,62,31,62,30,201,31,50,31,141,31,203,31,94,31,206,31,2,31,164,31,164,30,112,31,28,31,174,31,254,31,42,31,84,31,224,31,137,31,137,30,243,31,160,31,160,30,116,31,251,31,251,30,208,31,216,31,204,31,181,31,147,31,40,31,250,31,99,31,211,31,5,31,241,31,41,31,223,31,228,31,232,31,232,30,222,31,240,31,4,31,169,31,169,30,224,31,44,31,44,30,44,29,179,31,186,31,138,31,140,31,68,31,120,31,65,31,179,31,250,31,227,31,227,30,244,31,2,31,239,31,121,31,129,31,163,31,140,31,218,31,218,30,144,31,61,31,163,31,163,30,5,31,32,31,32,30,13,31,13,30,196,31,196,30,120,31,106,31,240,31,36,31,124,31,124,30,11,31,20,31,20,30,39,31,125,31,220,31,50,31,22,31,22,30,118,31,232,31,114,31,200,31,252,31,103,31,88,31,88,30,210,31,71,31,250,31,250,30,250,29,250,28,185,31,245,31,145,31,6,31,6,30,33,31,33,30,229,31,229,30,250,31,250,31,142,31,95,31,199,31,22,31,24,31,194,31,150,31,59,31,36,31,173,31,108,31,96,31,29,31,11,31,29,31,207,31,102,31,30,31,219,31,7,31,7,30,163,31,163,30,78,31,70,31,29,31,29,30,108,31,69,31,21,31,21,30,79,31,203,31,56,31,122,31,122,30,202,31,204,31,177,31,177,30,109,31,31,31,196,31,233,31,103,31,186,31,80,31,47,31,93,31,230,31,196,31,15,31,216,31,129,31,32,31,32,30,32,29,77,31,243,31,65,31,37,31,171,31,202,31,82,31,10,31,191,31,107,31,186,31,54,31,150,31,240,31,176,31,195,31,211,31,211,30,216,31,105,31,153,31,153,30,95,31,144,31,113,31,48,31,95,31,49,31,201,31,200,31,187,31,98,31,163,31,181,31,113,31,6,31,107,31,26,31,20,31,29,31,156,31,156,30,113,31,97,31,80,31,80,30,248,31,37,31,37,30,37,29,190,31,19,31,54,31,182,31,182,30,6,31,152,31,226,31,182,31,30,31,30,30,5,31,197,31,22,31,151,31,105,31,105,30,233,31,253,31,253,30,253,29,253,28,133,31,65,31,65,30,108,31,183,31,232,31,177,31,5,31,12,31,55,31,55,30,55,29,55,28,55,27,164,31,66,31,205,31,23,31,55,31,55,30,202,31,202,30,93,31,51,31,220,31,168,31,63,31,45,31,33,31,252,31,252,30,165,31,186,31,243,31,243,30,105,31,33,31,19,31,125,31,125,30,30,31,30,30,193,31,193,30,22,31,22,30,215,31,211,31,201,31,97,31,127,31,14,31,101,31,101,30,86,31,201,31,71,31,119,31,119,30,84,31,7,31,112,31,14,31,228,31,228,30,228,29,210,31,51,31,143,31,57,31,57,30,49,31,179,31,167,31,77,31,77,30,77,29,72,31,11,31,247,31,24,31,8,31,174,31,216,31,204,31,187,31,177,31,177,30,177,29,106,31,198,31,42,31,42,30,124,31,151,31,199,31,99,31,132,31,132,30,230,31,239,31,239,30,109,31,15,31,97,31,80,31,65,31,47,31,47,30,60,31,223,31,223,30,158,31,161,31,80,31,213,31,237,31,237,30,237,31,163,31,33,31,33,30,33,29,189,31,17,31,131,31,68,31,68,30,68,29,94,31,94,30,8,31,166,31,84,31,178,31,178,30,115,31,115,30,243,31,118,31,94,31,222,31,23,31,23,30,23,29,71,31,71,30,246,31,168,31,91,31,214,31,176,31,11,31,173,31,190,31,148,31,148,30,148,29,254,31,111,31,124,31,37,31,189,31,111,31,158,31,107,31,107,30,54,31,225,31,164,31,250,31,84,31,84,30,47,31,223,31,11,31,200,31,102,31,162,31,162,30,221,31,18,31,212,31,130,31,231,31,231,30,128,31,237,31,237,30,143,31,143,30,65,31,253,31,185,31,125,31,125,30,125,29,138,31,38,31,38,30,86,31,166,31,203,31,208,31,67,31,67,30,4,31,205,31,205,30,229,31,59,31,70,31,119,31,89,31,74,31,74,30,213,31,127,31,73,31,126,31,126,30,126,29,119,31,36,31,145,31,7,31,1,31,76,31,88,31,136,31,190,31,100,31,209,31,124,31,83,31,52,31,97,31,218,31,184,31,35,31,196,31,130,31,5,31,5,30,23,31,15,31,15,30,180,31,8,31,8,30,8,29,64,31,64,30,64,29,33,31,31,31,139,31,253,31,8,31,166,31,248,31,4,31,113,31,33,31,150,31,233,31,169,31,46,31,169,31,191,31,34,31,34,30,34,29,5,31,4,31,195,31,165,31,141,31,149,31,149,30,226,31,226,30,190,31,121,31,121,30,253,31,164,31,164,30,67,31,222,31,235,31,249,31,249,30,1,31,50,31,10,31,140,31,142,31,199,31,160,31,92,31,154,31,154,30,117,31,117,30,108,31,191,31,162,31,232,31,54,31,191,31,165,31,104,31,165,31,211,31,211,30,105,31,189,31,189,30,44,31,160,31,104,31,102,31,225,31,6,31,6,30,190,31,40,31,45,31,211,31,16,31,84,31,94,31,232,31,232,30,71,31,121,31,121,30,215,31,85,31,169,31,169,30,169,29,160,31,71,31,157,31,235,31,157,31,100,31,100,30,250,31,33,31,42,31,94,31,42,31,42,30,212,31,84,31,84,31,33,31,16,31,16,30,230,31,153,31,57,31,245,31,178,31,121,31,165,31,104,31,104,30,22,31,23,31,81,31,243,31,207,31,5,31,170,31,162,31,70,31,70,30,140,31,246,31,54,31,245,31,11,31,255,31,50,31,161,31,163,31,230,31,251,31,251,30,19,31,19,30,106,31,73,31,12,31,68,31,62,31,133,31,57,31,91,31,80,31,26,31,230,31,249,31,43,31,225,31,236,31,236,30,236,29,76,31,178,31,178,30,93,31,215,31,83,31,158,31,142,31,142,30,71,31,78,31,78,30,78,29,95,31,57,31,17,31,46,31,44,31,44,30,68,31,198,31,78,31,247,31,99,31,12,31,205,31,178,31,125,31,107,31,33,31,241,31,61,31,66,31,104,31,173,31,245,31,26,31,134,31,205,31,28,31,160,31,155,31,30,31,30,30,30,29,55,31,55,30,55,29,125,31,208,31,208,30,202,31,107,31,146,31,34,31,34,30,200,31,180,31,74,31,74,30,60,31,68,31,81,31,213,31,213,30,178,31,90,31,223,31,254,31,84,31,166,31,198,31,41,31,136,31,246,31,246,30,121,31,205,31,205,30,244,31,122,31,122,31,103,31,64,31,152,31,68,31,82,31,82,30,82,29,57,31,57,30,242,31,152,31,250,31,230,31,190,31,230,31,29,31,29,30,73,31,5,31,236,31,51,31,51,30,51,29,68,31,199,31,165,31,252,31,37,31,27,31,49,31,49,30,70,31,70,30,70,29,129,31,209,31,197,31,30,31,17,31,142,31,253,31,21,31,72,31,24,31,23,31,255,31,252,31,252,30,46,31,168,31,168,31,6,31,250,31,250,30,27,31,218,31,141,31,247,31,63,31,63,30,72,31,8,31,221,31,19,31,19,30,48,31,48,30,207,31,106,31,66,31,146,31,146,30,54,31,149,31,96,31,67,31,18,31,246,31,64,31,177,31,163,31,221,31,221,30,25,31,25,30,45,31,107,31,107,30,21,31,21,30,93,31,93,30,62,31,166,31,47,31,47,30,40,31,118,31,75,31,5,31,5,30,162,31,212,31,212,30,212,29,82,31,234,31,112,31,108,31,45,31,190,31,210,31,99,31,215,31,234,31,136,31,33,31,239,31,74,31,171,31,171,30,242,31,48,31,48,30,101,31,115,31,72,31,73,31,125,31,125,30,248,31,248,30,248,29,152,31,226,31,155,31,17,31,84,31,199,31,85,31,42,31,42,30,227,31,197,31,252,31,81,31,81,30,176,31,8,31,123,31,103,31,224,31,57,31,94,31,133,31,133,30,133,29,149,31,201,31,16,31,46,31,27,31,217,31,162,31,13,31,29,31,29,30,80,31,161,31,161,30,161,29,37,31,166,31,83,31,201,31,201,30,212,31,52,31,52,30,253,31,253,30,92,31,17,31,28,31,54,31,113,31,36,31,36,30,161,31,34,31,99,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
