-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_474 is
end project_tb_474;

architecture project_tb_arch_474 of project_tb_474 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 535;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (14,0,221,0,31,0,33,0,157,0,236,0,0,0,110,0,181,0,92,0,131,0,2,0,73,0,21,0,18,0,61,0,0,0,183,0,0,0,0,0,161,0,206,0,0,0,53,0,142,0,232,0,133,0,0,0,143,0,112,0,0,0,181,0,142,0,43,0,0,0,58,0,220,0,19,0,148,0,91,0,19,0,225,0,31,0,255,0,107,0,146,0,52,0,136,0,79,0,215,0,146,0,13,0,110,0,96,0,120,0,0,0,179,0,193,0,183,0,0,0,191,0,23,0,14,0,111,0,171,0,0,0,0,0,44,0,118,0,0,0,126,0,153,0,237,0,0,0,237,0,29,0,116,0,125,0,235,0,201,0,133,0,11,0,12,0,77,0,0,0,62,0,201,0,0,0,0,0,200,0,40,0,197,0,117,0,150,0,203,0,23,0,82,0,119,0,56,0,105,0,0,0,165,0,124,0,0,0,0,0,176,0,0,0,90,0,40,0,192,0,0,0,58,0,0,0,219,0,24,0,0,0,33,0,219,0,233,0,217,0,67,0,0,0,166,0,217,0,39,0,34,0,11,0,74,0,161,0,173,0,39,0,159,0,233,0,142,0,82,0,0,0,204,0,28,0,98,0,234,0,249,0,29,0,0,0,35,0,0,0,198,0,212,0,0,0,236,0,42,0,204,0,186,0,84,0,173,0,96,0,0,0,143,0,100,0,207,0,83,0,113,0,31,0,0,0,0,0,188,0,234,0,82,0,2,0,22,0,133,0,0,0,0,0,111,0,250,0,1,0,149,0,130,0,159,0,197,0,102,0,0,0,182,0,227,0,169,0,224,0,128,0,69,0,100,0,31,0,136,0,28,0,142,0,159,0,0,0,0,0,0,0,131,0,241,0,169,0,111,0,209,0,75,0,39,0,240,0,0,0,12,0,0,0,0,0,18,0,55,0,66,0,0,0,81,0,13,0,7,0,42,0,52,0,8,0,212,0,91,0,111,0,3,0,44,0,176,0,133,0,70,0,0,0,105,0,138,0,64,0,61,0,25,0,108,0,247,0,148,0,0,0,143,0,104,0,196,0,129,0,106,0,0,0,119,0,0,0,46,0,174,0,24,0,0,0,59,0,255,0,6,0,89,0,6,0,0,0,93,0,122,0,0,0,0,0,218,0,152,0,22,0,125,0,145,0,61,0,72,0,112,0,175,0,189,0,0,0,198,0,193,0,156,0,0,0,248,0,15,0,0,0,0,0,0,0,240,0,173,0,31,0,1,0,0,0,0,0,50,0,48,0,0,0,137,0,39,0,234,0,23,0,195,0,0,0,0,0,41,0,191,0,192,0,30,0,0,0,239,0,111,0,171,0,0,0,43,0,0,0,35,0,217,0,124,0,96,0,23,0,135,0,194,0,0,0,48,0,0,0,233,0,205,0,0,0,0,0,116,0,229,0,0,0,228,0,228,0,244,0,125,0,156,0,249,0,53,0,58,0,0,0,70,0,138,0,185,0,235,0,173,0,166,0,143,0,94,0,250,0,199,0,53,0,141,0,235,0,64,0,0,0,22,0,0,0,69,0,0,0,168,0,113,0,79,0,195,0,229,0,68,0,255,0,0,0,0,0,60,0,228,0,143,0,0,0,22,0,150,0,139,0,154,0,1,0,125,0,84,0,0,0,143,0,0,0,199,0,86,0,56,0,0,0,137,0,221,0,126,0,67,0,227,0,190,0,249,0,188,0,80,0,171,0,45,0,47,0,180,0,191,0,102,0,162,0,0,0,159,0,101,0,71,0,0,0,229,0,54,0,43,0,0,0,200,0,0,0,0,0,159,0,106,0,39,0,169,0,86,0,0,0,53,0,149,0,90,0,147,0,111,0,200,0,93,0,0,0,48,0,110,0,152,0,13,0,83,0,186,0,0,0,255,0,171,0,101,0,97,0,12,0,0,0,185,0,0,0,0,0,26,0,0,0,225,0,177,0,203,0,141,0,0,0,69,0,2,0,0,0,147,0,19,0,0,0,39,0,217,0,67,0,59,0,0,0,197,0,207,0,234,0,71,0,60,0,17,0,152,0,67,0,211,0,161,0,211,0,21,0,76,0,205,0,0,0,192,0,0,0,66,0,171,0,197,0,196,0,120,0,159,0,34,0,161,0,240,0,104,0,26,0,13,0,161,0,0,0,80,0,0,0,169,0,109,0,182,0,216,0,109,0,192,0,132,0,249,0,4,0,0,0,227,0,0,0,15,0,162,0,48,0,232,0,236,0,0,0,179,0,111,0,46,0,199,0,7,0,171,0,219,0,198,0,91,0,72,0,103,0,239,0,246,0,117,0,140,0,0,0,101,0,0,0,35,0,71,0,185,0,118,0,121,0,195,0,237,0,104,0,165,0,241,0,65,0,44,0,75,0);
signal scenario_full  : scenario_type := (14,31,221,31,31,31,33,31,157,31,236,31,236,30,110,31,181,31,92,31,131,31,2,31,73,31,21,31,18,31,61,31,61,30,183,31,183,30,183,29,161,31,206,31,206,30,53,31,142,31,232,31,133,31,133,30,143,31,112,31,112,30,181,31,142,31,43,31,43,30,58,31,220,31,19,31,148,31,91,31,19,31,225,31,31,31,255,31,107,31,146,31,52,31,136,31,79,31,215,31,146,31,13,31,110,31,96,31,120,31,120,30,179,31,193,31,183,31,183,30,191,31,23,31,14,31,111,31,171,31,171,30,171,29,44,31,118,31,118,30,126,31,153,31,237,31,237,30,237,31,29,31,116,31,125,31,235,31,201,31,133,31,11,31,12,31,77,31,77,30,62,31,201,31,201,30,201,29,200,31,40,31,197,31,117,31,150,31,203,31,23,31,82,31,119,31,56,31,105,31,105,30,165,31,124,31,124,30,124,29,176,31,176,30,90,31,40,31,192,31,192,30,58,31,58,30,219,31,24,31,24,30,33,31,219,31,233,31,217,31,67,31,67,30,166,31,217,31,39,31,34,31,11,31,74,31,161,31,173,31,39,31,159,31,233,31,142,31,82,31,82,30,204,31,28,31,98,31,234,31,249,31,29,31,29,30,35,31,35,30,198,31,212,31,212,30,236,31,42,31,204,31,186,31,84,31,173,31,96,31,96,30,143,31,100,31,207,31,83,31,113,31,31,31,31,30,31,29,188,31,234,31,82,31,2,31,22,31,133,31,133,30,133,29,111,31,250,31,1,31,149,31,130,31,159,31,197,31,102,31,102,30,182,31,227,31,169,31,224,31,128,31,69,31,100,31,31,31,136,31,28,31,142,31,159,31,159,30,159,29,159,28,131,31,241,31,169,31,111,31,209,31,75,31,39,31,240,31,240,30,12,31,12,30,12,29,18,31,55,31,66,31,66,30,81,31,13,31,7,31,42,31,52,31,8,31,212,31,91,31,111,31,3,31,44,31,176,31,133,31,70,31,70,30,105,31,138,31,64,31,61,31,25,31,108,31,247,31,148,31,148,30,143,31,104,31,196,31,129,31,106,31,106,30,119,31,119,30,46,31,174,31,24,31,24,30,59,31,255,31,6,31,89,31,6,31,6,30,93,31,122,31,122,30,122,29,218,31,152,31,22,31,125,31,145,31,61,31,72,31,112,31,175,31,189,31,189,30,198,31,193,31,156,31,156,30,248,31,15,31,15,30,15,29,15,28,240,31,173,31,31,31,1,31,1,30,1,29,50,31,48,31,48,30,137,31,39,31,234,31,23,31,195,31,195,30,195,29,41,31,191,31,192,31,30,31,30,30,239,31,111,31,171,31,171,30,43,31,43,30,35,31,217,31,124,31,96,31,23,31,135,31,194,31,194,30,48,31,48,30,233,31,205,31,205,30,205,29,116,31,229,31,229,30,228,31,228,31,244,31,125,31,156,31,249,31,53,31,58,31,58,30,70,31,138,31,185,31,235,31,173,31,166,31,143,31,94,31,250,31,199,31,53,31,141,31,235,31,64,31,64,30,22,31,22,30,69,31,69,30,168,31,113,31,79,31,195,31,229,31,68,31,255,31,255,30,255,29,60,31,228,31,143,31,143,30,22,31,150,31,139,31,154,31,1,31,125,31,84,31,84,30,143,31,143,30,199,31,86,31,56,31,56,30,137,31,221,31,126,31,67,31,227,31,190,31,249,31,188,31,80,31,171,31,45,31,47,31,180,31,191,31,102,31,162,31,162,30,159,31,101,31,71,31,71,30,229,31,54,31,43,31,43,30,200,31,200,30,200,29,159,31,106,31,39,31,169,31,86,31,86,30,53,31,149,31,90,31,147,31,111,31,200,31,93,31,93,30,48,31,110,31,152,31,13,31,83,31,186,31,186,30,255,31,171,31,101,31,97,31,12,31,12,30,185,31,185,30,185,29,26,31,26,30,225,31,177,31,203,31,141,31,141,30,69,31,2,31,2,30,147,31,19,31,19,30,39,31,217,31,67,31,59,31,59,30,197,31,207,31,234,31,71,31,60,31,17,31,152,31,67,31,211,31,161,31,211,31,21,31,76,31,205,31,205,30,192,31,192,30,66,31,171,31,197,31,196,31,120,31,159,31,34,31,161,31,240,31,104,31,26,31,13,31,161,31,161,30,80,31,80,30,169,31,109,31,182,31,216,31,109,31,192,31,132,31,249,31,4,31,4,30,227,31,227,30,15,31,162,31,48,31,232,31,236,31,236,30,179,31,111,31,46,31,199,31,7,31,171,31,219,31,198,31,91,31,72,31,103,31,239,31,246,31,117,31,140,31,140,30,101,31,101,30,35,31,71,31,185,31,118,31,121,31,195,31,237,31,104,31,165,31,241,31,65,31,44,31,75,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
