-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_137 is
end project_tb_137;

architecture project_tb_arch_137 of project_tb_137 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 1023;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (70,0,252,0,237,0,73,0,238,0,28,0,222,0,130,0,0,0,0,0,0,0,76,0,72,0,203,0,104,0,3,0,18,0,0,0,181,0,232,0,227,0,0,0,239,0,5,0,0,0,254,0,204,0,116,0,186,0,56,0,129,0,88,0,0,0,0,0,42,0,0,0,155,0,0,0,9,0,60,0,224,0,3,0,0,0,132,0,24,0,227,0,107,0,27,0,105,0,44,0,16,0,114,0,126,0,181,0,80,0,29,0,93,0,0,0,0,0,185,0,42,0,168,0,41,0,98,0,0,0,137,0,194,0,91,0,185,0,71,0,179,0,205,0,135,0,177,0,223,0,16,0,148,0,159,0,193,0,0,0,79,0,0,0,222,0,157,0,0,0,216,0,136,0,209,0,0,0,232,0,42,0,74,0,116,0,231,0,0,0,0,0,9,0,245,0,209,0,0,0,218,0,0,0,6,0,184,0,175,0,227,0,76,0,48,0,41,0,18,0,93,0,0,0,17,0,110,0,6,0,0,0,214,0,105,0,245,0,20,0,0,0,176,0,0,0,59,0,0,0,228,0,247,0,63,0,138,0,77,0,156,0,0,0,34,0,74,0,19,0,97,0,212,0,246,0,105,0,6,0,237,0,193,0,100,0,0,0,124,0,135,0,107,0,174,0,118,0,231,0,166,0,0,0,236,0,205,0,105,0,128,0,92,0,185,0,0,0,0,0,198,0,115,0,167,0,71,0,218,0,0,0,153,0,138,0,37,0,32,0,29,0,0,0,28,0,58,0,142,0,0,0,92,0,110,0,245,0,34,0,240,0,0,0,185,0,132,0,90,0,212,0,81,0,243,0,166,0,0,0,220,0,195,0,67,0,157,0,83,0,91,0,116,0,0,0,0,0,115,0,0,0,219,0,160,0,166,0,5,0,0,0,0,0,178,0,72,0,255,0,154,0,192,0,154,0,140,0,197,0,183,0,0,0,218,0,56,0,38,0,227,0,195,0,214,0,141,0,254,0,68,0,0,0,40,0,0,0,0,0,85,0,0,0,35,0,149,0,77,0,210,0,21,0,175,0,159,0,0,0,206,0,125,0,216,0,228,0,252,0,0,0,144,0,43,0,60,0,186,0,143,0,0,0,0,0,0,0,163,0,54,0,22,0,140,0,74,0,58,0,132,0,56,0,0,0,131,0,231,0,168,0,242,0,0,0,61,0,251,0,7,0,12,0,96,0,213,0,0,0,79,0,150,0,33,0,99,0,192,0,0,0,128,0,0,0,140,0,30,0,0,0,99,0,0,0,0,0,42,0,0,0,123,0,131,0,0,0,77,0,144,0,51,0,0,0,0,0,67,0,238,0,0,0,217,0,100,0,67,0,74,0,158,0,101,0,128,0,49,0,49,0,0,0,28,0,125,0,224,0,109,0,180,0,0,0,0,0,199,0,132,0,28,0,59,0,31,0,84,0,127,0,14,0,199,0,0,0,234,0,223,0,239,0,0,0,25,0,178,0,90,0,171,0,204,0,82,0,165,0,212,0,0,0,72,0,0,0,0,0,82,0,61,0,0,0,4,0,176,0,163,0,39,0,210,0,90,0,114,0,4,0,77,0,123,0,83,0,100,0,238,0,44,0,45,0,0,0,120,0,170,0,14,0,171,0,0,0,70,0,219,0,41,0,234,0,183,0,243,0,58,0,199,0,0,0,182,0,0,0,140,0,188,0,238,0,197,0,11,0,254,0,0,0,230,0,33,0,0,0,206,0,0,0,44,0,0,0,191,0,137,0,0,0,93,0,83,0,0,0,43,0,0,0,181,0,107,0,129,0,0,0,0,0,109,0,7,0,6,0,171,0,252,0,50,0,61,0,172,0,251,0,64,0,103,0,136,0,0,0,179,0,4,0,104,0,0,0,91,0,0,0,56,0,190,0,220,0,1,0,83,0,184,0,0,0,104,0,75,0,150,0,49,0,43,0,157,0,51,0,158,0,39,0,157,0,196,0,91,0,49,0,107,0,96,0,161,0,219,0,209,0,15,0,60,0,60,0,113,0,242,0,249,0,0,0,0,0,11,0,0,0,0,0,31,0,180,0,47,0,156,0,49,0,110,0,23,0,196,0,20,0,178,0,51,0,96,0,22,0,156,0,227,0,0,0,252,0,220,0,69,0,0,0,0,0,18,0,214,0,77,0,0,0,44,0,0,0,110,0,103,0,154,0,144,0,129,0,3,0,0,0,232,0,76,0,244,0,12,0,243,0,69,0,35,0,0,0,5,0,139,0,0,0,1,0,0,0,69,0,19,0,131,0,148,0,80,0,109,0,185,0,232,0,170,0,155,0,167,0,13,0,111,0,255,0,39,0,28,0,187,0,191,0,0,0,134,0,138,0,0,0,0,0,174,0,34,0,0,0,0,0,169,0,96,0,0,0,24,0,115,0,65,0,219,0,55,0,195,0,16,0,87,0,176,0,17,0,35,0,0,0,158,0,230,0,39,0,232,0,31,0,252,0,83,0,0,0,69,0,0,0,98,0,11,0,0,0,147,0,0,0,249,0,165,0,0,0,126,0,246,0,93,0,0,0,122,0,134,0,28,0,140,0,235,0,69,0,97,0,248,0,183,0,204,0,51,0,0,0,0,0,237,0,200,0,124,0,100,0,181,0,0,0,170,0,0,0,0,0,177,0,13,0,243,0,170,0,127,0,25,0,159,0,174,0,255,0,27,0,58,0,114,0,86,0,160,0,168,0,94,0,41,0,230,0,102,0,66,0,0,0,8,0,0,0,0,0,217,0,107,0,211,0,0,0,221,0,216,0,194,0,35,0,27,0,0,0,200,0,0,0,48,0,176,0,72,0,255,0,170,0,0,0,40,0,208,0,81,0,3,0,204,0,226,0,217,0,98,0,197,0,0,0,188,0,204,0,192,0,148,0,186,0,0,0,0,0,131,0,239,0,0,0,208,0,0,0,29,0,116,0,0,0,192,0,47,0,160,0,0,0,222,0,83,0,0,0,21,0,54,0,132,0,244,0,93,0,91,0,178,0,214,0,191,0,0,0,226,0,103,0,22,0,43,0,69,0,144,0,228,0,68,0,31,0,83,0,214,0,193,0,202,0,0,0,250,0,75,0,233,0,55,0,212,0,0,0,147,0,14,0,93,0,249,0,141,0,255,0,112,0,66,0,56,0,225,0,155,0,98,0,127,0,149,0,78,0,15,0,138,0,0,0,219,0,12,0,83,0,0,0,5,0,0,0,249,0,203,0,216,0,177,0,103,0,95,0,0,0,76,0,125,0,190,0,211,0,3,0,208,0,0,0,61,0,158,0,122,0,5,0,39,0,34,0,0,0,194,0,149,0,96,0,0,0,6,0,115,0,201,0,61,0,254,0,87,0,187,0,0,0,88,0,175,0,0,0,250,0,135,0,0,0,160,0,197,0,113,0,79,0,187,0,0,0,234,0,0,0,71,0,230,0,249,0,151,0,0,0,77,0,194,0,53,0,24,0,0,0,43,0,240,0,162,0,234,0,3,0,37,0,38,0,0,0,198,0,145,0,4,0,184,0,234,0,224,0,158,0,222,0,193,0,185,0,235,0,112,0,0,0,232,0,111,0,28,0,0,0,91,0,106,0,59,0,105,0,9,0,141,0,78,0,17,0,118,0,0,0,0,0,147,0,249,0,235,0,159,0,253,0,37,0,0,0,92,0,80,0,0,0,0,0,0,0,0,0,247,0,53,0,44,0,34,0,34,0,216,0,83,0,50,0,118,0,211,0,46,0,0,0,70,0,66,0,56,0,185,0,3,0,66,0,0,0,67,0,118,0,98,0,206,0,208,0,0,0,0,0,239,0,243,0,243,0,124,0,137,0,35,0,55,0,41,0,80,0,87,0,167,0,163,0,20,0,132,0,82,0,180,0,170,0,200,0,0,0,103,0,162,0,191,0,0,0,248,0,211,0,247,0,250,0,252,0,203,0,35,0,145,0,0,0,0,0,243,0,0,0,150,0,231,0,0,0,154,0,94,0,0,0,164,0,90,0,167,0,197,0,206,0,0,0,0,0,197,0,58,0,3,0,33,0,125,0,15,0,121,0,147,0,159,0,100,0,172,0,137,0,77,0,10,0,44,0,96,0,229,0,188,0,200,0,14,0,244,0,0,0,23,0,117,0,8,0,93,0,13,0,140,0,135,0,91,0,65,0,8,0,71,0,194,0,0,0,0,0,113,0,22,0,251,0,0,0,2,0,0,0,143,0,42,0,97,0,213,0,174,0,98,0,180,0,97,0,209,0,221,0,135,0,221,0,179,0,115,0,160,0,48,0,152,0,0,0,85,0,60,0,112,0,0,0,118,0,162,0,0,0,0,0,0,0,47,0,63,0,23,0,254,0,202,0,103,0,174,0,227,0,114,0,53,0,110,0,198,0,73,0,91,0,0,0,0,0,0,0,94,0,157,0,82,0,8,0,253,0,200,0,209,0,159,0,200,0,121,0,230,0,0,0,0,0,130,0,0,0,26,0,18,0,143,0,87,0,65,0,126,0,169,0,1,0,124,0,0,0,133,0,126,0,54,0,0,0,250,0,0,0,41,0,91,0,0,0);
signal scenario_full  : scenario_type := (70,31,252,31,237,31,73,31,238,31,28,31,222,31,130,31,130,30,130,29,130,28,76,31,72,31,203,31,104,31,3,31,18,31,18,30,181,31,232,31,227,31,227,30,239,31,5,31,5,30,254,31,204,31,116,31,186,31,56,31,129,31,88,31,88,30,88,29,42,31,42,30,155,31,155,30,9,31,60,31,224,31,3,31,3,30,132,31,24,31,227,31,107,31,27,31,105,31,44,31,16,31,114,31,126,31,181,31,80,31,29,31,93,31,93,30,93,29,185,31,42,31,168,31,41,31,98,31,98,30,137,31,194,31,91,31,185,31,71,31,179,31,205,31,135,31,177,31,223,31,16,31,148,31,159,31,193,31,193,30,79,31,79,30,222,31,157,31,157,30,216,31,136,31,209,31,209,30,232,31,42,31,74,31,116,31,231,31,231,30,231,29,9,31,245,31,209,31,209,30,218,31,218,30,6,31,184,31,175,31,227,31,76,31,48,31,41,31,18,31,93,31,93,30,17,31,110,31,6,31,6,30,214,31,105,31,245,31,20,31,20,30,176,31,176,30,59,31,59,30,228,31,247,31,63,31,138,31,77,31,156,31,156,30,34,31,74,31,19,31,97,31,212,31,246,31,105,31,6,31,237,31,193,31,100,31,100,30,124,31,135,31,107,31,174,31,118,31,231,31,166,31,166,30,236,31,205,31,105,31,128,31,92,31,185,31,185,30,185,29,198,31,115,31,167,31,71,31,218,31,218,30,153,31,138,31,37,31,32,31,29,31,29,30,28,31,58,31,142,31,142,30,92,31,110,31,245,31,34,31,240,31,240,30,185,31,132,31,90,31,212,31,81,31,243,31,166,31,166,30,220,31,195,31,67,31,157,31,83,31,91,31,116,31,116,30,116,29,115,31,115,30,219,31,160,31,166,31,5,31,5,30,5,29,178,31,72,31,255,31,154,31,192,31,154,31,140,31,197,31,183,31,183,30,218,31,56,31,38,31,227,31,195,31,214,31,141,31,254,31,68,31,68,30,40,31,40,30,40,29,85,31,85,30,35,31,149,31,77,31,210,31,21,31,175,31,159,31,159,30,206,31,125,31,216,31,228,31,252,31,252,30,144,31,43,31,60,31,186,31,143,31,143,30,143,29,143,28,163,31,54,31,22,31,140,31,74,31,58,31,132,31,56,31,56,30,131,31,231,31,168,31,242,31,242,30,61,31,251,31,7,31,12,31,96,31,213,31,213,30,79,31,150,31,33,31,99,31,192,31,192,30,128,31,128,30,140,31,30,31,30,30,99,31,99,30,99,29,42,31,42,30,123,31,131,31,131,30,77,31,144,31,51,31,51,30,51,29,67,31,238,31,238,30,217,31,100,31,67,31,74,31,158,31,101,31,128,31,49,31,49,31,49,30,28,31,125,31,224,31,109,31,180,31,180,30,180,29,199,31,132,31,28,31,59,31,31,31,84,31,127,31,14,31,199,31,199,30,234,31,223,31,239,31,239,30,25,31,178,31,90,31,171,31,204,31,82,31,165,31,212,31,212,30,72,31,72,30,72,29,82,31,61,31,61,30,4,31,176,31,163,31,39,31,210,31,90,31,114,31,4,31,77,31,123,31,83,31,100,31,238,31,44,31,45,31,45,30,120,31,170,31,14,31,171,31,171,30,70,31,219,31,41,31,234,31,183,31,243,31,58,31,199,31,199,30,182,31,182,30,140,31,188,31,238,31,197,31,11,31,254,31,254,30,230,31,33,31,33,30,206,31,206,30,44,31,44,30,191,31,137,31,137,30,93,31,83,31,83,30,43,31,43,30,181,31,107,31,129,31,129,30,129,29,109,31,7,31,6,31,171,31,252,31,50,31,61,31,172,31,251,31,64,31,103,31,136,31,136,30,179,31,4,31,104,31,104,30,91,31,91,30,56,31,190,31,220,31,1,31,83,31,184,31,184,30,104,31,75,31,150,31,49,31,43,31,157,31,51,31,158,31,39,31,157,31,196,31,91,31,49,31,107,31,96,31,161,31,219,31,209,31,15,31,60,31,60,31,113,31,242,31,249,31,249,30,249,29,11,31,11,30,11,29,31,31,180,31,47,31,156,31,49,31,110,31,23,31,196,31,20,31,178,31,51,31,96,31,22,31,156,31,227,31,227,30,252,31,220,31,69,31,69,30,69,29,18,31,214,31,77,31,77,30,44,31,44,30,110,31,103,31,154,31,144,31,129,31,3,31,3,30,232,31,76,31,244,31,12,31,243,31,69,31,35,31,35,30,5,31,139,31,139,30,1,31,1,30,69,31,19,31,131,31,148,31,80,31,109,31,185,31,232,31,170,31,155,31,167,31,13,31,111,31,255,31,39,31,28,31,187,31,191,31,191,30,134,31,138,31,138,30,138,29,174,31,34,31,34,30,34,29,169,31,96,31,96,30,24,31,115,31,65,31,219,31,55,31,195,31,16,31,87,31,176,31,17,31,35,31,35,30,158,31,230,31,39,31,232,31,31,31,252,31,83,31,83,30,69,31,69,30,98,31,11,31,11,30,147,31,147,30,249,31,165,31,165,30,126,31,246,31,93,31,93,30,122,31,134,31,28,31,140,31,235,31,69,31,97,31,248,31,183,31,204,31,51,31,51,30,51,29,237,31,200,31,124,31,100,31,181,31,181,30,170,31,170,30,170,29,177,31,13,31,243,31,170,31,127,31,25,31,159,31,174,31,255,31,27,31,58,31,114,31,86,31,160,31,168,31,94,31,41,31,230,31,102,31,66,31,66,30,8,31,8,30,8,29,217,31,107,31,211,31,211,30,221,31,216,31,194,31,35,31,27,31,27,30,200,31,200,30,48,31,176,31,72,31,255,31,170,31,170,30,40,31,208,31,81,31,3,31,204,31,226,31,217,31,98,31,197,31,197,30,188,31,204,31,192,31,148,31,186,31,186,30,186,29,131,31,239,31,239,30,208,31,208,30,29,31,116,31,116,30,192,31,47,31,160,31,160,30,222,31,83,31,83,30,21,31,54,31,132,31,244,31,93,31,91,31,178,31,214,31,191,31,191,30,226,31,103,31,22,31,43,31,69,31,144,31,228,31,68,31,31,31,83,31,214,31,193,31,202,31,202,30,250,31,75,31,233,31,55,31,212,31,212,30,147,31,14,31,93,31,249,31,141,31,255,31,112,31,66,31,56,31,225,31,155,31,98,31,127,31,149,31,78,31,15,31,138,31,138,30,219,31,12,31,83,31,83,30,5,31,5,30,249,31,203,31,216,31,177,31,103,31,95,31,95,30,76,31,125,31,190,31,211,31,3,31,208,31,208,30,61,31,158,31,122,31,5,31,39,31,34,31,34,30,194,31,149,31,96,31,96,30,6,31,115,31,201,31,61,31,254,31,87,31,187,31,187,30,88,31,175,31,175,30,250,31,135,31,135,30,160,31,197,31,113,31,79,31,187,31,187,30,234,31,234,30,71,31,230,31,249,31,151,31,151,30,77,31,194,31,53,31,24,31,24,30,43,31,240,31,162,31,234,31,3,31,37,31,38,31,38,30,198,31,145,31,4,31,184,31,234,31,224,31,158,31,222,31,193,31,185,31,235,31,112,31,112,30,232,31,111,31,28,31,28,30,91,31,106,31,59,31,105,31,9,31,141,31,78,31,17,31,118,31,118,30,118,29,147,31,249,31,235,31,159,31,253,31,37,31,37,30,92,31,80,31,80,30,80,29,80,28,80,27,247,31,53,31,44,31,34,31,34,31,216,31,83,31,50,31,118,31,211,31,46,31,46,30,70,31,66,31,56,31,185,31,3,31,66,31,66,30,67,31,118,31,98,31,206,31,208,31,208,30,208,29,239,31,243,31,243,31,124,31,137,31,35,31,55,31,41,31,80,31,87,31,167,31,163,31,20,31,132,31,82,31,180,31,170,31,200,31,200,30,103,31,162,31,191,31,191,30,248,31,211,31,247,31,250,31,252,31,203,31,35,31,145,31,145,30,145,29,243,31,243,30,150,31,231,31,231,30,154,31,94,31,94,30,164,31,90,31,167,31,197,31,206,31,206,30,206,29,197,31,58,31,3,31,33,31,125,31,15,31,121,31,147,31,159,31,100,31,172,31,137,31,77,31,10,31,44,31,96,31,229,31,188,31,200,31,14,31,244,31,244,30,23,31,117,31,8,31,93,31,13,31,140,31,135,31,91,31,65,31,8,31,71,31,194,31,194,30,194,29,113,31,22,31,251,31,251,30,2,31,2,30,143,31,42,31,97,31,213,31,174,31,98,31,180,31,97,31,209,31,221,31,135,31,221,31,179,31,115,31,160,31,48,31,152,31,152,30,85,31,60,31,112,31,112,30,118,31,162,31,162,30,162,29,162,28,47,31,63,31,23,31,254,31,202,31,103,31,174,31,227,31,114,31,53,31,110,31,198,31,73,31,91,31,91,30,91,29,91,28,94,31,157,31,82,31,8,31,253,31,200,31,209,31,159,31,200,31,121,31,230,31,230,30,230,29,130,31,130,30,26,31,18,31,143,31,87,31,65,31,126,31,169,31,1,31,124,31,124,30,133,31,126,31,54,31,54,30,250,31,250,30,41,31,91,31,91,30);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
