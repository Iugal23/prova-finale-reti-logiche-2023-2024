-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb is
end project_tb;

architecture project_tb_arch of project_tb is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 221;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (244,0,0,0,0,0,25,0,6,0,132,0,0,0,0,0,156,0,211,0,6,0,184,0,58,0,251,0,70,0,7,0,0,0,161,0,138,0,0,0,193,0,148,0,205,0,0,0,98,0,159,0,157,0,0,0,0,0,204,0,24,0,0,0,197,0,223,0,101,0,58,0,178,0,204,0,0,0,105,0,139,0,109,0,207,0,97,0,219,0,115,0,192,0,0,0,86,0,17,0,131,0,150,0,133,0,0,0,205,0,172,0,212,0,0,0,93,0,31,0,0,0,0,0,0,0,0,0,146,0,152,0,77,0,81,0,78,0,0,0,78,0,180,0,51,0,24,0,194,0,7,0,147,0,0,0,189,0,231,0,163,0,76,0,143,0,100,0,67,0,41,0,84,0,60,0,255,0,44,0,134,0,28,0,33,0,149,0,0,0,247,0,134,0,69,0,163,0,141,0,207,0,204,0,186,0,168,0,215,0,0,0,226,0,39,0,0,0,255,0,153,0,136,0,249,0,0,0,0,0,5,0,98,0,173,0,96,0,161,0,136,0,0,0,162,0,248,0,117,0,149,0,87,0,0,0,0,0,43,0,67,0,28,0,0,0,42,0,115,0,201,0,253,0,238,0,143,0,0,0,190,0,0,0,35,0,111,0,25,0,172,0,61,0,127,0,13,0,173,0,3,0,0,0,91,0,0,0,236,0,0,0,217,0,0,0,25,0,131,0,190,0,111,0,239,0,170,0,45,0,160,0,100,0,89,0,0,0,101,0,194,0,122,0,11,0,0,0,158,0,0,0,206,0,0,0,104,0,0,0,76,0,133,0,48,0,155,0,235,0,45,0,192,0,82,0,0,0,0,0,35,0,21,0,142,0,221,0,0,0,0,0,160,0,165,0,127,0,168,0,175,0,156,0,25,0,223,0,104,0,0,0,13,0,166,0,113,0,0,0,54,0,164,0,0,0,174,0,0,0,49,0,12,0,63,0,120,0,92,0,222,0);
signal scenario_full  : scenario_type := (244,31,244,30,244,29,25,31,6,31,132,31,132,30,132,29,156,31,211,31,6,31,184,31,58,31,251,31,70,31,7,31,7,30,161,31,138,31,138,30,193,31,148,31,205,31,205,30,98,31,159,31,157,31,157,30,157,29,204,31,24,31,24,30,197,31,223,31,101,31,58,31,178,31,204,31,204,30,105,31,139,31,109,31,207,31,97,31,219,31,115,31,192,31,192,30,86,31,17,31,131,31,150,31,133,31,133,30,205,31,172,31,212,31,212,30,93,31,31,31,31,30,31,29,31,28,31,27,146,31,152,31,77,31,81,31,78,31,78,30,78,31,180,31,51,31,24,31,194,31,7,31,147,31,147,30,189,31,231,31,163,31,76,31,143,31,100,31,67,31,41,31,84,31,60,31,255,31,44,31,134,31,28,31,33,31,149,31,149,30,247,31,134,31,69,31,163,31,141,31,207,31,204,31,186,31,168,31,215,31,215,30,226,31,39,31,39,30,255,31,153,31,136,31,249,31,249,30,249,29,5,31,98,31,173,31,96,31,161,31,136,31,136,30,162,31,248,31,117,31,149,31,87,31,87,30,87,29,43,31,67,31,28,31,28,30,42,31,115,31,201,31,253,31,238,31,143,31,143,30,190,31,190,30,35,31,111,31,25,31,172,31,61,31,127,31,13,31,173,31,3,31,3,30,91,31,91,30,236,31,236,30,217,31,217,30,25,31,131,31,190,31,111,31,239,31,170,31,45,31,160,31,100,31,89,31,89,30,101,31,194,31,122,31,11,31,11,30,158,31,158,30,206,31,206,30,104,31,104,30,76,31,133,31,48,31,155,31,235,31,45,31,192,31,82,31,82,30,82,29,35,31,21,31,142,31,221,31,221,30,221,29,160,31,165,31,127,31,168,31,175,31,156,31,25,31,223,31,104,31,104,30,13,31,166,31,113,31,113,30,54,31,164,31,164,30,174,31,174,30,49,31,12,31,63,31,120,31,92,31,222,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
