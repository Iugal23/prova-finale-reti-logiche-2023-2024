-- TB EXAMPLE PFRL 2023-2024

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;

entity project_tb_911 is
end project_tb_911;

architecture project_tb_arch_911 of project_tb_911 is
    constant CLOCK_PERIOD : time := 20 ns;
    signal tb_clk : std_logic := '0';
    signal tb_rst, tb_start, tb_done : std_logic;
    signal tb_add : std_logic_vector(15 downto 0);
    signal tb_k   : std_logic_vector(9 downto 0);

    signal tb_o_mem_addr, exc_o_mem_addr, init_o_mem_addr : std_logic_vector(15 downto 0);
    signal tb_o_mem_data, exc_o_mem_data, init_o_mem_data : std_logic_vector(7 downto 0);
    signal tb_i_mem_data : std_logic_vector(7 downto 0);
    signal tb_o_mem_we, tb_o_mem_en, exc_o_mem_we, exc_o_mem_en, init_o_mem_we, init_o_mem_en : std_logic;

    type ram_type is array (65535 downto 0) of std_logic_vector(7 downto 0);
    signal RAM : ram_type := (OTHERS => "00000000");

constant SCENARIO_LENGTH : integer := 745;
    type scenario_type is array (0 to SCENARIO_LENGTH*2-1) of integer;

signal scenario_input : scenario_type := (69,0,95,0,99,0,58,0,2,0,89,0,90,0,86,0,48,0,92,0,117,0,0,0,98,0,0,0,170,0,0,0,104,0,141,0,0,0,244,0,15,0,15,0,54,0,130,0,131,0,100,0,113,0,161,0,254,0,179,0,0,0,224,0,0,0,161,0,0,0,195,0,61,0,85,0,70,0,54,0,170,0,0,0,0,0,109,0,141,0,0,0,0,0,64,0,147,0,21,0,9,0,211,0,207,0,118,0,140,0,177,0,139,0,0,0,0,0,43,0,73,0,159,0,197,0,0,0,43,0,0,0,89,0,207,0,8,0,234,0,134,0,107,0,112,0,0,0,106,0,255,0,176,0,233,0,0,0,2,0,125,0,156,0,210,0,86,0,132,0,212,0,129,0,64,0,0,0,0,0,0,0,146,0,14,0,104,0,216,0,25,0,82,0,159,0,221,0,0,0,124,0,97,0,102,0,148,0,58,0,54,0,108,0,155,0,23,0,19,0,17,0,0,0,106,0,67,0,247,0,0,0,174,0,105,0,234,0,0,0,116,0,212,0,19,0,0,0,223,0,48,0,30,0,217,0,168,0,242,0,49,0,0,0,139,0,0,0,184,0,200,0,199,0,117,0,199,0,39,0,189,0,191,0,19,0,111,0,166,0,147,0,22,0,0,0,41,0,250,0,221,0,0,0,126,0,0,0,0,0,93,0,121,0,115,0,138,0,47,0,204,0,0,0,63,0,0,0,252,0,0,0,0,0,208,0,0,0,252,0,72,0,0,0,0,0,0,0,165,0,154,0,176,0,87,0,215,0,222,0,120,0,6,0,102,0,0,0,222,0,0,0,0,0,0,0,60,0,111,0,90,0,204,0,187,0,43,0,71,0,172,0,208,0,95,0,202,0,77,0,108,0,137,0,105,0,11,0,0,0,53,0,60,0,76,0,129,0,246,0,0,0,65,0,24,0,55,0,0,0,0,0,0,0,95,0,0,0,97,0,211,0,218,0,237,0,0,0,223,0,26,0,81,0,55,0,68,0,207,0,32,0,30,0,60,0,0,0,3,0,22,0,11,0,87,0,141,0,49,0,0,0,239,0,6,0,0,0,0,0,92,0,89,0,132,0,187,0,112,0,100,0,82,0,202,0,136,0,91,0,122,0,242,0,231,0,145,0,227,0,40,0,17,0,136,0,166,0,235,0,41,0,187,0,2,0,182,0,47,0,87,0,0,0,55,0,238,0,0,0,213,0,0,0,218,0,132,0,162,0,102,0,3,0,127,0,27,0,24,0,67,0,218,0,193,0,0,0,113,0,142,0,31,0,159,0,32,0,0,0,229,0,89,0,0,0,0,0,53,0,64,0,83,0,143,0,45,0,58,0,229,0,100,0,95,0,78,0,182,0,165,0,0,0,0,0,241,0,15,0,0,0,0,0,29,0,80,0,36,0,38,0,120,0,77,0,0,0,226,0,0,0,192,0,121,0,233,0,208,0,190,0,0,0,0,0,10,0,72,0,193,0,0,0,129,0,0,0,50,0,199,0,183,0,72,0,139,0,0,0,240,0,117,0,228,0,133,0,194,0,42,0,252,0,116,0,203,0,0,0,199,0,196,0,58,0,184,0,178,0,94,0,9,0,43,0,21,0,0,0,156,0,2,0,0,0,159,0,226,0,0,0,211,0,11,0,90,0,122,0,120,0,14,0,188,0,225,0,235,0,0,0,10,0,38,0,201,0,0,0,118,0,0,0,0,0,143,0,0,0,18,0,250,0,184,0,3,0,16,0,80,0,230,0,212,0,242,0,188,0,0,0,0,0,54,0,193,0,18,0,32,0,114,0,191,0,169,0,0,0,68,0,81,0,0,0,200,0,48,0,98,0,0,0,99,0,2,0,190,0,106,0,0,0,60,0,0,0,27,0,10,0,79,0,207,0,186,0,0,0,86,0,0,0,33,0,18,0,76,0,162,0,1,0,157,0,233,0,221,0,112,0,0,0,174,0,0,0,185,0,23,0,72,0,0,0,193,0,178,0,99,0,229,0,0,0,0,0,185,0,101,0,177,0,0,0,131,0,0,0,255,0,186,0,213,0,189,0,0,0,79,0,172,0,125,0,75,0,116,0,218,0,228,0,0,0,116,0,170,0,50,0,32,0,225,0,0,0,225,0,102,0,68,0,143,0,250,0,224,0,163,0,118,0,11,0,251,0,0,0,0,0,210,0,0,0,73,0,246,0,45,0,61,0,221,0,33,0,227,0,72,0,149,0,217,0,38,0,0,0,65,0,176,0,161,0,17,0,200,0,85,0,0,0,0,0,95,0,0,0,0,0,224,0,0,0,180,0,225,0,69,0,190,0,78,0,186,0,111,0,171,0,25,0,98,0,192,0,0,0,164,0,0,0,121,0,136,0,201,0,19,0,226,0,123,0,0,0,116,0,0,0,243,0,139,0,165,0,0,0,92,0,241,0,56,0,119,0,170,0,184,0,120,0,79,0,0,0,0,0,49,0,62,0,77,0,0,0,5,0,130,0,0,0,0,0,0,0,11,0,237,0,0,0,0,0,90,0,30,0,148,0,247,0,32,0,79,0,116,0,0,0,137,0,15,0,120,0,0,0,189,0,108,0,87,0,75,0,254,0,0,0,40,0,212,0,0,0,159,0,7,0,70,0,208,0,198,0,5,0,169,0,139,0,59,0,203,0,93,0,173,0,101,0,21,0,0,0,0,0,209,0,226,0,0,0,79,0,183,0,168,0,227,0,231,0,112,0,1,0,45,0,222,0,160,0,238,0,157,0,71,0,210,0,16,0,112,0,213,0,75,0,216,0,128,0,254,0,138,0,241,0,204,0,229,0,156,0,234,0,54,0,0,0,26,0,112,0,233,0,0,0,157,0,168,0,149,0,0,0,246,0,41,0,165,0,196,0,184,0,238,0,202,0,127,0,219,0,96,0,86,0,50,0,138,0,253,0,237,0,220,0,34,0,87,0,44,0,58,0,0,0,41,0,126,0,255,0,98,0,147,0,116,0,206,0,90,0,114,0,40,0,242,0,76,0,205,0,0,0,205,0,0,0,0,0,0,0,192,0,55,0,132,0,91,0,120,0,72,0,77,0,46,0,215,0,92,0,37,0,22,0,133,0,126,0,109,0,9,0,39,0,238,0,29,0,179,0,64,0,188,0,0,0,3,0,135,0,141,0,209,0,0,0,139,0,87,0,0,0,75,0,0,0,246,0,0,0,0,0,0,0,208,0,230,0,23,0,65,0,0,0,62,0,153,0,95,0,48,0,0,0,119,0,156,0,252,0,0,0,215,0,222,0,166,0,52,0,95,0,241,0,143,0,0,0,0,0,107,0);
signal scenario_full  : scenario_type := (69,31,95,31,99,31,58,31,2,31,89,31,90,31,86,31,48,31,92,31,117,31,117,30,98,31,98,30,170,31,170,30,104,31,141,31,141,30,244,31,15,31,15,31,54,31,130,31,131,31,100,31,113,31,161,31,254,31,179,31,179,30,224,31,224,30,161,31,161,30,195,31,61,31,85,31,70,31,54,31,170,31,170,30,170,29,109,31,141,31,141,30,141,29,64,31,147,31,21,31,9,31,211,31,207,31,118,31,140,31,177,31,139,31,139,30,139,29,43,31,73,31,159,31,197,31,197,30,43,31,43,30,89,31,207,31,8,31,234,31,134,31,107,31,112,31,112,30,106,31,255,31,176,31,233,31,233,30,2,31,125,31,156,31,210,31,86,31,132,31,212,31,129,31,64,31,64,30,64,29,64,28,146,31,14,31,104,31,216,31,25,31,82,31,159,31,221,31,221,30,124,31,97,31,102,31,148,31,58,31,54,31,108,31,155,31,23,31,19,31,17,31,17,30,106,31,67,31,247,31,247,30,174,31,105,31,234,31,234,30,116,31,212,31,19,31,19,30,223,31,48,31,30,31,217,31,168,31,242,31,49,31,49,30,139,31,139,30,184,31,200,31,199,31,117,31,199,31,39,31,189,31,191,31,19,31,111,31,166,31,147,31,22,31,22,30,41,31,250,31,221,31,221,30,126,31,126,30,126,29,93,31,121,31,115,31,138,31,47,31,204,31,204,30,63,31,63,30,252,31,252,30,252,29,208,31,208,30,252,31,72,31,72,30,72,29,72,28,165,31,154,31,176,31,87,31,215,31,222,31,120,31,6,31,102,31,102,30,222,31,222,30,222,29,222,28,60,31,111,31,90,31,204,31,187,31,43,31,71,31,172,31,208,31,95,31,202,31,77,31,108,31,137,31,105,31,11,31,11,30,53,31,60,31,76,31,129,31,246,31,246,30,65,31,24,31,55,31,55,30,55,29,55,28,95,31,95,30,97,31,211,31,218,31,237,31,237,30,223,31,26,31,81,31,55,31,68,31,207,31,32,31,30,31,60,31,60,30,3,31,22,31,11,31,87,31,141,31,49,31,49,30,239,31,6,31,6,30,6,29,92,31,89,31,132,31,187,31,112,31,100,31,82,31,202,31,136,31,91,31,122,31,242,31,231,31,145,31,227,31,40,31,17,31,136,31,166,31,235,31,41,31,187,31,2,31,182,31,47,31,87,31,87,30,55,31,238,31,238,30,213,31,213,30,218,31,132,31,162,31,102,31,3,31,127,31,27,31,24,31,67,31,218,31,193,31,193,30,113,31,142,31,31,31,159,31,32,31,32,30,229,31,89,31,89,30,89,29,53,31,64,31,83,31,143,31,45,31,58,31,229,31,100,31,95,31,78,31,182,31,165,31,165,30,165,29,241,31,15,31,15,30,15,29,29,31,80,31,36,31,38,31,120,31,77,31,77,30,226,31,226,30,192,31,121,31,233,31,208,31,190,31,190,30,190,29,10,31,72,31,193,31,193,30,129,31,129,30,50,31,199,31,183,31,72,31,139,31,139,30,240,31,117,31,228,31,133,31,194,31,42,31,252,31,116,31,203,31,203,30,199,31,196,31,58,31,184,31,178,31,94,31,9,31,43,31,21,31,21,30,156,31,2,31,2,30,159,31,226,31,226,30,211,31,11,31,90,31,122,31,120,31,14,31,188,31,225,31,235,31,235,30,10,31,38,31,201,31,201,30,118,31,118,30,118,29,143,31,143,30,18,31,250,31,184,31,3,31,16,31,80,31,230,31,212,31,242,31,188,31,188,30,188,29,54,31,193,31,18,31,32,31,114,31,191,31,169,31,169,30,68,31,81,31,81,30,200,31,48,31,98,31,98,30,99,31,2,31,190,31,106,31,106,30,60,31,60,30,27,31,10,31,79,31,207,31,186,31,186,30,86,31,86,30,33,31,18,31,76,31,162,31,1,31,157,31,233,31,221,31,112,31,112,30,174,31,174,30,185,31,23,31,72,31,72,30,193,31,178,31,99,31,229,31,229,30,229,29,185,31,101,31,177,31,177,30,131,31,131,30,255,31,186,31,213,31,189,31,189,30,79,31,172,31,125,31,75,31,116,31,218,31,228,31,228,30,116,31,170,31,50,31,32,31,225,31,225,30,225,31,102,31,68,31,143,31,250,31,224,31,163,31,118,31,11,31,251,31,251,30,251,29,210,31,210,30,73,31,246,31,45,31,61,31,221,31,33,31,227,31,72,31,149,31,217,31,38,31,38,30,65,31,176,31,161,31,17,31,200,31,85,31,85,30,85,29,95,31,95,30,95,29,224,31,224,30,180,31,225,31,69,31,190,31,78,31,186,31,111,31,171,31,25,31,98,31,192,31,192,30,164,31,164,30,121,31,136,31,201,31,19,31,226,31,123,31,123,30,116,31,116,30,243,31,139,31,165,31,165,30,92,31,241,31,56,31,119,31,170,31,184,31,120,31,79,31,79,30,79,29,49,31,62,31,77,31,77,30,5,31,130,31,130,30,130,29,130,28,11,31,237,31,237,30,237,29,90,31,30,31,148,31,247,31,32,31,79,31,116,31,116,30,137,31,15,31,120,31,120,30,189,31,108,31,87,31,75,31,254,31,254,30,40,31,212,31,212,30,159,31,7,31,70,31,208,31,198,31,5,31,169,31,139,31,59,31,203,31,93,31,173,31,101,31,21,31,21,30,21,29,209,31,226,31,226,30,79,31,183,31,168,31,227,31,231,31,112,31,1,31,45,31,222,31,160,31,238,31,157,31,71,31,210,31,16,31,112,31,213,31,75,31,216,31,128,31,254,31,138,31,241,31,204,31,229,31,156,31,234,31,54,31,54,30,26,31,112,31,233,31,233,30,157,31,168,31,149,31,149,30,246,31,41,31,165,31,196,31,184,31,238,31,202,31,127,31,219,31,96,31,86,31,50,31,138,31,253,31,237,31,220,31,34,31,87,31,44,31,58,31,58,30,41,31,126,31,255,31,98,31,147,31,116,31,206,31,90,31,114,31,40,31,242,31,76,31,205,31,205,30,205,31,205,30,205,29,205,28,192,31,55,31,132,31,91,31,120,31,72,31,77,31,46,31,215,31,92,31,37,31,22,31,133,31,126,31,109,31,9,31,39,31,238,31,29,31,179,31,64,31,188,31,188,30,3,31,135,31,141,31,209,31,209,30,139,31,87,31,87,30,75,31,75,30,246,31,246,30,246,29,246,28,208,31,230,31,23,31,65,31,65,30,62,31,153,31,95,31,48,31,48,30,119,31,156,31,252,31,252,30,215,31,222,31,166,31,52,31,95,31,241,31,143,31,143,30,143,29,107,31);

    signal memory_control : std_logic := '0';
    
    constant SCENARIO_ADDRESS : integer := 1234;

    component project_reti_logiche is
        port (
                i_clk : in std_logic;
                i_rst : in std_logic;
                i_start : in std_logic;
                i_add : in std_logic_vector(15 downto 0);
                i_k   : in std_logic_vector(9 downto 0);
                
                o_done : out std_logic;
                
                o_mem_addr : out std_logic_vector(15 downto 0);
                i_mem_data : in  std_logic_vector(7 downto 0);
                o_mem_data : out std_logic_vector(7 downto 0);
                o_mem_we   : out std_logic;
                o_mem_en   : out std_logic
        );
    end component project_reti_logiche;

begin
    UUT : project_reti_logiche
    port map(
                i_clk   => tb_clk,
                i_rst   => tb_rst,
                i_start => tb_start,
                i_add   => tb_add,
                i_k     => tb_k,
                
                o_done => tb_done,
                
                o_mem_addr => exc_o_mem_addr,
                i_mem_data => tb_i_mem_data,
                o_mem_data => exc_o_mem_data,
                o_mem_we   => exc_o_mem_we,
                o_mem_en   => exc_o_mem_en
    );

    -- Clock generation
    tb_clk <= not tb_clk after CLOCK_PERIOD/2;

    -- Process related to the memory
    MEM : process (tb_clk)
    begin
        if tb_clk'event and tb_clk = '1' then
            if tb_o_mem_en = '1' then
                if tb_o_mem_we = '1' then
                    RAM(to_integer(unsigned(tb_o_mem_addr))) <= tb_o_mem_data after 1 ns;
                    tb_i_mem_data <= tb_o_mem_data after 1 ns;
                else
                    tb_i_mem_data <= RAM(to_integer(unsigned(tb_o_mem_addr))) after 1 ns;
                end if;
            end if;
        end if;
    end process;
    
    memory_signal_swapper : process(memory_control, init_o_mem_addr, init_o_mem_data,
                                    init_o_mem_en,  init_o_mem_we,   exc_o_mem_addr,
                                    exc_o_mem_data, exc_o_mem_en, exc_o_mem_we)
    begin
        -- This is necessary for the testbench to work: we swap the memory
        -- signals from the component to the testbench when needed.
    
        tb_o_mem_addr <= init_o_mem_addr;
        tb_o_mem_data <= init_o_mem_data;
        tb_o_mem_en   <= init_o_mem_en;
        tb_o_mem_we   <= init_o_mem_we;

        if memory_control = '1' then
            tb_o_mem_addr <= exc_o_mem_addr;
            tb_o_mem_data <= exc_o_mem_data;
            tb_o_mem_en   <= exc_o_mem_en;
            tb_o_mem_we   <= exc_o_mem_we;
        end if;
    end process;
    
    -- This process provides the correct scenario on the signal controlled by the TB
    create_scenario : process
    begin
        wait for 50 ns;

        -- Signal initialization and reset of the component
        tb_start <= '0';
        tb_add <= (others=>'0');
        tb_k   <= (others=>'0');
        tb_rst <= '1';
        
        -- Wait some time for the component to reset...
        wait for 50 ns;
        
        tb_rst <= '0';
        memory_control <= '0';  -- Memory controlled by the testbench
        
        wait until falling_edge(tb_clk); -- Skew the testbench transitions with respect to the clock

        -- Configure the memory        
        for i in 0 to SCENARIO_LENGTH*2-1 loop
            init_o_mem_addr<= std_logic_vector(to_unsigned(SCENARIO_ADDRESS+i, 16));
            init_o_mem_data<= std_logic_vector(to_unsigned(scenario_input(i),8));
            init_o_mem_en  <= '1';
            init_o_mem_we  <= '1';
            wait until rising_edge(tb_clk);   
        end loop;
        
        wait until falling_edge(tb_clk);

        memory_control <= '1';  -- Memory controlled by the component
        
        tb_add <= std_logic_vector(to_unsigned(SCENARIO_ADDRESS, 16));
        tb_k   <= std_logic_vector(to_unsigned(SCENARIO_LENGTH, 10));
        
        tb_start <= '1';

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        wait for 5 ns;
        
        tb_start <= '0';
        
        wait;
        
    end process;

    -- Process without sensitivity list designed to test the actual component.
    test_routine : process
    begin

        wait until tb_rst = '1';
        wait for 25 ns;
        assert tb_done = '0' report "TEST FALLITO o_done !=0 during reset" severity failure;
        wait until tb_rst = '0';

        wait until falling_edge(tb_clk);
        assert tb_done = '0' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        
        wait until rising_edge(tb_start);

        while tb_done /= '1' loop                
            wait until rising_edge(tb_clk);
        end loop;

        assert tb_o_mem_en = '0' or tb_o_mem_we = '0' report "TEST FALLITO o_mem_en !=0 memory should not be written after done." severity failure;

        for i in 0 to SCENARIO_LENGTH*2-1 loop
            assert RAM(SCENARIO_ADDRESS+i) = std_logic_vector(to_unsigned(scenario_full(i),8)) report "TEST FALLITO @ OFFSET=" & integer'image(i) & " expected= " & integer'image(scenario_full(i)) & " actual=" & integer'image(to_integer(unsigned(RAM(i)))) severity failure;
        end loop;

        wait until falling_edge(tb_start);
        assert tb_done = '1' report "TEST FALLITO o_done !=0 after reset before start" severity failure;
        wait until falling_edge(tb_done);

        assert false report "Simulation Ended! TEST PASSATO (EXAMPLE)" severity failure;
    end process;

end architecture;
